-- Xilinx Vhdl netlist produced by netgen application (version G.25a)
-- Command       : -intstyle ise -s 6 -pcf network.pcf -ngm network.ngm -fn -rpw 100 -tpw 0 -ar Structure -xon false -w -ofmt vhdl -sim network.ncd testsuite_PR.vhd 
-- Input file    : network.ncd
-- Output file   : testsuite_PR.vhd
-- Design name   : network
-- # of Entities : 1
-- Xilinx        : C:/Xilinx
-- Device        : 2s200epq208-6 (PRODUCTION 1.17 2003-09-30)

-- This vhdl netlist is a simulation model and uses simulation 
-- primitives which may not represent the true implementation of the 
-- device, however the netlist is functionally correct and should not 
-- be modified. This file cannot be synthesized and should only be used 
-- with supported simulation tools.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library SIMPRIM;
use SIMPRIM.VCOMPONENTS.ALL;
use SIMPRIM.VPACKAGE.ALL;

entity network is
  port (
    DOUTEN : out STD_LOGIC; 
    MCLK : out STD_LOGIC; 
    LED100 : out STD_LOGIC; 
    LED1000 : out STD_LOGIC; 
    PHYRESET : out STD_LOGIC; 
    GTX_CLK : out STD_LOGIC; 
    LEDACT : out STD_LOGIC; 
    SOUT : out STD_LOGIC; 
    MWE : out STD_LOGIC; 
    TX_EN : out STD_LOGIC; 
    LEDDPX : out STD_LOGIC; 
    LEDTX : out STD_LOGIC; 
    LEDRX : out STD_LOGIC; 
    LEDPOWER : out STD_LOGIC; 
    MDC : out STD_LOGIC; 
    MDIO : inout STD_LOGIC; 
    SCS : in STD_LOGIC := 'X'; 
    NEXTFRAME : in STD_LOGIC := 'X'; 
    SCLK : in STD_LOGIC := 'X'; 
    DINEN : in STD_LOGIC := 'X'; 
    CLKIOIN : in STD_LOGIC := 'X'; 
    RX_CLK : in STD_LOGIC := 'X'; 
    NEWFRAME : in STD_LOGIC := 'X'; 
    RESET : in STD_LOGIC := 'X'; 
    CLKIN : in STD_LOGIC := 'X'; 
    RX_ER : in STD_LOGIC := 'X'; 
    RX_DV : in STD_LOGIC := 'X'; 
    SIN : in STD_LOGIC := 'X'; 
    DOUT : out STD_LOGIC_VECTOR ( 15 downto 0 ); 
    TXD : out STD_LOGIC_VECTOR ( 7 downto 0 ); 
    MA : out STD_LOGIC_VECTOR ( 16 downto 0 ); 
    MD : inout STD_LOGIC_VECTOR ( 31 downto 0 ); 
    RXD : in STD_LOGIC_VECTOR ( 7 downto 0 ); 
    DIN : in STD_LOGIC_VECTOR ( 15 downto 0 ) 
  );
end network;

architecture Structure of network is
  signal rx_input_fifo_fifo_N2444 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2443 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2442 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2441 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5329 : STD_LOGIC; 
  signal rx_input_ince : STD_LOGIC; 
  signal rx_input_fifo_fifo_full : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2364 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4912 : STD_LOGIC; 
  signal rx_input_fifo_fifo_BU431_O : STD_LOGIC; 
  signal clkrx : STD_LOGIC; 
  signal rx_input_fifo_RESET_1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2417 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2362 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4903 : STD_LOGIC; 
  signal GTX_CLK_OBUF : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2478 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2418 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2428 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2477 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2427 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3982 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2397 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2398 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2419 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4905 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2480 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2420 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2430 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2479 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2429 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2438 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2437 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2467 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2468 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6355 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2448 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2447 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3972 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2400 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2399 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2421 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4907 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2482 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2422 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2432 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2481 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2431 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2439 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2440 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2469 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2470 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6347 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2450 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2449 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5330 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3962 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2401 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2402 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2423 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4909 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2484 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2424 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2434 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2483 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2433 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2472 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2471 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6339 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2452 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2451 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3952 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2403 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2404 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2486 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2426 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2436 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2485 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2425 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2435 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2473 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2474 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6331 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2454 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2453 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2405 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2406 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2445 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2446 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2475 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2476 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2456 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2455 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N23 : STD_LOGIC; 
  signal rx_input_rx_nearf : STD_LOGIC; 
  signal rx_input_fifo_rd_en : STD_LOGIC; 
  signal rx_input_fifo_fifo_empty : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3646 : STD_LOGIC; 
  signal rx_input_fifo_fifo_BU216_O : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3637 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2498 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2497 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2852 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3639 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2500 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2499 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2842 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3641 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2502 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2501 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N16 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N17 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2832 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3643 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2504 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2503 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N19 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N18 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2822 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2506 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2505 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N21 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N20 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N22 : STD_LOGIC; 
  signal slowclock_n0002 : STD_LOGIC; 
  signal slowclock_n0005 : STD_LOGIC; 
  signal RESET_IBUF_2 : STD_LOGIC; 
  signal tx_input_n0021 : STD_LOGIC; 
  signal mac_control_CHOICE1616 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_153 : STD_LOGIC; 
  signal mac_control_CHOICE1609 : STD_LOGIC; 
  signal mac_control_N81797 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_152 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_150 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151 : STD_LOGIC; 
  signal mac_control_n0039 : STD_LOGIC; 
  signal rx_input_GMII_rx_dvl : STD_LOGIC; 
  signal rx_input_GMII_ro : STD_LOGIC; 
  signal rx_input_GMII_rx_dvll : STD_LOGIC; 
  signal rx_input_GMII_dvdelta : STD_LOGIC; 
  signal tx_input_n0020 : STD_LOGIC; 
  signal tx_input_addr_27 : STD_LOGIC; 
  signal tx_input_addr_26 : STD_LOGIC; 
  signal tx_input_n0023 : STD_LOGIC; 
  signal tx_input_addr_29 : STD_LOGIC; 
  signal tx_input_addr_28 : STD_LOGIC; 
  signal tx_input_addr_31 : STD_LOGIC; 
  signal tx_input_addr_30 : STD_LOGIC; 
  signal mac_control_CHOICE1593 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_165 : STD_LOGIC; 
  signal mac_control_CHOICE1586 : STD_LOGIC; 
  signal mac_control_N81777 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_164 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_162 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163 : STD_LOGIC; 
  signal mac_control_n0041 : STD_LOGIC; 
  signal rx_input_endf : STD_LOGIC; 
  signal rx_input_invalid : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd2 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd1 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16 : STD_LOGIC; 
  signal rx_input_memio_brdy : STD_LOGIC; 
  signal rx_input_RESET_1 : STD_LOGIC; 
  signal rxucast : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxucastl : STD_LOGIC; 
  signal mac_control_n0029 : STD_LOGIC; 
  signal mac_control_n0030 : STD_LOGIC; 
  signal mac_control_n0031 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_11_58 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_10_59 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_13_56 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_12_57 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_15_54 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_14_55 : STD_LOGIC; 
  signal rx_output_denll : STD_LOGIC; 
  signal rx_output_fifo_empty : STD_LOGIC; 
  signal rx_output_fifo_N2579 : STD_LOGIC; 
  signal rx_output_fifo_N18 : STD_LOGIC; 
  signal clkio : STD_LOGIC; 
  signal rx_output_fifo_reset : STD_LOGIC; 
  signal rx_output_invalid : STD_LOGIC; 
  signal rx_output_fifo_N1515 : STD_LOGIC; 
  signal memcontroller_n0005 : STD_LOGIC; 
  signal mac_control_bitcnt_104 : STD_LOGIC; 
  signal mac_control_bitcnt_106 : STD_LOGIC; 
  signal mac_control_bitcnt_105 : STD_LOGIC; 
  signal mac_control_Ker52136_2 : STD_LOGIC; 
  signal memcontroller_n0006 : STD_LOGIC; 
  signal RESET_IBUF : STD_LOGIC; 
  signal slowclock_rxfifowerrl : STD_LOGIC; 
  signal clkslen : STD_LOGIC; 
  signal rxfifowerrsr : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2 : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_25_Xo_1_1_2 : STD_LOGIC; 
  signal slowclock_rxoferrl : STD_LOGIC; 
  signal rxoferrsr : STD_LOGIC; 
  signal tx_output_cs_FFd9 : STD_LOGIC; 
  signal tx_output_cs_FFd10 : STD_LOGIC; 
  signal tx_output_cs_FFd11 : STD_LOGIC; 
  signal tx_output_cs_FFd13 : STD_LOGIC; 
  signal tx_output_cs_FFd14 : STD_LOGIC; 
  signal tx_output_cs_Out1160_2 : STD_LOGIC; 
  signal tx_output_CHOICE1641 : STD_LOGIC; 
  signal tx_output_cs_Out1160_SW0_1 : STD_LOGIC; 
  signal tx_output_CHOICE1634 : STD_LOGIC; 
  signal txfifowerr : STD_LOGIC; 
  signal slowclock_txfifowerrl : STD_LOGIC; 
  signal rxfifofull : STD_LOGIC; 
  signal rx_input_memio_fifofulll : STD_LOGIC; 
  signal rx_input_memio_n0032 : STD_LOGIC; 
  signal rx_output_nf : STD_LOGIC; 
  signal rx_output_nfl : STD_LOGIC; 
  signal mac_control_Mshreg_sinlll_102 : STD_LOGIC; 
  signal mac_control_n0010 : STD_LOGIC; 
  signal tx_input_CHOICE1710 : STD_LOGIC; 
  signal tx_input_CHOICE1729 : STD_LOGIC; 
  signal tx_input_CHOICE1717 : STD_LOGIC; 
  signal tx_input_CHOICE1732 : STD_LOGIC; 
  signal tx_input_Ker34480137_2 : STD_LOGIC; 
  signal tx_input_N81681 : STD_LOGIC; 
  signal tx_input_cs_FFd11 : STD_LOGIC; 
  signal tx_input_cs_FFd6 : STD_LOGIC; 
  signal tx_input_N69350 : STD_LOGIC; 
  signal tx_input_N73800 : STD_LOGIC; 
  signal RESET_IBUF_1 : STD_LOGIC; 
  signal tx_input_cs_FFd10 : STD_LOGIC; 
  signal mac_control_n0011 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_34 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_32 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n001124_2 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81705 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2526 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd10 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1451 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1447 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd15 : STD_LOGIC; 
  signal rx_input_memio_N81863 : STD_LOGIC; 
  signal tx_output_n0025 : STD_LOGIC; 
  signal tx_output_cs_FFd16 : STD_LOGIC; 
  signal tx_output_crc_3_Q : STD_LOGIC; 
  signal mac_control_PHY_status_n00151_1 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0016 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2546 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2532 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N82069 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N82067 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2555 : STD_LOGIC; 
  signal rx_input_memio_n0030 : STD_LOGIC; 
  signal rx_input_memio_N70785 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd3 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd1 : STD_LOGIC; 
  signal mac_control_n0103 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_18_42_SW0_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_20_42_SW0_1 : STD_LOGIC; 
  signal rxf : STD_LOGIC; 
  signal mac_control_n0025 : STD_LOGIC; 
  signal rxoferr : STD_LOGIC; 
  signal rx_input_memio_crcrst : STD_LOGIC; 
  signal mac_control_sclkl : STD_LOGIC; 
  signal mac_control_N52198 : STD_LOGIC; 
  signal mac_control_sclkll : STD_LOGIC; 
  signal rx_input_memio_n0044 : STD_LOGIC; 
  signal rx_input_memio_n0045 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N37245 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd5 : STD_LOGIC; 
  signal MDC_OBUF : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_37 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0010 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N37240 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2562 : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2 : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_18_Xo_2_1_2 : STD_LOGIC; 
  signal tx_output_ltxen3 : STD_LOGIC; 
  signal tx_output_ltxen2 : STD_LOGIC; 
  signal txf : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd2 : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd1 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1462 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1455 : STD_LOGIC; 
  signal rx_input_fifo_control_n0008 : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4 : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd3 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1458 : STD_LOGIC; 
  signal rx_output_cs_FFd1 : STD_LOGIC; 
  signal rx_output_cs_FFd11 : STD_LOGIC; 
  signal rx_output_cs_FFd5 : STD_LOGIC; 
  signal rx_output_n0018 : STD_LOGIC; 
  signal rx_output_N33107 : STD_LOGIC; 
  signal rx_output_cs_FFd9 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1483 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1518 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1465 : STD_LOGIC; 
  signal tx_output_bcnt_42 : STD_LOGIC; 
  signal tx_output_bcnt_43 : STD_LOGIC; 
  signal tx_output_bcnt_44 : STD_LOGIC; 
  signal tx_output_bcnt_45 : STD_LOGIC; 
  signal tx_output_CHOICE1656 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1490 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1511 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1521 : STD_LOGIC; 
  signal tx_output_bcnt_50 : STD_LOGIC; 
  signal tx_output_bcnt_51 : STD_LOGIC; 
  signal tx_output_bcnt_52 : STD_LOGIC; 
  signal tx_output_bcnt_53 : STD_LOGIC; 
  signal tx_output_bcnt_41 : STD_LOGIC; 
  signal tx_output_CHOICE1664 : STD_LOGIC; 
  signal tx_output_CHOICE1671 : STD_LOGIC; 
  signal tx_output_N81677 : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4_In_2 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1497 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1514 : STD_LOGIC; 
  signal tx_output_bcnt_46 : STD_LOGIC; 
  signal tx_output_bcnt_47 : STD_LOGIC; 
  signal tx_output_bcnt_48 : STD_LOGIC; 
  signal tx_output_bcnt_49 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1476 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1504 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1500 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1507 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1493 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1486 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1469 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1479 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1472 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81600 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N69488 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd3 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd4 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1550 : STD_LOGIC; 
  signal tx_output_crc_6_Q : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd5 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd7 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd6 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1551 : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_4_Xo_1_1_2 : STD_LOGIC; 
  signal mac_control_newcmd : STD_LOGIC; 
  signal mac_control_N69420 : STD_LOGIC; 
  signal mac_control_N52220 : STD_LOGIC; 
  signal mac_control_N52153 : STD_LOGIC; 
  signal mac_control_n0034 : STD_LOGIC; 
  signal mac_control_bitcnt_108 : STD_LOGIC; 
  signal mac_control_bitcnt_107 : STD_LOGIC; 
  signal mac_control_n001220_1 : STD_LOGIC; 
  signal mac_control_CHOICE1171 : STD_LOGIC; 
  signal mac_control_n001220_SW0_1 : STD_LOGIC; 
  signal mac_control_N52138 : STD_LOGIC; 
  signal mac_control_N70898 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0004_2 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0004 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd3 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd2 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0079 : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_2 : STD_LOGIC; 
  signal tx_input_den : STD_LOGIC; 
  signal tx_input_N34493 : STD_LOGIC; 
  signal tx_input_cs_FFd12 : STD_LOGIC; 
  signal rx_output_cs_FFd19 : STD_LOGIC; 
  signal rx_output_N69253 : STD_LOGIC; 
  signal rx_output_cs_FFd17 : STD_LOGIC; 
  signal rx_output_n0043 : STD_LOGIC; 
  signal tx_output_crc_7_Q : STD_LOGIC; 
  signal mac_control_PHY_status_n0011 : STD_LOGIC; 
  signal mac_control_N52111 : STD_LOGIC; 
  signal mac_control_N52132 : STD_LOGIC; 
  signal mac_control_N82133 : STD_LOGIC; 
  signal mac_control_N82121 : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_25_42_SW0_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_30_42_SW0_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_28_42_SW0_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_22_42_SW0_1 : STD_LOGIC; 
  signal txfifofull : STD_LOGIC; 
  signal tx_input_fifofulll : STD_LOGIC; 
  signal tx_output_crc_8_Q : STD_LOGIC; 
  signal rx_input_memio_CHOICE2946 : STD_LOGIC; 
  signal rx_input_memio_n0059143_2 : STD_LOGIC; 
  signal rx_input_memio_n0059143_SW0_2 : STD_LOGIC; 
  signal rx_input_memio_CHOICE2951 : STD_LOGIC; 
  signal rx_input_memio_crcequal : STD_LOGIC; 
  signal mac_control_CHOICE2449 : STD_LOGIC; 
  signal mac_control_CHOICE2432 : STD_LOGIC; 
  signal mac_control_n0085 : STD_LOGIC; 
  signal mac_control_n0060 : STD_LOGIC; 
  signal mac_control_N81665 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd1 : STD_LOGIC; 
  signal mac_control_PHY_status_n0015 : STD_LOGIC; 
  signal mac_control_PHY_status_phyaddrws : STD_LOGIC; 
  signal mac_control_bitcnt_109 : STD_LOGIC; 
  signal mac_control_sclkdeltall : STD_LOGIC; 
  signal mac_control_N82019 : STD_LOGIC; 
  signal mac_control_N82013 : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2 : STD_LOGIC; 
  signal rx_output_fifo_nearfull : STD_LOGIC; 
  signal tx_output_crc_9_Q : STD_LOGIC; 
  signal tx_input_addr_17 : STD_LOGIC; 
  signal tx_input_addr_16 : STD_LOGIC; 
  signal tx_input_mrw : STD_LOGIC; 
  signal tx_input_addr_19 : STD_LOGIC; 
  signal tx_input_addr_18 : STD_LOGIC; 
  signal tx_input_addr_21 : STD_LOGIC; 
  signal tx_input_addr_20 : STD_LOGIC; 
  signal tx_input_addr_23 : STD_LOGIC; 
  signal tx_input_addr_22 : STD_LOGIC; 
  signal tx_input_addr_25 : STD_LOGIC; 
  signal tx_input_addr_24 : STD_LOGIC; 
  signal rx_output_cs_FFd13 : STD_LOGIC; 
  signal rx_output_cs_FFd12 : STD_LOGIC; 
  signal rx_output_cs_FFd15 : STD_LOGIC; 
  signal rx_output_cs_FFd14 : STD_LOGIC; 
  signal rx_output_cs_FFd16 : STD_LOGIC; 
  signal rx_output_cs_FFd8 : STD_LOGIC; 
  signal rx_output_cs_FFd7 : STD_LOGIC; 
  signal rx_output_ceinl : STD_LOGIC; 
  signal rx_output_n0033 : STD_LOGIC; 
  signal rx_output_cs_FFd10 : STD_LOGIC; 
  signal rx_output_n0034 : STD_LOGIC; 
  signal rxfsr : STD_LOGIC; 
  signal mac_control_rxf_cross : STD_LOGIC; 
  signal tx_input_cs_FFd7 : STD_LOGIC; 
  signal tx_input_cs_FFd2 : STD_LOGIC; 
  signal mac_control_N52251 : STD_LOGIC; 
  signal mac_control_sclkdelta : STD_LOGIC; 
  signal mac_control_phyrstcnt_129 : STD_LOGIC; 
  signal mac_control_phyrstcnt_111 : STD_LOGIC; 
  signal mac_control_phyrstcnt_130 : STD_LOGIC; 
  signal mac_control_phyrstcnt_131 : STD_LOGIC; 
  signal mac_control_CHOICE2746 : STD_LOGIC; 
  signal mac_control_CHOICE2966 : STD_LOGIC; 
  signal mac_control_phyrstcnt_125 : STD_LOGIC; 
  signal mac_control_phyrstcnt_126 : STD_LOGIC; 
  signal mac_control_phyrstcnt_127 : STD_LOGIC; 
  signal mac_control_phyrstcnt_128 : STD_LOGIC; 
  signal mac_control_CHOICE2739 : STD_LOGIC; 
  signal mac_control_CHOICE2963 : STD_LOGIC; 
  signal mac_control_phyrstcnt_136 : STD_LOGIC; 
  signal mac_control_phyrstcnt_137 : STD_LOGIC; 
  signal mac_control_phyrstcnt_138 : STD_LOGIC; 
  signal mac_control_phyrstcnt_139 : STD_LOGIC; 
  signal mac_control_CHOICE2762 : STD_LOGIC; 
  signal mac_control_CHOICE2974 : STD_LOGIC; 
  signal mac_control_phyrstcnt_121 : STD_LOGIC; 
  signal mac_control_phyrstcnt_122 : STD_LOGIC; 
  signal mac_control_phyrstcnt_123 : STD_LOGIC; 
  signal mac_control_phyrstcnt_124 : STD_LOGIC; 
  signal mac_control_CHOICE2731 : STD_LOGIC; 
  signal mac_control_phyrstcnt_120 : STD_LOGIC; 
  signal mac_control_phyrstcnt_119 : STD_LOGIC; 
  signal mac_control_phyrstcnt_110 : STD_LOGIC; 
  signal mac_control_CHOICE2732 : STD_LOGIC; 
  signal mac_control_phyrstcnt_132 : STD_LOGIC; 
  signal mac_control_phyrstcnt_133 : STD_LOGIC; 
  signal mac_control_phyrstcnt_134 : STD_LOGIC; 
  signal mac_control_phyrstcnt_135 : STD_LOGIC; 
  signal mac_control_CHOICE2971 : STD_LOGIC; 
  signal mac_control_phyrstcnt_112 : STD_LOGIC; 
  signal mac_control_phyrstcnt_140 : STD_LOGIC; 
  signal mac_control_phyrstcnt_113 : STD_LOGIC; 
  signal mac_control_phyrstcnt_114 : STD_LOGIC; 
  signal mac_control_CHOICE2770 : STD_LOGIC; 
  signal mac_control_CHOICE2978 : STD_LOGIC; 
  signal mac_control_phyrstcnt_115 : STD_LOGIC; 
  signal mac_control_phyrstcnt_116 : STD_LOGIC; 
  signal mac_control_phyrstcnt_117 : STD_LOGIC; 
  signal mac_control_phyrstcnt_118 : STD_LOGIC; 
  signal mac_control_CHOICE2777 : STD_LOGIC; 
  signal mac_control_CHOICE2981 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N72822 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_142 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_144 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145 : STD_LOGIC; 
  signal mac_control_ledtx_rst : STD_LOGIC; 
  signal mac_control_N73201 : STD_LOGIC; 
  signal mac_control_n0038 : STD_LOGIC; 
  signal tx_output_crc_0_Q : STD_LOGIC; 
  signal mac_control_ledrx_cnt_154 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_156 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_146 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_148 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149 : STD_LOGIC; 
  signal mac_control_CHOICE2755 : STD_LOGIC; 
  signal mac_control_n0035194_SW0_2 : STD_LOGIC; 
  signal mac_control_ledrx_rst : STD_LOGIC; 
  signal mac_control_N73084 : STD_LOGIC; 
  signal mac_control_n0040 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_158 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_160 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161 : STD_LOGIC; 
  signal slowclock_rxfl : STD_LOGIC; 
  signal slowclock_txfl : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_14_Xo_3_1_2 : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_5_Xo_1_1_2 : STD_LOGIC; 
  signal mac_control_N52125 : STD_LOGIC; 
  signal mac_control_N52244 : STD_LOGIC; 
  signal mac_control_CHOICE2442 : STD_LOGIC; 
  signal mac_control_CHOICE2436 : STD_LOGIC; 
  signal mac_control_CHOICE2448 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_1_68 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_0_69 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_3_66 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_2_67 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_5_64 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_4_65 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_7_62 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_6_63 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_9_60 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_8_61 : STD_LOGIC; 
  signal mac_control_N82117 : STD_LOGIC; 
  signal mac_control_CHOICE2480 : STD_LOGIC; 
  signal mac_control_CHOICE2474 : STD_LOGIC; 
  signal mac_control_CHOICE2486 : STD_LOGIC; 
  signal mac_control_CHOICE2487 : STD_LOGIC; 
  signal mac_control_N82129 : STD_LOGIC; 
  signal rx_output_N69852 : STD_LOGIC; 
  signal rx_input_memio_n0034 : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_25_Xo_1_1_2 : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_4_Xo_1_1_2 : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_5_Xo_1_1_2 : STD_LOGIC; 
  signal txfsr : STD_LOGIC; 
  signal mac_control_txf_cross : STD_LOGIC; 
  signal rx_output_cs_FFd6 : STD_LOGIC; 
  signal rx_output_fifo_full : STD_LOGIC; 
  signal rx_output_N70424 : STD_LOGIC; 
  signal rx_output_N69800 : STD_LOGIC; 
  signal rx_output_N69904 : STD_LOGIC; 
  signal rx_output_cs_FFd4 : STD_LOGIC; 
  signal rx_output_cs_FFd3 : STD_LOGIC; 
  signal rx_output_cs_FFd2 : STD_LOGIC; 
  signal rx_output_CHOICE1557 : STD_LOGIC; 
  signal rx_output_CHOICE1525 : STD_LOGIC; 
  signal rx_output_CHOICE1528 : STD_LOGIC; 
  signal rx_output_denl : STD_LOGIC; 
  signal rx_output_N69956 : STD_LOGIC; 
  signal mac_control_lrxbcast : STD_LOGIC; 
  signal rxbcast : STD_LOGIC; 
  signal rx_output_N70008 : STD_LOGIC; 
  signal mac_control_CHOICE2470 : STD_LOGIC; 
  signal mac_control_N81637 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2503 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2497 : STD_LOGIC; 
  signal tx_output_crc_1_Q : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2511 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2512 : STD_LOGIC; 
  signal rx_output_N70112 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2513 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_sout498_2 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_3_108_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_3_96_1 : STD_LOGIC; 
  signal mac_control_CHOICE1821 : STD_LOGIC; 
  signal mac_control_CHOICE1814 : STD_LOGIC; 
  signal mac_control_CHOICE1817 : STD_LOGIC; 
  signal mac_control_N82074 : STD_LOGIC; 
  signal mac_control_CHOICE1877 : STD_LOGIC; 
  signal mac_control_CHOICE1870 : STD_LOGIC; 
  signal mac_control_CHOICE1873 : STD_LOGIC; 
  signal mac_control_N82082 : STD_LOGIC; 
  signal rx_output_N70060 : STD_LOGIC; 
  signal tx_input_cs_FFd4 : STD_LOGIC; 
  signal rx_output_N70164 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1403 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1392 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1399 : STD_LOGIC; 
  signal tx_output_CHOICE1303 : STD_LOGIC; 
  signal tx_output_CHOICE1380 : STD_LOGIC; 
  signal tx_output_CHOICE1385 : STD_LOGIC; 
  signal tx_output_CHOICE1336 : STD_LOGIC; 
  signal tx_output_CHOICE1369 : STD_LOGIC; 
  signal tx_output_CHOICE1374 : STD_LOGIC; 
  signal mac_control_N52163 : STD_LOGIC; 
  signal mac_control_N82001 : STD_LOGIC; 
  signal tx_output_CHOICE1314 : STD_LOGIC; 
  signal tx_output_CHOICE1358 : STD_LOGIC; 
  signal tx_output_CHOICE1363 : STD_LOGIC; 
  signal tx_output_CHOICE1341 : STD_LOGIC; 
  signal tx_output_CHOICE1325 : STD_LOGIC; 
  signal tx_output_CHOICE1347 : STD_LOGIC; 
  signal tx_output_CHOICE1352 : STD_LOGIC; 
  signal tx_output_CHOICE1330 : STD_LOGIC; 
  signal tx_output_CHOICE1319 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0051_2 : STD_LOGIC; 
  signal rx_input_memio_addrchk_validbcast : STD_LOGIC; 
  signal tx_output_CHOICE1308 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0052_2 : STD_LOGIC; 
  signal rx_input_memio_addrchk_validucast : STD_LOGIC; 
  signal mac_control_lrxmcast : STD_LOGIC; 
  signal rxmcast : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1774 : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1781 : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1796 : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1789 : STD_LOGIC; 
  signal rx_fifocheck_n0003 : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1797 : STD_LOGIC; 
  signal rx_fifocheck_N74128 : STD_LOGIC; 
  signal mac_control_lrxucast : STD_LOGIC; 
  signal tx_output_cs_FFd8 : STD_LOGIC; 
  signal tx_output_crcenl : STD_LOGIC; 
  signal tx_output_cs_FFd6 : STD_LOGIC; 
  signal tx_output_cs_FFd15 : STD_LOGIC; 
  signal tx_output_cs_FFd17 : STD_LOGIC; 
  signal tx_output_cs_FFd12 : STD_LOGIC; 
  signal tx_output_CHOICE1679 : STD_LOGIC; 
  signal tx_output_cs_FFd5 : STD_LOGIC; 
  signal tx_output_cs_FFd4 : STD_LOGIC; 
  signal tx_output_cs_FFd7 : STD_LOGIC; 
  signal tx_output_cs_FFd3 : STD_LOGIC; 
  signal tx_output_N81625 : STD_LOGIC; 
  signal tx_output_CHOICE1683 : STD_LOGIC; 
  signal tx_output_cs_FFd2 : STD_LOGIC; 
  signal tx_output_cs_FFd1 : STD_LOGIC; 
  signal tx_output_CHOICE1686 : STD_LOGIC; 
  signal tx_output_cs_Out13_2 : STD_LOGIC; 
  signal mac_control_phyrstcnt_141 : STD_LOGIC; 
  signal mac_control_N81689 : STD_LOGIC; 
  signal mac_control_N79380 : STD_LOGIC; 
  signal mac_control_PHY_status_rwl : STD_LOGIC; 
  signal rx_input_GMII_rx_of : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2 : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_30_Xo_1_1_2 : STD_LOGIC; 
  signal rx_input_memio_CHOICE2922 : STD_LOGIC; 
  signal rx_input_memio_CHOICE2913 : STD_LOGIC; 
  signal rx_input_memio_CHOICE2917 : STD_LOGIC; 
  signal rx_input_memio_CHOICE2926 : STD_LOGIC; 
  signal slowclock_lclken : STD_LOGIC; 
  signal rx_input_memio_CHOICE2941 : STD_LOGIC; 
  signal rx_input_memio_CHOICE2934 : STD_LOGIC; 
  signal rx_input_memio_crc_0_Q : STD_LOGIC; 
  signal mac_control_PHY_status_n0021 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_29_42_SW0_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_26_42_SW0_1 : STD_LOGIC; 
  signal tx_output_N81669 : STD_LOGIC; 
  signal mac_control_N52100 : STD_LOGIC; 
  signal mac_control_N52143 : STD_LOGIC; 
  signal mac_control_n0013 : STD_LOGIC; 
  signal mac_control_N52236 : STD_LOGIC; 
  signal mac_control_CHOICE2186 : STD_LOGIC; 
  signal mac_control_CHOICE2183 : STD_LOGIC; 
  signal mac_control_N81789 : STD_LOGIC; 
  signal mac_control_n0016 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_292 : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_103 : STD_LOGIC; 
  signal mac_control_rxphyerr_rst : STD_LOGIC; 
  signal mac_control_n0050 : STD_LOGIC; 
  signal mac_control_txf_rst : STD_LOGIC; 
  signal mac_control_n0042 : STD_LOGIC; 
  signal rxphyerrsr : STD_LOGIC; 
  signal mac_control_n0051 : STD_LOGIC; 
  signal mac_control_n0043 : STD_LOGIC; 
  signal mac_control_CHOICE2959 : STD_LOGIC; 
  signal mac_control_CHOICE2960 : STD_LOGIC; 
  signal mac_control_rxoferr_rst : STD_LOGIC; 
  signal mac_control_n0052 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_26_77_1 : STD_LOGIC; 
  signal mac_control_n0037 : STD_LOGIC; 
  signal mac_control_n0036 : STD_LOGIC; 
  signal mac_control_rxf_rst : STD_LOGIC; 
  signal mac_control_n0044 : STD_LOGIC; 
  signal tx_input_DONE : STD_LOGIC; 
  signal mac_control_n0053 : STD_LOGIC; 
  signal mac_control_n0045 : STD_LOGIC; 
  signal mac_control_rxcrcerr_rst : STD_LOGIC; 
  signal mac_control_n0054 : STD_LOGIC; 
  signal mac_control_txfifowerr_rst : STD_LOGIC; 
  signal mac_control_n0046 : STD_LOGIC; 
  signal rxcrcerrsr : STD_LOGIC; 
  signal mac_control_n0055 : STD_LOGIC; 
  signal txfifowerrsr : STD_LOGIC; 
  signal mac_control_n0047 : STD_LOGIC; 
  signal mac_control_rxfifowerr_rst : STD_LOGIC; 
  signal mac_control_n0048 : STD_LOGIC; 
  signal mac_control_N81693 : STD_LOGIC; 
  signal mac_control_CHOICE2801 : STD_LOGIC; 
  signal mac_control_n0080 : STD_LOGIC; 
  signal mac_control_CHOICE2810 : STD_LOGIC; 
  signal mac_control_n0049 : STD_LOGIC; 
  signal mac_control_N52228 : STD_LOGIC; 
  signal mac_control_n0073 : STD_LOGIC; 
  signal mac_control_n0081 : STD_LOGIC; 
  signal mac_control_CHOICE2054 : STD_LOGIC; 
  signal mac_control_n0074 : STD_LOGIC; 
  signal mac_control_sclkdeltal : STD_LOGIC; 
  signal mac_control_N52118 : STD_LOGIC; 
  signal mac_control_n0082 : STD_LOGIC; 
  signal mac_control_CHOICE2645 : STD_LOGIC; 
  signal mac_control_n0083 : STD_LOGIC; 
  signal mac_control_n0076 : STD_LOGIC; 
  signal mac_control_CHOICE2064 : STD_LOGIC; 
  signal mac_control_n0084 : STD_LOGIC; 
  signal mac_control_CHOICE2711 : STD_LOGIC; 
  signal mac_control_n0077 : STD_LOGIC; 
  signal mac_control_CHOICE2790 : STD_LOGIC; 
  signal mac_control_n0087 : STD_LOGIC; 
  signal mac_control_n0086 : STD_LOGIC; 
  signal mac_control_n0078 : STD_LOGIC; 
  signal mac_control_n0079 : STD_LOGIC; 
  signal mac_control_CHOICE2793 : STD_LOGIC; 
  signal slowclock_rxcrcerrl : STD_LOGIC; 
  signal mac_control_CHOICE2857 : STD_LOGIC; 
  signal mac_control_CHOICE2854 : STD_LOGIC; 
  signal mac_control_CHOICE2600 : STD_LOGIC; 
  signal mac_control_N81785 : STD_LOGIC; 
  signal mac_control_CHOICE1905 : STD_LOGIC; 
  signal mac_control_CHOICE1898 : STD_LOGIC; 
  signal mac_control_CHOICE1901 : STD_LOGIC; 
  signal mac_control_N82086 : STD_LOGIC; 
  signal mac_control_CHOICE1849 : STD_LOGIC; 
  signal mac_control_CHOICE1842 : STD_LOGIC; 
  signal mac_control_CHOICE1845 : STD_LOGIC; 
  signal mac_control_N82078 : STD_LOGIC; 
  signal mac_control_PHY_status_miirw : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE1201 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_sts : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd4 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n001124_SW0_2 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE1541 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0030 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0031 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0032 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1424 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0027 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0028 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1431 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0029 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1427 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1417 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1406 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1434 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1438 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1420 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1410 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1441 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1413 : STD_LOGIC; 
  signal rx_output_ldouten2 : STD_LOGIC; 
  signal tx_output_n0006 : STD_LOGIC; 
  signal rx_input_memio_crc_1_Q : STD_LOGIC; 
  signal tx_output_N81617 : STD_LOGIC; 
  signal tx_output_N81613 : STD_LOGIC; 
  signal mac_control_CHOICE2825 : STD_LOGIC; 
  signal mac_control_CHOICE2822 : STD_LOGIC; 
  signal mac_control_CHOICE2162 : STD_LOGIC; 
  signal mac_control_CHOICE2159 : STD_LOGIC; 
  signal mac_control_N81817 : STD_LOGIC; 
  signal mac_control_N81813 : STD_LOGIC; 
  signal rx_input_ce : STD_LOGIC; 
  signal rx_input_memio_crcen : STD_LOGIC; 
  signal rx_input_memio_n0102 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd5 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd2 : STD_LOGIC; 
  signal rx_input_memio_cs_Out916_2 : STD_LOGIC; 
  signal rx_input_memio_bpen : STD_LOGIC; 
  signal rx_input_memio_n0031 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd13 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd9 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd8 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd7 : STD_LOGIC; 
  signal rx_input_memio_men : STD_LOGIC; 
  signal rx_input_memio_menl : STD_LOGIC; 
  signal rx_input_memio_n0033 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd14 : STD_LOGIC; 
  signal rx_input_memio_n0046 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd12 : STD_LOGIC; 
  signal rx_input_memio_n0047 : STD_LOGIC; 
  signal mac_control_N52268 : STD_LOGIC; 
  signal mac_control_N70611 : STD_LOGIC; 
  signal mac_control_CHOICE2889 : STD_LOGIC; 
  signal mac_control_CHOICE2886 : STD_LOGIC; 
  signal mac_control_CHOICE2662 : STD_LOGIC; 
  signal mac_control_N81757 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd4 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd2 : STD_LOGIC; 
  signal mac_control_PHY_status_n0019_2 : STD_LOGIC; 
  signal tx_output_N81605 : STD_LOGIC; 
  signal tx_output_N81609 : STD_LOGIC; 
  signal mac_control_N81753 : STD_LOGIC; 
  signal mac_control_CHOICE2223 : STD_LOGIC; 
  signal rx_output_fifo_N10 : STD_LOGIC; 
  signal rx_output_fifo_N11 : STD_LOGIC; 
  signal rx_output_fifo_N1546 : STD_LOGIC; 
  signal rx_output_fifo_N1547 : STD_LOGIC; 
  signal rx_output_fifo_N2 : STD_LOGIC; 
  signal rx_output_fifo_N1517 : STD_LOGIC; 
  signal rx_output_fifo_N3 : STD_LOGIC; 
  signal rx_output_fifo_N1610 : STD_LOGIC; 
  signal rx_output_fifo_N1611 : STD_LOGIC; 
  signal rx_output_fifo_N1563 : STD_LOGIC; 
  signal rx_output_fifo_N1562 : STD_LOGIC; 
  signal rx_output_fifo_N1551 : STD_LOGIC; 
  signal rx_output_fifo_N1550 : STD_LOGIC; 
  signal rx_output_fifo_N1567 : STD_LOGIC; 
  signal rx_output_fifo_N1566 : STD_LOGIC; 
  signal rx_output_fifo_N1627 : STD_LOGIC; 
  signal rx_output_fifo_N1626 : STD_LOGIC; 
  signal rx_output_ceinll : STD_LOGIC; 
  signal rx_output_fifo_full_0 : STD_LOGIC; 
  signal rx_output_fifo_N19 : STD_LOGIC; 
  signal rx_output_fifo_N3617 : STD_LOGIC; 
  signal rx_output_fifo_N1549 : STD_LOGIC; 
  signal rx_output_fifo_N1548 : STD_LOGIC; 
  signal rx_output_fifo_N1565 : STD_LOGIC; 
  signal rx_output_fifo_N1564 : STD_LOGIC; 
  signal rx_output_fifo_N1553 : STD_LOGIC; 
  signal rx_output_fifo_N1552 : STD_LOGIC; 
  signal rx_output_fifo_N1569 : STD_LOGIC; 
  signal rx_output_fifo_N1568 : STD_LOGIC; 
  signal rx_output_fifo_N1613 : STD_LOGIC; 
  signal rx_output_fifo_N1612 : STD_LOGIC; 
  signal rx_output_fifo_N1629 : STD_LOGIC; 
  signal rx_output_fifo_N1628 : STD_LOGIC; 
  signal rx_output_fifo_N1617 : STD_LOGIC; 
  signal rx_output_fifo_N1616 : STD_LOGIC; 
  signal rx_output_fifo_N1633 : STD_LOGIC; 
  signal rx_output_fifo_N1632 : STD_LOGIC; 
  signal rx_output_fifo_N1615 : STD_LOGIC; 
  signal rx_output_fifo_N1614 : STD_LOGIC; 
  signal rx_output_fifo_N1631 : STD_LOGIC; 
  signal rx_output_fifo_N1630 : STD_LOGIC; 
  signal rx_output_fifo_N1573 : STD_LOGIC; 
  signal rx_output_fifo_N1572 : STD_LOGIC; 
  signal rx_output_fifo_N1577 : STD_LOGIC; 
  signal rx_output_fifo_N1576 : STD_LOGIC; 
  signal mac_control_PHY_status_n0019 : STD_LOGIC; 
  signal rx_output_fifo_N1575 : STD_LOGIC; 
  signal rx_output_fifo_N1574 : STD_LOGIC; 
  signal rx_output_cs_FFd18_In_2 : STD_LOGIC; 
  signal rx_output_n0017 : STD_LOGIC; 
  signal rx_output_cs_FFd18 : STD_LOGIC; 
  signal clken3 : STD_LOGIC; 
  signal rx_output_fifo_N5 : STD_LOGIC; 
  signal rx_output_fifo_N4 : STD_LOGIC; 
  signal rx_output_fifo_N1605 : STD_LOGIC; 
  signal rx_output_fifo_N1604 : STD_LOGIC; 
  signal rx_output_fifo_N9 : STD_LOGIC; 
  signal rx_output_fifo_N8 : STD_LOGIC; 
  signal rx_output_fifo_N1609 : STD_LOGIC; 
  signal rx_output_fifo_N1608 : STD_LOGIC; 
  signal mac_control_PHY_status_n0020 : STD_LOGIC; 
  signal rx_output_fifo_N1585 : STD_LOGIC; 
  signal rx_output_fifo_N1584 : STD_LOGIC; 
  signal rx_output_fifo_N1571 : STD_LOGIC; 
  signal rx_output_fifo_N1570 : STD_LOGIC; 
  signal rx_output_fifo_N1578 : STD_LOGIC; 
  signal rx_output_fifo_N1579 : STD_LOGIC; 
  signal rx_output_fifo_N1586 : STD_LOGIC; 
  signal rx_output_fifo_N1587 : STD_LOGIC; 
  signal rx_output_fifo_N3959 : STD_LOGIC; 
  signal rx_output_fifo_N1582 : STD_LOGIC; 
  signal rx_output_fifo_N1583 : STD_LOGIC; 
  signal rx_output_fifo_N1591 : STD_LOGIC; 
  signal rx_output_fifo_N3958 : STD_LOGIC; 
  signal rx_output_fifo_N1603 : STD_LOGIC; 
  signal rx_output_fifo_N1602 : STD_LOGIC; 
  signal rx_output_fifo_N7 : STD_LOGIC; 
  signal rx_output_fifo_N6 : STD_LOGIC; 
  signal rx_output_fifo_N1607 : STD_LOGIC; 
  signal rx_output_fifo_N1606 : STD_LOGIC; 
  signal memcontroller_oe : STD_LOGIC; 
  signal rx_output_fifo_N1581 : STD_LOGIC; 
  signal rx_output_fifo_N1580 : STD_LOGIC; 
  signal clken2 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0013 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N69539 : STD_LOGIC; 
  signal tx_output_crc_10_Q : STD_LOGIC; 
  signal mac_control_CHOICE2114 : STD_LOGIC; 
  signal mac_control_CHOICE2111 : STD_LOGIC; 
  signal mac_control_CHOICE2693 : STD_LOGIC; 
  signal mac_control_N81793 : STD_LOGIC; 
  signal rx_output_lmasell : STD_LOGIC; 
  signal tx_output_bcnt_40 : STD_LOGIC; 
  signal tx_output_bcnt_38 : STD_LOGIC; 
  signal tx_output_bcnt_39 : STD_LOGIC; 
  signal tx_output_N73488 : STD_LOGIC; 
  signal tx_input_enable : STD_LOGIC; 
  signal rx_input_memio_crc_3_Q : STD_LOGIC; 
  signal mac_control_N82125 : STD_LOGIC; 
  signal mac_control_N82137 : STD_LOGIC; 
  signal tx_fifocheck_N73964 : STD_LOGIC; 
  signal mac_control_CHOICE2138 : STD_LOGIC; 
  signal mac_control_CHOICE2135 : STD_LOGIC; 
  signal mac_control_CHOICE2631 : STD_LOGIC; 
  signal mac_control_N81749 : STD_LOGIC; 
  signal tx_output_crc_11_Q : STD_LOGIC; 
  signal mac_control_CHOICE2259 : STD_LOGIC; 
  signal mac_control_CHOICE2242 : STD_LOGIC; 
  signal mac_control_N81657 : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_2 : STD_LOGIC; 
  signal tx_output_N70584 : STD_LOGIC; 
  signal rx_input_GMII_endf : STD_LOGIC; 
  signal mac_control_n00561_2 : STD_LOGIC; 
  signal mac_control_N82113 : STD_LOGIC; 
  signal tx_output_N70557 : STD_LOGIC; 
  signal tx_output_N70530 : STD_LOGIC; 
  signal tx_output_CHOICE1289 : STD_LOGIC; 
  signal tx_output_CHOICE1297 : STD_LOGIC; 
  signal tx_output_CHOICE1277 : STD_LOGIC; 
  signal tx_output_CHOICE1285 : STD_LOGIC; 
  signal tx_output_CHOICE1253 : STD_LOGIC; 
  signal tx_output_CHOICE1261 : STD_LOGIC; 
  signal tx_output_CHOICE1265 : STD_LOGIC; 
  signal tx_output_CHOICE1273 : STD_LOGIC; 
  signal mac_control_CHOICE2297 : STD_LOGIC; 
  signal mac_control_CHOICE2280 : STD_LOGIC; 
  signal mac_control_N81645 : STD_LOGIC; 
  signal tx_output_CHOICE1241 : STD_LOGIC; 
  signal tx_output_CHOICE1249 : STD_LOGIC; 
  signal tx_output_N70503 : STD_LOGIC; 
  signal tx_output_CHOICE1229 : STD_LOGIC; 
  signal tx_output_CHOICE1237 : STD_LOGIC; 
  signal tx_output_CHOICE1217 : STD_LOGIC; 
  signal tx_output_CHOICE1225 : STD_LOGIC; 
  signal tx_output_CHOICE1205 : STD_LOGIC; 
  signal tx_output_CHOICE1213 : STD_LOGIC; 
  signal tx_output_N69304 : STD_LOGIC; 
  signal tx_input_cs_FFd5 : STD_LOGIC; 
  signal tx_input_cs_FFd9 : STD_LOGIC; 
  signal tx_input_n0033 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_sout : STD_LOGIC; 
  signal SCS_IBUF : STD_LOGIC; 
  signal SIN_IBUF : STD_LOGIC; 
  signal MCLK_OBUF : STD_LOGIC; 
  signal tx_input_newframel : STD_LOGIC; 
  signal CLKIN_IBUFG : STD_LOGIC; 
  signal memcontroller_n0116 : STD_LOGIC; 
  signal RX_CLK_IBUFG : STD_LOGIC; 
  signal rx_input_GMII_rx_erl : STD_LOGIC; 
  signal memcontroller_oel : STD_LOGIC; 
  signal CLKIOIN_IBUFG : STD_LOGIC; 
  signal clkio_to_bufg : STD_LOGIC; 
  signal clk_to_bufg : STD_LOGIC; 
  signal clkrx_to_bufg : STD_LOGIC; 
  signal GLOBAL_LOGIC0 : STD_LOGIC; 
  signal rx_input_endfin : STD_LOGIC; 
  signal rx_output_fifo_N12 : STD_LOGIC; 
  signal rx_output_fifo_N13 : STD_LOGIC; 
  signal rx_output_fifo_N14 : STD_LOGIC; 
  signal rx_output_fifo_N15 : STD_LOGIC; 
  signal rx_output_fifo_N16 : STD_LOGIC; 
  signal rx_output_fifo_N17 : STD_LOGIC; 
  signal mac_control_CHOICE1813 : STD_LOGIC; 
  signal mac_control_CHOICE1869 : STD_LOGIC; 
  signal mac_control_CHOICE1841 : STD_LOGIC; 
  signal mac_control_CHOICE1897 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2588 : STD_LOGIC; 
  signal tx_output_addrinc : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_1 : STD_LOGIC; 
  signal GLOBAL_LOGIC1 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_3 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_5 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_7 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_9 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_11 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_13 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_271 : STD_LOGIC; 
  signal rx_input_memio_bcnt_86 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_273 : STD_LOGIC; 
  signal rx_input_memio_bcnt_87 : STD_LOGIC; 
  signal rx_input_memio_bcnt_88 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_275 : STD_LOGIC; 
  signal rx_input_memio_bcnt_89 : STD_LOGIC; 
  signal rx_input_memio_bcnt_90 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_277 : STD_LOGIC; 
  signal rx_input_memio_bcnt_91 : STD_LOGIC; 
  signal rx_input_memio_bcnt_92 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_279 : STD_LOGIC; 
  signal rx_input_memio_bcnt_93 : STD_LOGIC; 
  signal rx_input_memio_bcnt_94 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_281 : STD_LOGIC; 
  signal rx_input_memio_bcnt_95 : STD_LOGIC; 
  signal rx_input_memio_bcnt_96 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_283 : STD_LOGIC; 
  signal rx_input_memio_bcnt_97 : STD_LOGIC; 
  signal rx_input_memio_bcnt_98 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_285 : STD_LOGIC; 
  signal rx_input_memio_bcnt_99 : STD_LOGIC; 
  signal rx_input_memio_bcnt_100 : STD_LOGIC; 
  signal rx_input_memio_bcnt_101 : STD_LOGIC; 
  signal rx_input_memio_cs_Out916_SW0_2 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_49 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_51 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_53 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_55 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_57 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_59 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_61 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_222 : STD_LOGIC; 
  signal rx_input_memio_macnt_70 : STD_LOGIC; 
  signal rx_input_memio_macnt_71 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_224 : STD_LOGIC; 
  signal rx_input_memio_macnt_72 : STD_LOGIC; 
  signal rx_input_memio_macnt_73 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_226 : STD_LOGIC; 
  signal rx_input_memio_macnt_74 : STD_LOGIC; 
  signal rx_input_memio_macnt_75 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_228 : STD_LOGIC; 
  signal rx_input_memio_macnt_76 : STD_LOGIC; 
  signal rx_input_memio_macnt_77 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_230 : STD_LOGIC; 
  signal rx_input_memio_macnt_78 : STD_LOGIC; 
  signal rx_input_memio_macnt_79 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_232 : STD_LOGIC; 
  signal rx_input_memio_macnt_80 : STD_LOGIC; 
  signal rx_input_memio_macnt_81 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_234 : STD_LOGIC; 
  signal rx_input_memio_macnt_82 : STD_LOGIC; 
  signal rx_input_memio_macnt_83 : STD_LOGIC; 
  signal rx_input_memio_macnt_84 : STD_LOGIC; 
  signal rx_input_memio_macnt_85 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_341 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_343 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_345 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_347 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_349 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_351 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_195 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_197 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_199 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_201 : STD_LOGIC; 
  signal tx_output_n0035 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_87 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_89 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_91 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_93 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_95 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_97 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_99 : STD_LOGIC; 
  signal tx_output_n0033 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_205 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_207 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_209 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_211 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_213 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_215 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_217 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_219 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_79 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_81 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_83 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_162 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_164 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_166 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_168 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_170 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_172 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_174 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_162 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_164 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_166 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_168 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_170 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_172 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_174 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_328 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_330 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_332 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_334 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_336 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_338 : STD_LOGIC; 
  signal rx_output_fifo_N1919 : STD_LOGIC; 
  signal rx_output_fifo_N1929 : STD_LOGIC; 
  signal rx_output_fifo_N1939 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_119 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_121 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_123 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_125 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_127 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_129 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_131 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_188 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_190 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_192 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_36 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_79 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_81 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_83 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_102 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_104 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_106 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_108 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_110 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_112 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_114 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_116 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_152 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_154 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_156 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_158 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_152 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_154 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_156 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_158 : STD_LOGIC; 
  signal tx_fifocheck_n0003 : STD_LOGIC; 
  signal mac_control_N80441 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_295 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_297 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_299 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_301 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_303 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_305 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_307 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_309 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_311 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_313 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_315 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_317 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_319 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_321 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_323 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_325 : STD_LOGIC; 
  signal rx_input_memio_n0101 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_254 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_256 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_258 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_260 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_262 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_264 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_266 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_268 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_64 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_66 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_68 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_70 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_72 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_74 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_76 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_79 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_81 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_83 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_238 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_240 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_242 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_244 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_246 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_248 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_250 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_135 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_137 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_139 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_141 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_143 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_145 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_147 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_149 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_182 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_184 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178 : STD_LOGIC; 
  signal rx_output_fifo_N2847 : STD_LOGIC; 
  signal rx_output_fifo_N2857 : STD_LOGIC; 
  signal rx_output_fifo_N2867 : STD_LOGIC; 
  signal rx_output_fifo_N2576 : STD_LOGIC; 
  signal rx_output_fifo_N2574 : STD_LOGIC; 
  signal rx_output_fifo_N2572 : STD_LOGIC; 
  signal rx_output_fifo_BU172_O : STD_LOGIC; 
  signal rx_output_fifo_N3614 : STD_LOGIC; 
  signal rx_output_fifo_N3612 : STD_LOGIC; 
  signal rx_output_fifo_N3610 : STD_LOGIC; 
  signal rx_output_fifo_BU351_O : STD_LOGIC; 
  signal rx_output_fifo_N4763 : STD_LOGIC; 
  signal rx_output_fifo_N1593 : STD_LOGIC; 
  signal rx_output_fifo_N1592 : STD_LOGIC; 
  signal rx_output_fifo_N4771 : STD_LOGIC; 
  signal rx_output_fifo_N1590 : STD_LOGIC; 
  signal rx_output_fifo_N4779 : STD_LOGIC; 
  signal rx_output_fifo_N1589 : STD_LOGIC; 
  signal rx_output_fifo_N1588 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_288 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_290 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd11 : STD_LOGIC; 
  signal rx_input_memio_wbpl : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd6 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd8 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd6 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd3 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1570 : STD_LOGIC; 
  signal tx_input_enableint : STD_LOGIC; 
  signal tx_input_enableintl : STD_LOGIC; 
  signal mac_control_PHY_status_done : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd5 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd7 : STD_LOGIC; 
  signal tx_output_decbcnt : STD_LOGIC; 
  signal rxfifowerr : STD_LOGIC; 
  signal rxcrcerr : STD_LOGIC; 
  signal rxphyerr : STD_LOGIC; 
  signal tx_input_newfint : STD_LOGIC; 
  signal tx_input_cs_FFd8 : STD_LOGIC; 
  signal mac_control_PHY_status_n0017 : STD_LOGIC; 
  signal mac_control_PHY_status_n0018 : STD_LOGIC; 
  signal mac_control_CHOICE2197 : STD_LOGIC; 
  signal mac_control_CHOICE2423 : STD_LOGIC; 
  signal mac_control_CHOICE2277 : STD_LOGIC; 
  signal mac_control_CHOICE2429 : STD_LOGIC; 
  signal mac_control_CHOICE2021 : STD_LOGIC; 
  signal mac_control_CHOICE2874 : STD_LOGIC; 
  signal mac_control_CHOICE2859 : STD_LOGIC; 
  signal mac_control_CHOICE2420 : STD_LOGIC; 
  signal mac_control_CHOICE2431 : STD_LOGIC; 
  signal mac_control_CHOICE2665 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_12_94_1 : STD_LOGIC; 
  signal mac_control_CHOICE2872 : STD_LOGIC; 
  signal mac_control_CHOICE2869 : STD_LOGIC; 
  signal mac_control_N81769 : STD_LOGIC; 
  signal mac_control_CHOICE1939 : STD_LOGIC; 
  signal mac_control_CHOICE1942 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_20_66_1 : STD_LOGIC; 
  signal mac_control_CHOICE2322 : STD_LOGIC; 
  signal mac_control_CHOICE2366 : STD_LOGIC; 
  signal mac_control_CHOICE2676 : STD_LOGIC; 
  signal mac_control_CHOICE2668 : STD_LOGIC; 
  signal mac_control_CHOICE2673 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_12_94_SW0_2 : STD_LOGIC; 
  signal mac_control_CHOICE2833 : STD_LOGIC; 
  signal mac_control_CHOICE2865 : STD_LOGIC; 
  signal mac_control_CHOICE2606 : STD_LOGIC; 
  signal mac_control_CHOICE2290 : STD_LOGIC; 
  signal mac_control_CHOICE1952 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_20_42_1 : STD_LOGIC; 
  signal mac_control_CHOICE1949 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_20_77_1 : STD_LOGIC; 
  signal mac_control_CHOICE1954 : STD_LOGIC; 
  signal mac_control_CHOICE2148 : STD_LOGIC; 
  signal mac_control_CHOICE2151 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_21_69_1 : STD_LOGIC; 
  signal mac_control_CHOICE2696 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_13_94_1 : STD_LOGIC; 
  signal mac_control_CHOICE2124 : STD_LOGIC; 
  signal mac_control_CHOICE2018 : STD_LOGIC; 
  signal mac_control_CHOICE2680 : STD_LOGIC; 
  signal mac_control_CHOICE2683 : STD_LOGIC; 
  signal mac_control_CHOICE2684 : STD_LOGIC; 
  signal mac_control_CHOICE2707 : STD_LOGIC; 
  signal mac_control_CHOICE2699 : STD_LOGIC; 
  signal mac_control_CHOICE2704 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_13_94_SW0_2 : STD_LOGIC; 
  signal mac_control_CHOICE2618 : STD_LOGIC; 
  signal mac_control_CHOICE2637 : STD_LOGIC; 
  signal mac_control_CHOICE2385 : STD_LOGIC; 
  signal mac_control_CHOICE2461 : STD_LOGIC; 
  signal mac_control_CHOICE2057 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_30_66_1 : STD_LOGIC; 
  signal mac_control_CHOICE1962 : STD_LOGIC; 
  signal mac_control_CHOICE1965 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_22_66_1 : STD_LOGIC; 
  signal mac_control_CHOICE2614 : STD_LOGIC; 
  signal mac_control_CHOICE2687 : STD_LOGIC; 
  signal mac_control_CHOICE2714 : STD_LOGIC; 
  signal mac_control_CHOICE2715 : STD_LOGIC; 
  signal mac_control_N52081 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_21_80_1 : STD_LOGIC; 
  signal mac_control_CHOICE2164 : STD_LOGIC; 
  signal mac_control_CHOICE2391 : STD_LOGIC; 
  signal mac_control_CHOICE2467 : STD_LOGIC; 
  signal mac_control_CHOICE2067 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_30_42_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_30_77_1 : STD_LOGIC; 
  signal mac_control_CHOICE2069 : STD_LOGIC; 
  signal mac_control_CHOICE1929 : STD_LOGIC; 
  signal mac_control_CHOICE1975 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_22_42_1 : STD_LOGIC; 
  signal mac_control_CHOICE1972 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_22_77_1 : STD_LOGIC; 
  signal mac_control_CHOICE1977 : STD_LOGIC; 
  signal mac_control_CHOICE1998 : STD_LOGIC; 
  signal mac_control_CHOICE2044 : STD_LOGIC; 
  signal mac_control_CHOICE1926 : STD_LOGIC; 
  signal mac_control_CHOICE2906 : STD_LOGIC; 
  signal mac_control_CHOICE2891 : STD_LOGIC; 
  signal mac_control_CHOICE2718 : STD_LOGIC; 
  signal mac_control_CHOICE2458 : STD_LOGIC; 
  signal mac_control_CHOICE2469 : STD_LOGIC; 
  signal mac_control_CHOICE1995 : STD_LOGIC; 
  signal mac_control_CHOICE2216 : STD_LOGIC; 
  signal mac_control_CHOICE2210 : STD_LOGIC; 
  signal mac_control_CHOICE2206 : STD_LOGIC; 
  signal mac_control_CHOICE2224 : STD_LOGIC; 
  signal mac_control_CHOICE1802 : STD_LOGIC; 
  signal mac_control_CHOICE1805 : STD_LOGIC; 
  signal mac_control_CHOICE2309 : STD_LOGIC; 
  signal mac_control_CHOICE2100 : STD_LOGIC; 
  signal mac_control_CHOICE2103 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_16_69_1 : STD_LOGIC; 
  signal mac_control_CHOICE1858 : STD_LOGIC; 
  signal mac_control_CHOICE1861 : STD_LOGIC; 
  signal mac_control_CHOICE2233 : STD_LOGIC; 
  signal mac_control_CHOICE2904 : STD_LOGIC; 
  signal mac_control_CHOICE2901 : STD_LOGIC; 
  signal mac_control_N81745 : STD_LOGIC; 
  signal mac_control_CHOICE2172 : STD_LOGIC; 
  signal mac_control_CHOICE2175 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_24_69_1 : STD_LOGIC; 
  signal mac_control_CHOICE2347 : STD_LOGIC; 
  signal mac_control_CHOICE2649 : STD_LOGIC; 
  signal mac_control_CHOICE2897 : STD_LOGIC; 
  signal mac_control_CHOICE1833 : STD_LOGIC; 
  signal mac_control_CHOICE1830 : STD_LOGIC; 
  signal mac_control_CHOICE2404 : STD_LOGIC; 
  signal mac_control_CHOICE2077 : STD_LOGIC; 
  signal tx_output_crc_13_Q : STD_LOGIC; 
  signal mac_control_CHOICE2127 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_17_69_1 : STD_LOGIC; 
  signal mac_control_CHOICE1985 : STD_LOGIC; 
  signal mac_control_CHOICE1988 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_25_66_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_16_80_1 : STD_LOGIC; 
  signal mac_control_CHOICE2116 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_24_80_1 : STD_LOGIC; 
  signal mac_control_CHOICE2188 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_25_42_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_25_77_1 : STD_LOGIC; 
  signal mac_control_CHOICE2000 : STD_LOGIC; 
  signal mac_control_CHOICE2252 : STD_LOGIC; 
  signal mac_control_CHOICE2246 : STD_LOGIC; 
  signal mac_control_CHOICE2258 : STD_LOGIC; 
  signal mac_control_CHOICE2008 : STD_LOGIC; 
  signal mac_control_CHOICE2011 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_26_66_1 : STD_LOGIC; 
  signal mac_control_CHOICE1916 : STD_LOGIC; 
  signal mac_control_CHOICE1919 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_18_66_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_17_80_1 : STD_LOGIC; 
  signal mac_control_CHOICE2140 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_18_42_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_18_77_1 : STD_LOGIC; 
  signal mac_control_CHOICE1931 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_26_42_1 : STD_LOGIC; 
  signal mac_control_CHOICE2023 : STD_LOGIC; 
  signal mac_control_CHOICE2284 : STD_LOGIC; 
  signal mac_control_CHOICE2296 : STD_LOGIC; 
  signal mac_control_CHOICE1886 : STD_LOGIC; 
  signal mac_control_CHOICE1889 : STD_LOGIC; 
  signal mac_control_CHOICE2031 : STD_LOGIC; 
  signal mac_control_CHOICE2034 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_28_66_1 : STD_LOGIC; 
  signal mac_control_CHOICE2360 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_28_42_1 : STD_LOGIC; 
  signal mac_control_CHOICE2041 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_28_77_1 : STD_LOGIC; 
  signal mac_control_CHOICE2046 : STD_LOGIC; 
  signal mac_control_CHOICE2080 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_29_66_1 : STD_LOGIC; 
  signal mac_control_CHOICE2087 : STD_LOGIC; 
  signal mac_control_CHOICE2090 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_29_42_1 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_29_77_1 : STD_LOGIC; 
  signal mac_control_CHOICE2092 : STD_LOGIC; 
  signal mac_control_CHOICE2372 : STD_LOGIC; 
  signal mac_control_CHOICE2373 : STD_LOGIC; 
  signal rx_input_memio_crc_6_Q : STD_LOGIC; 
  signal mac_control_CHOICE2328 : STD_LOGIC; 
  signal mac_control_CHOICE2334 : STD_LOGIC; 
  signal mac_control_CHOICE2335 : STD_LOGIC; 
  signal mac_control_CHOICE2398 : STD_LOGIC; 
  signal mac_control_CHOICE2410 : STD_LOGIC; 
  signal mac_control_CHOICE2411 : STD_LOGIC; 
  signal tx_input_CHOICE1695 : STD_LOGIC; 
  signal tx_input_CHOICE1702 : STD_LOGIC; 
  signal slowclock_rxphyerrl : STD_LOGIC; 
  signal rx_input_memio_crc_7_Q : STD_LOGIC; 
  signal rx_input_memio_cs_FFd4 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd6 : STD_LOGIC; 
  signal tx_output_crc_15_Q : STD_LOGIC; 
  signal mac_control_CHOICE2356 : STD_LOGIC; 
  signal mac_control_N81649 : STD_LOGIC; 
  signal rx_input_memio_crc_10_Q : STD_LOGIC; 
  signal rx_input_memio_crc_8_Q : STD_LOGIC; 
  signal mac_control_CHOICE2382 : STD_LOGIC; 
  signal mac_control_CHOICE2194 : STD_LOGIC; 
  signal mac_control_CHOICE2230 : STD_LOGIC; 
  signal mac_control_CHOICE2306 : STD_LOGIC; 
  signal mac_control_CHOICE2268 : STD_LOGIC; 
  signal mac_control_CHOICE2344 : STD_LOGIC; 
  signal tx_output_crc_24_Q : STD_LOGIC; 
  signal tx_output_crc_16_Q : STD_LOGIC; 
  signal mac_control_CHOICE2318 : STD_LOGIC; 
  signal mac_control_N81661 : STD_LOGIC; 
  signal rx_input_memio_crc_11_Q : STD_LOGIC; 
  signal mac_control_n0238 : STD_LOGIC; 
  signal rx_input_memio_crc_9_Q : STD_LOGIC; 
  signal rx_output_cs_FFd10_In11_1 : STD_LOGIC; 
  signal tx_output_crc_17_Q : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxbcastl : STD_LOGIC; 
  signal rx_input_memio_addrchk_validmcast : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxmcastl : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxallfl : STD_LOGIC; 
  signal rx_input_memio_addrchk_N70965 : STD_LOGIC; 
  signal rx_input_memio_destok : STD_LOGIC; 
  signal mac_control_n0033102_SW0_2 : STD_LOGIC; 
  signal mac_control_N81729 : STD_LOGIC; 
  signal rx_output_CHOICE1560 : STD_LOGIC; 
  signal tx_output_crc_26_Q : STD_LOGIC; 
  signal mac_control_lrxallf : STD_LOGIC; 
  signal mac_control_CHOICE2394 : STD_LOGIC; 
  signal mac_control_N81653 : STD_LOGIC; 
  signal rx_input_memio_crc_13_Q : STD_LOGIC; 
  signal mac_control_CHOICE2315 : STD_LOGIC; 
  signal mac_control_CHOICE2203 : STD_LOGIC; 
  signal mac_control_CHOICE2840 : STD_LOGIC; 
  signal mac_control_CHOICE2205 : STD_LOGIC; 
  signal mac_control_CHOICE2239 : STD_LOGIC; 
  signal mac_control_CHOICE2241 : STD_LOGIC; 
  signal mac_control_N81741 : STD_LOGIC; 
  signal mac_control_CHOICE2795 : STD_LOGIC; 
  signal mac_control_CHOICE2271 : STD_LOGIC; 
  signal mac_control_CHOICE2279 : STD_LOGIC; 
  signal mac_control_CHOICE2603 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_4_94_1 : STD_LOGIC; 
  signal mac_control_CHOICE2808 : STD_LOGIC; 
  signal mac_control_CHOICE2805 : STD_LOGIC; 
  signal mac_control_CHOICE2611 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_4_94_SW0_2 : STD_LOGIC; 
  signal mac_control_CHOICE2621 : STD_LOGIC; 
  signal mac_control_CHOICE2622 : STD_LOGIC; 
  signal mac_control_CHOICE2353 : STD_LOGIC; 
  signal mac_control_CHOICE2625 : STD_LOGIC; 
  signal mac_control_CHOICE2355 : STD_LOGIC; 
  signal mac_control_CHOICE2842 : STD_LOGIC; 
  signal mac_control_CHOICE2827 : STD_LOGIC; 
  signal mac_control_CHOICE2317 : STD_LOGIC; 
  signal mac_control_CHOICE2837 : STD_LOGIC; 
  signal mac_control_N81809 : STD_LOGIC; 
  signal mac_control_CHOICE2634 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_9_94_1 : STD_LOGIC; 
  signal mac_control_CHOICE2393 : STD_LOGIC; 
  signal mac_control_CHOICE2642 : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_9_94_SW0_2 : STD_LOGIC; 
  signal mac_control_CHOICE2652 : STD_LOGIC; 
  signal mac_control_CHOICE2653 : STD_LOGIC; 
  signal mac_control_CHOICE2656 : STD_LOGIC; 
  signal tx_output_crc_27_Q : STD_LOGIC; 
  signal tx_input_N69386 : STD_LOGIC; 
  signal tx_output_crc_28_Q : STD_LOGIC; 
  signal rx_input_memio_crc_15_Q : STD_LOGIC; 
  signal rxallf : STD_LOGIC; 
  signal tx_output_crc_29_Q : STD_LOGIC; 
  signal rx_input_memio_crc_24_Q : STD_LOGIC; 
  signal rx_input_memio_crc_16_Q : STD_LOGIC; 
  signal mac_control_n0028 : STD_LOGIC; 
  signal mac_control_n0026 : STD_LOGIC; 
  signal mac_control_n0027 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd3_In_1 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2593 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2564 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2574 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2575 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd4_In_2 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2591 : STD_LOGIC; 
  signal tx_output_N69282 : STD_LOGIC; 
  signal tx_input_CHOICE1722 : STD_LOGIC; 
  signal tx_output_N70823 : STD_LOGIC; 
  signal rx_input_memio_crc_17_Q : STD_LOGIC; 
  signal mac_control_PHY_status_n0019_SW0_2 : STD_LOGIC; 
  signal tx_input_CHOICE1725 : STD_LOGIC; 
  signal mac_control_PHY_status_start : STD_LOGIC; 
  signal rx_input_memio_crc_26_Q : STD_LOGIC; 
  signal rx_input_fifo_control_celll : STD_LOGIC; 
  signal rx_input_memio_crc_27_Q : STD_LOGIC; 
  signal mac_control_PHY_status_N41765 : STD_LOGIC; 
  signal rx_input_fifo_control_cell : STD_LOGIC; 
  signal rx_input_memio_crc_28_Q : STD_LOGIC; 
  signal mac_control_PHY_status_N41773 : STD_LOGIC; 
  signal rx_input_memio_crccomb_N82101 : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1742 : STD_LOGIC; 
  signal rx_input_memio_crc_29_Q : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1749 : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1764 : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1757 : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1765 : STD_LOGIC; 
  signal rx_input_memio_cs_Out8_2 : STD_LOGIC; 
  signal rx_output_N70216 : STD_LOGIC; 
  signal rx_output_N70268 : STD_LOGIC; 
  signal rx_output_N70320 : STD_LOGIC; 
  signal rx_output_N69748 : STD_LOGIC; 
  signal mac_control_CHOICE2986 : STD_LOGIC; 
  signal rx_output_N70372 : STD_LOGIC; 
  signal rx_output_N69696 : STD_LOGIC; 
  signal tx_output_crc_loigc_N81880 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_0 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_1 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_2 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_3 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_4 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_5 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_6 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_7 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_8 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_9 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_10 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_11 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_12 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_13 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_14 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_15 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_16 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_17 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_18 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_19 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_20 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_21 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_22 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_23 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_24 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_25 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_26 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_27 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_28 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_29 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_30 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_31 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_32 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_33 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_34 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_35 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_36 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_37 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_0 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_1 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_2 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_3 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_4 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_5 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_6 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_7 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_8 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_9 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_10 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_11 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_12 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_13 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_14 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_15 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_16 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_17 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_18 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_19 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_20 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_21 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_22 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_23 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_24 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_25 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_26 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_27 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_28 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_29 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_30 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_31 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_32 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_33 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_34 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_35 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_36 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_37 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_38 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_39 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_40 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_41 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_42 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_43 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_44 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_45 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_46 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_47 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_48 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_49 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_50 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_51 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_52 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_53 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_54 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_55 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_56 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_57 : STD_LOGIC; 
  signal GSR : STD_LOGIC; 
  signal GTS : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5329_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2364_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2364_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_full_FFX_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_full_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4913 : STD_LOGIC; 
  signal rx_input_fifo_fifo_full_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2427_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4892 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2427_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4891 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4902 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2427_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2427_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2478_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2478_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4690 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4730 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3985 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3943 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3990 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3987 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3944 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2417_FFX_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2417_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2428_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4894 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2428_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4893 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4904 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2428_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2428_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2438_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2467_FFY_SET : STD_LOGIC; 
  signal rx_input_rx_nearf_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6356 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6362 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6359 : STD_LOGIC; 
  signal rx_input_rx_nearf_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6323 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5349 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4610 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4650 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3975 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3941 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3980 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3977 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3942 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4896 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2431_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4895 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4906 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2431_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2431_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2469_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6348 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6355_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6352 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6351 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6355_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5348 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2449_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2428_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4530 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4570 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3965 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3939 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N7_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3970 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3967 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N7_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3940 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4898 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2432_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4897 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4908 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2432_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2432_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6340 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6347_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6344 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6343 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6347_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5346 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5345 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4490 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4450 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3955 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3937 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N9_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3960 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3957 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N9_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3938 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4900 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2434_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4899 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4910 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2434_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2434_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2443_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6332 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6339_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6336 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6335 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6339_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2438_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5344 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5343 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4370 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4410 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3945 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3935 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3950 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3947 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3936 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2436_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2475_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6324 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6331_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6328 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6327 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6331_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5342 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5341 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2467_FFX_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2362_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2362_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2447_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2724 : STD_LOGIC; 
  signal rx_input_fifo_fifo_empty_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3647 : STD_LOGIC; 
  signal rx_input_fifo_fifo_empty_CYINIT : STD_LOGIC; 
  signal mac_control_lmacaddr_27_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_37_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_45_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_29_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_39_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_47_FFY_RST : STD_LOGIC; 
  signal rxbp_11_FFY_RST : STD_LOGIC; 
  signal rxbp_11_CEMUXNOT : STD_LOGIC; 
  signal rxbp_13_FFY_RST : STD_LOGIC; 
  signal rxbp_13_CEMUXNOT : STD_LOGIC; 
  signal rxbp_15_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifo_N2579_FROM : STD_LOGIC; 
  signal rx_output_fifo_N2579_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1835 : STD_LOGIC; 
  signal rx_output_invalid_GROM : STD_LOGIC; 
  signal q2_1_FFY_RST : STD_LOGIC; 
  signal mac_control_Ker52136_2_GROM : STD_LOGIC; 
  signal q3_1_FFY_RST : STD_LOGIC; 
  signal q2_7_FFY_RST : STD_LOGIC; 
  signal q3_3_FFY_RST : STD_LOGIC; 
  signal q2_9_FFY_RST : STD_LOGIC; 
  signal q3_5_FFY_RST : STD_LOGIC; 
  signal rxfbbp_11_FFY_RST : STD_LOGIC; 
  signal rxfbbp_11_CEMUXNOT : STD_LOGIC; 
  signal q3_7_FFY_RST : STD_LOGIC; 
  signal rxfbbp_13_FFY_RST : STD_LOGIC; 
  signal rxfbbp_13_CEMUXNOT : STD_LOGIC; 
  signal q3_9_FFY_RST : STD_LOGIC; 
  signal rxfbbp_15_FFY_RST : STD_LOGIC; 
  signal rxfbbp_15_CEMUXNOT : STD_LOGIC; 
  signal rxfifowerrsr_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_11_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_11_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_13_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_13_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_15_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_15_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5_FFX_RST : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2_GROM : STD_LOGIC; 
  signal tx_output_outsell_2_FFY_RST : STD_LOGIC; 
  signal tx_output_outsell_2_FROM : STD_LOGIC; 
  signal tx_output_outsel_3_Q : STD_LOGIC; 
  signal tx_output_outsell_2_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2420_FFY_RST : STD_LOGIC; 
  signal slowclock_txfifowerrl_LOGIC_ZERO : STD_LOGIC; 
  signal slowclock_txfifowerrl_GROM : STD_LOGIC; 
  signal rx_input_memio_fifofulll_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_fifofulll_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_endbyte_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_endbyte_2_FFY_RST : STD_LOGIC; 
  signal rx_output_nfl_FFY_RST : STD_LOGIC; 
  signal rx_output_nfl_CEMUXNOT : STD_LOGIC; 
  signal mac_control_addr_1_FFY_RST : STD_LOGIC; 
  signal mac_control_addr_3_FFY_RST : STD_LOGIC; 
  signal mac_control_addr_5_FFY_RST : STD_LOGIC; 
  signal mac_control_addr_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2431_FFY_RST : STD_LOGIC; 
  signal tx_input_CHOICE1710_FROM : STD_LOGIC; 
  signal tx_input_CHOICE1710_GROM : STD_LOGIC; 
  signal tx_input_CHOICE1717_FROM : STD_LOGIC; 
  signal tx_input_CHOICE1717_GROM : STD_LOGIC; 
  signal tx_input_cs_FFd10_FROM : STD_LOGIC; 
  signal tx_input_cs_FFd10_In : STD_LOGIC; 
  signal mac_control_din_11_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3626 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2497_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3625 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3636 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2497_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2497_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3600 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3560 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2855 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2813 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2860 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2857 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N13_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2814 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3628 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2499_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3627 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3638 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2499_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2499_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3480 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3520 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2845 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2811 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2850 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2847 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2812 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3630 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2500_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3629 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3640 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2500_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2500_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3440 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3400 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2835 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2809 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N17_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2840 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2837 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N17_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2810 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3632 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2502_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3631 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3642 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2502_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2502_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3320 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3360 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2825 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2807 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N19_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2830 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2827 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N19_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2808 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3634 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2504_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3633 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3644 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2504_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2504_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3240 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3280 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2815 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2805 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N21_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2820 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2817 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N21_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N21_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2806 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2505_GROM : STD_LOGIC; 
  signal slowclock_n0002_FROM : STD_LOGIC; 
  signal slowclock_n0002_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_9_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dh_13_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_15_FFY_RST : STD_LOGIC; 
  signal mac_control_N81797_FROM : STD_LOGIC; 
  signal mac_control_N81797_GROM : STD_LOGIC; 
  signal rx_input_GMII_lince : STD_LOGIC; 
  signal rx_input_ince_GROM : STD_LOGIC; 
  signal txbp_11_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_13_FFY_RST : STD_LOGIC; 
  signal txbp_13_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2447_FFX_SET : STD_LOGIC; 
  signal txbp_15_FFY_RST : STD_LOGIC; 
  signal mac_control_N81777_FROM : STD_LOGIC; 
  signal mac_control_N81777_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd1_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd1_In : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxucastl_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2480_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_11_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_21_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_13_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_23_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_31_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_15_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_33_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_41_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_17_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_25_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_35_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2480_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_43_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_19_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1797_FROM : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1797_GROM : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1789_GROM : STD_LOGIC; 
  signal tx_output_cs_Out1160_SW0_1_FROM : STD_LOGIC; 
  signal tx_output_cs_Out1160_SW0_1_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1679_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1679_GROM : STD_LOGIC; 
  signal tx_output_N81625_FROM : STD_LOGIC; 
  signal tx_output_N81625_GROM : STD_LOGIC; 
  signal tx_output_crcl_5_GROM : STD_LOGIC; 
  signal tx_output_crcl_4_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_n0007_Xo_0_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_n0007_Xo_0_GROM : STD_LOGIC; 
  signal tx_output_outsell_0_FROM : STD_LOGIC; 
  signal tx_output_outsel_0_Q : STD_LOGIC; 
  signal tx_output_outsell_0_CEMUXNOT : STD_LOGIC; 
  signal mac_control_N81689_FROM : STD_LOGIC; 
  signal mac_control_N81689_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1447_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1451_GROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE2917_FROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE2917_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE2922_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE2926_GROM : STD_LOGIC; 
  signal slowclock_lclken_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_CHOICE2934_FROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE2934_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_CHOICE2941_GROM : STD_LOGIC; 
  signal mac_control_n001220_1_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_0_FROM : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_3_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_5_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_7_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_11_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_13_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_15_FFY_RST : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_29_42_SW0_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_29_42_SW0_1_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2434_FFY_RST : STD_LOGIC; 
  signal tx_output_ltxen3_FROM : STD_LOGIC; 
  signal tx_output_ltxen : STD_LOGIC; 
  signal tx_output_ltxen3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_n0030_FROM : STD_LOGIC; 
  signal mac_control_n0030_GROM : STD_LOGIC; 
  signal mac_control_n0103_FROM : STD_LOGIC; 
  signal mac_control_n0103_GROM : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_191 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_256 : STD_LOGIC; 
  signal mac_control_bitcnt_109_GROM : STD_LOGIC; 
  signal mac_control_bitcnt_109_CYINIT : STD_LOGIC; 
  signal mac_control_n0050_GROM : STD_LOGIC; 
  signal mac_control_n0042_GROM : STD_LOGIC; 
  signal mac_control_n0051_GROM : STD_LOGIC; 
  signal mac_control_n0043_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2423_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE2959_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2959_GROM : STD_LOGIC; 
  signal mac_control_n0052_GROM : STD_LOGIC; 
  signal mac_control_n0060_FROM : STD_LOGIC; 
  signal mac_control_n0060_GROM : STD_LOGIC; 
  signal mac_control_din_15_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2420_FFX_RST : STD_LOGIC; 
  signal mac_control_din_31_FFY_RST : STD_LOGIC; 
  signal mac_control_din_17_FFY_RST : STD_LOGIC; 
  signal mac_control_din_19_FFY_RST : STD_LOGIC; 
  signal mac_control_din_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crccomb_n0118_0_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_n0118_0_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n001124_2_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2439_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81705_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81705_GROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd15_FROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd15_In : STD_LOGIC; 
  signal tx_output_crcl_3_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2439_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_n00151_1_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_dout_3_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_5_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_7_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_9_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N82067_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N82067_GROM : STD_LOGIC; 
  signal rx_input_memio_bpl_13_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_FROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_In : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2431_FFX_RST : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_18_42_SW0_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_18_42_SW0_1_GROM : STD_LOGIC; 
  signal rx_input_fifo_RESET_1_GROM : STD_LOGIC; 
  signal rxf_CEMUXNOT : STD_LOGIC; 
  signal mac_control_phyaddr_3_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_5_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_7_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_9_FFY_RST : STD_LOGIC; 
  signal slowclock_rxoferrl_LOGIC_ZERO : STD_LOGIC; 
  signal slowclock_rxoferrl_GROM : STD_LOGIC; 
  signal rx_input_memio_crcrst_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_dout_1_FFY_RST : STD_LOGIC; 
  signal txfbbp_11_FFY_RST : STD_LOGIC; 
  signal txfbbp_11_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_dout_3_FFY_RST : STD_LOGIC; 
  signal txfbbp_13_FFY_RST : STD_LOGIC; 
  signal txfbbp_13_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_15_FFY_RST : STD_LOGIC; 
  signal txfbbp_15_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_dout_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_9_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N37245_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N37245_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N37240_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N37240_GROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2_GROM : STD_LOGIC; 
  signal txf_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1462_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1462_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2469_FFX_SET : STD_LOGIC; 
  signal rx_input_data_0_FROM : STD_LOGIC; 
  signal rx_output_cs_FFd9_FROM : STD_LOGIC; 
  signal rx_output_cs_FFd9_In : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1483_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1483_GROM : STD_LOGIC; 
  signal rx_input_data_1_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1656_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1490_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1490_GROM : STD_LOGIC; 
  signal rx_input_data_2_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1671_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1671_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4_In_2_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4_In_2_GROM : STD_LOGIC; 
  signal rx_input_data_3_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1664_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1476_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1476_GROM : STD_LOGIC; 
  signal rx_input_data_4_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2449_FFY_SET : STD_LOGIC; 
  signal rx_input_data_5_FROM : STD_LOGIC; 
  signal rx_input_data_6_FROM : STD_LOGIC; 
  signal rx_input_data_7_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1469_GROM : STD_LOGIC; 
  signal rx_input_endf_FROM : STD_LOGIC; 
  signal rx_input_invalid_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81600_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81600_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd2_In : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd2_GROM : STD_LOGIC; 
  signal tx_output_crcl_6_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd6_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd6_In : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_7_Xo_1_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_7_Xo_1_GROM : STD_LOGIC; 
  signal mac_control_N52153_FROM : STD_LOGIC; 
  signal mac_control_N52153_GROM : STD_LOGIC; 
  signal mac_control_N52138_FROM : STD_LOGIC; 
  signal mac_control_N52138_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd2_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd2_In : STD_LOGIC; 
  signal rx_input_fifo_fifo_N7_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_1_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2482_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2449_FFX_SET : STD_LOGIC; 
  signal macaddr_3_FFY_RST : STD_LOGIC; 
  signal macaddr_5_FFY_RST : STD_LOGIC; 
  signal macaddr_7_FFY_RST : STD_LOGIC; 
  signal macaddr_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_2_GROM : STD_LOGIC; 
  signal tx_input_N34493_FROM : STD_LOGIC; 
  signal tx_input_N34493_GROM : STD_LOGIC; 
  signal rx_output_N69253_FROM : STD_LOGIC; 
  signal rx_output_N69253_GROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0122_1_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0122_1_GROM : STD_LOGIC; 
  signal tx_output_crcl_7_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_din_3_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_5_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2432_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_9_FFY_RST : STD_LOGIC; 
  signal mac_control_N82133_FROM : STD_LOGIC; 
  signal mac_control_N82133_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2482_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2_GROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_25_42_SW0_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_25_42_SW0_1_GROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_28_42_SW0_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_28_42_SW0_1_GROM : STD_LOGIC; 
  signal tx_input_fifofulll_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_8_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_8_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2421_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_CHOICE2946_GROM : STD_LOGIC; 
  signal rx_input_memio_crcequal_FROM : STD_LOGIC; 
  signal rx_input_memio_N80267 : STD_LOGIC; 
  signal rx_input_memio_crcequal_CEMUXNOT : STD_LOGIC; 
  signal mac_control_dout_10_FROM : STD_LOGIC; 
  signal mac_control_N77583 : STD_LOGIC; 
  signal mac_control_PHY_status_phyaddrws_BYMUXNOT : STD_LOGIC; 
  signal mac_control_N82019_FROM : STD_LOGIC; 
  signal mac_control_N82019_GROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_26_Xo_1_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_26_Xo_1_GROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2_GROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0122_0_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0122_0_GROM : STD_LOGIC; 
  signal rx_output_fifo_nearfull_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_9_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_9_FROM : STD_LOGIC; 
  signal addr4ext_3_FFY_RST : STD_LOGIC; 
  signal addr4ext_5_FFY_RST : STD_LOGIC; 
  signal addr4ext_7_FFY_RST : STD_LOGIC; 
  signal addr4ext_9_FFY_RST : STD_LOGIC; 
  signal d4_3_FFY_RST : STD_LOGIC; 
  signal d4_5_FFY_RST : STD_LOGIC; 
  signal d4_7_FFY_RST : STD_LOGIC; 
  signal d4_9_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_11_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_13_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_15_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd12_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd14_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd16_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N7_FFX_RST : STD_LOGIC; 
  signal rx_output_cein : STD_LOGIC; 
  signal rx_output_ceinl_CEMUXNOT : STD_LOGIC; 
  signal rx_output_ceinl_GROM : STD_LOGIC; 
  signal rx_output_fifo_reset_FROM : STD_LOGIC; 
  signal rx_output_fifo_reset_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2441_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd6_In : STD_LOGIC; 
  signal tx_input_cs_FFd6_GROM : STD_LOGIC; 
  signal tx_input_n0023_GROM : STD_LOGIC; 
  signal mac_control_n0010_FROM : STD_LOGIC; 
  signal mac_control_n0010_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2746_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2746_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2739_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2739_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2762_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2762_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2731_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2731_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2971_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2770_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2770_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2777_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2777_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1609_GROM : STD_LOGIC; 
  signal mac_control_N73201_FROM : STD_LOGIC; 
  signal mac_control_N73201_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2421_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_0_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1586_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1616_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2755_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2755_GROM : STD_LOGIC; 
  signal mac_control_N73084_FROM : STD_LOGIC; 
  signal mac_control_N73084_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1593_GROM : STD_LOGIC; 
  signal slowclock_rxfl_LOGIC_ZERO : STD_LOGIC; 
  signal slowclock_rxfl_GROM : STD_LOGIC; 
  signal slowclock_txfl_LOGIC_ZERO : STD_LOGIC; 
  signal slowclock_txfl_GROM : STD_LOGIC; 
  signal tx_input_dh_3_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crccomb_n0118_1_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_n0118_1_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2472_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_crccomb_n0124_0_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_n0124_0_GROM : STD_LOGIC; 
  signal tx_input_dh_9_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_1_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_3_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_5_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2432_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_9_FFY_RST : STD_LOGIC; 
  signal txbp_9_FFX_RST : STD_LOGIC; 
  signal MDC_OBUF_FFY_RST : STD_LOGIC; 
  signal mac_control_CHOICE2448_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2448_GROM : STD_LOGIC; 
  signal mac_control_lmacaddr_1_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_1_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_3_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2441_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_5_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_5_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_7_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_7_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_9_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_9_FFY_RST : STD_LOGIC; 
  signal rxbp_1_FFX_RST : STD_LOGIC; 
  signal rxbp_1_FFY_RST : STD_LOGIC; 
  signal rxbp_1_CEMUXNOT : STD_LOGIC; 
  signal rxbp_3_FFY_RST : STD_LOGIC; 
  signal rxbp_3_CEMUXNOT : STD_LOGIC; 
  signal rxbp_5_FFY_RST : STD_LOGIC; 
  signal rxbp_5_CEMUXNOT : STD_LOGIC; 
  signal rxbp_7_FFY_RST : STD_LOGIC; 
  signal rxbp_7_CEMUXNOT : STD_LOGIC; 
  signal rxbp_9_FFY_RST : STD_LOGIC; 
  signal rxbp_9_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_1_FFY_RST : STD_LOGIC; 
  signal rxfbbp_1_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_3_FFY_RST : STD_LOGIC; 
  signal rxfbbp_3_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_5_FFY_RST : STD_LOGIC; 
  signal rxfbbp_5_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_7_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_9_FFY_RST : STD_LOGIC; 
  signal rxfbbp_9_CEMUXNOT : STD_LOGIC; 
  signal mac_control_CHOICE2486_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2486_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_3_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_5_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2472_FFX_SET : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_7_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2451_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_9_CEMUXNOT : STD_LOGIC; 
  signal mac_control_N82129_FROM : STD_LOGIC; 
  signal mac_control_N82129_GROM : STD_LOGIC; 
  signal rx_output_lenr_2_FROM : STD_LOGIC; 
  signal rx_output_lenr_2_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcl_25_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_9_Xo_0_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_9_Xo_0_GROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0118_1_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0118_1_GROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0124_0_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0124_0_GROM : STD_LOGIC; 
  signal rx_output_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd6_FROM : STD_LOGIC; 
  signal rx_output_cs_FFd6_In : STD_LOGIC; 
  signal rx_output_lenr_3_FROM : STD_LOGIC; 
  signal rx_output_lenr_3_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_4_FROM : STD_LOGIC; 
  signal rx_output_lenr_4_CEMUXNOT : STD_LOGIC; 
  signal rx_output_CHOICE1557_FROM : STD_LOGIC; 
  signal rx_output_CHOICE1557_GROM : STD_LOGIC; 
  signal rx_output_denl_FROM : STD_LOGIC; 
  signal rx_output_denl_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_CHOICE1529 : STD_LOGIC; 
  signal rx_output_lenr_5_FROM : STD_LOGIC; 
  signal rx_output_lenr_5_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_6_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_6_FROM : STD_LOGIC; 
  signal rx_output_lenr_6_CEMUXNOT : STD_LOGIC; 
  signal mac_control_dout_14_FROM : STD_LOGIC; 
  signal mac_control_N77791 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2503_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2503_GROM : STD_LOGIC; 
  signal tx_output_crcl_1_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2511_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2511_GROM : STD_LOGIC; 
  signal rx_output_lenr_7_FROM : STD_LOGIC; 
  signal rx_output_lenr_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2513_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2513_GROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_3_108_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_3_108_1_GROM : STD_LOGIC; 
  signal mac_control_dout_31_FROM : STD_LOGIC; 
  signal mac_control_N74276 : STD_LOGIC; 
  signal mac_control_dout_23_FROM : STD_LOGIC; 
  signal mac_control_N74572 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2451_FFX_SET : STD_LOGIC; 
  signal rx_output_lenr_8_FROM : STD_LOGIC; 
  signal rx_output_lenr_8_CEMUXNOT : STD_LOGIC; 
  signal tx_input_mrw_GROM : STD_LOGIC; 
  signal rx_output_lenr_9_FROM : STD_LOGIC; 
  signal rx_output_lenr_9_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1403_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1403_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_mcast_0_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_mcast_0_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2483_FFY_RST : STD_LOGIC; 
  signal tx_output_CHOICE1303_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1303_GROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_0_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_0_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_dout_15_FFY_RST : STD_LOGIC; 
  signal tx_output_CHOICE1336_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1336_GROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_1_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_N52163_FROM : STD_LOGIC; 
  signal mac_control_N52163_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1314_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1314_GROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_2_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_2_CEMUXNOT : STD_LOGIC; 
  signal tx_output_ncrcbytel_3_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_3_CEMUXNOT : STD_LOGIC; 
  signal tx_output_CHOICE1325_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1325_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_4_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_4_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_4_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2483_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_25_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2423_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_5_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_ncrcbytel_6_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_6_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_validbcast_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0051 : STD_LOGIC; 
  signal rx_input_memio_addrchk_validbcast_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N9_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_7_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_7_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_validucast_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0052 : STD_LOGIC; 
  signal rx_input_memio_addrchk_validucast_CEMUXNOT : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1774_GROM : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1781_GROM : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1796_GROM : STD_LOGIC; 
  signal LEDDPX_ENABLE : STD_LOGIC; 
  signal LEDDPX_TORGTS : STD_LOGIC; 
  signal LEDDPX_OUTMUX : STD_LOGIC; 
  signal mac_control_LEDDPX_OBUF : STD_LOGIC; 
  signal LEDDPX_OD : STD_LOGIC; 
  signal rx_input_GMII_RXD_0_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_1_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_2_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_3_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_4_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_5_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_6_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_7_IBUF : STD_LOGIC; 
  signal tx_input_DIN_10_IBUF : STD_LOGIC; 
  signal tx_input_DIN_11_IBUF : STD_LOGIC; 
  signal tx_input_DIN_12_IBUF : STD_LOGIC; 
  signal tx_input_DIN_13_IBUF : STD_LOGIC; 
  signal tx_input_DIN_14_IBUF : STD_LOGIC; 
  signal tx_input_DIN_15_IBUF : STD_LOGIC; 
  signal DOUT_0_ENABLE : STD_LOGIC; 
  signal DOUT_0_TORGTS : STD_LOGIC; 
  signal DOUT_0_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_0_OBUF : STD_LOGIC; 
  signal DOUT_0_OD : STD_LOGIC; 
  signal DOUT_1_ENABLE : STD_LOGIC; 
  signal DOUT_1_TORGTS : STD_LOGIC; 
  signal DOUT_1_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_1_OBUF : STD_LOGIC; 
  signal DOUT_1_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2397_FFX_SET : STD_LOGIC; 
  signal DOUT_2_ENABLE : STD_LOGIC; 
  signal DOUT_2_TORGTS : STD_LOGIC; 
  signal DOUT_2_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_2_OBUF : STD_LOGIC; 
  signal DOUT_2_OD : STD_LOGIC; 
  signal DOUT_3_ENABLE : STD_LOGIC; 
  signal DOUT_3_TORGTS : STD_LOGIC; 
  signal DOUT_3_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_3_OBUF : STD_LOGIC; 
  signal DOUT_3_OD : STD_LOGIC; 
  signal DOUT_4_ENABLE : STD_LOGIC; 
  signal DOUT_4_TORGTS : STD_LOGIC; 
  signal DOUT_4_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_4_OBUF : STD_LOGIC; 
  signal DOUT_4_OD : STD_LOGIC; 
  signal DOUT_5_ENABLE : STD_LOGIC; 
  signal DOUT_5_TORGTS : STD_LOGIC; 
  signal DOUT_5_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_5_OBUF : STD_LOGIC; 
  signal DOUT_5_OD : STD_LOGIC; 
  signal DOUT_6_ENABLE : STD_LOGIC; 
  signal DOUT_6_TORGTS : STD_LOGIC; 
  signal DOUT_6_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_6_OBUF : STD_LOGIC; 
  signal DOUT_6_OD : STD_LOGIC; 
  signal DOUT_7_ENABLE : STD_LOGIC; 
  signal DOUT_7_TORGTS : STD_LOGIC; 
  signal DOUT_7_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_7_OBUF : STD_LOGIC; 
  signal DOUT_7_OD : STD_LOGIC; 
  signal DOUT_8_ENABLE : STD_LOGIC; 
  signal DOUT_8_TORGTS : STD_LOGIC; 
  signal DOUT_8_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_8_OBUF : STD_LOGIC; 
  signal DOUT_8_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2499_FFY_RST : STD_LOGIC; 
  signal DOUT_9_ENABLE : STD_LOGIC; 
  signal DOUT_9_TORGTS : STD_LOGIC; 
  signal DOUT_9_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_9_OBUF : STD_LOGIC; 
  signal DOUT_9_OD : STD_LOGIC; 
  signal SOUT_ENABLE : STD_LOGIC; 
  signal SOUT_TORGTS : STD_LOGIC; 
  signal SOUT_OUTMUX : STD_LOGIC; 
  signal mac_control_SOUT_OBUF : STD_LOGIC; 
  signal SOUT_OD : STD_LOGIC; 
  signal mac_control_SCLK_IBUF : STD_LOGIC; 
  signal LEDRX_ENABLE : STD_LOGIC; 
  signal LEDRX_TORGTS : STD_LOGIC; 
  signal LEDRX_OUTMUX : STD_LOGIC; 
  signal mac_control_LEDRX_OBUF : STD_LOGIC; 
  signal LEDRX_OD : STD_LOGIC; 
  signal LEDTX_ENABLE : STD_LOGIC; 
  signal LEDTX_TORGTS : STD_LOGIC; 
  signal LEDTX_OUTMUX : STD_LOGIC; 
  signal mac_control_LEDTX_OBUF : STD_LOGIC; 
  signal LEDTX_OD : STD_LOGIC; 
  signal tx_input_DIN_0_IBUF : STD_LOGIC; 
  signal tx_input_DIN_1_IBUF : STD_LOGIC; 
  signal tx_input_DIN_2_IBUF : STD_LOGIC; 
  signal tx_input_DIN_3_IBUF : STD_LOGIC; 
  signal tx_input_DIN_4_IBUF : STD_LOGIC; 
  signal tx_input_DIN_5_IBUF : STD_LOGIC; 
  signal tx_input_DIN_6_IBUF : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2400_FFY_RST : STD_LOGIC; 
  signal tx_input_DIN_7_IBUF : STD_LOGIC; 
  signal tx_input_DIN_8_IBUF : STD_LOGIC; 
  signal tx_input_DIN_9_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RX_ER_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RX_DV_IBUF : STD_LOGIC; 
  signal MA_10_ENABLE : STD_LOGIC; 
  signal MA_10_TORGTS : STD_LOGIC; 
  signal MA_10_OUTMUX : STD_LOGIC; 
  signal MA_10_OCEMUXNOT : STD_LOGIC; 
  signal MA_10_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N13_FFX_RST : STD_LOGIC; 
  signal MA_11_ENABLE : STD_LOGIC; 
  signal MA_11_TORGTS : STD_LOGIC; 
  signal MA_11_OUTMUX : STD_LOGIC; 
  signal MA_11_OCEMUXNOT : STD_LOGIC; 
  signal MA_11_OD : STD_LOGIC; 
  signal MA_12_ENABLE : STD_LOGIC; 
  signal MA_12_TORGTS : STD_LOGIC; 
  signal MA_12_OUTMUX : STD_LOGIC; 
  signal MA_12_OCEMUXNOT : STD_LOGIC; 
  signal MA_12_OD : STD_LOGIC; 
  signal mac_control_n0037_FROM : STD_LOGIC; 
  signal mac_control_n0037_GROM : STD_LOGIC; 
  signal mac_control_n0044_GROM : STD_LOGIC; 
  signal mac_control_n0053_GROM : STD_LOGIC; 
  signal mac_control_n0045_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2473_FFY_SET : STD_LOGIC; 
  signal mac_control_n0054_GROM : STD_LOGIC; 
  signal mac_control_n0046_GROM : STD_LOGIC; 
  signal mac_control_n0055_GROM : STD_LOGIC; 
  signal mac_control_n0047_GROM : STD_LOGIC; 
  signal mac_control_n0048_GROM : STD_LOGIC; 
  signal mac_control_n0080_FROM : STD_LOGIC; 
  signal mac_control_n0080_GROM : STD_LOGIC; 
  signal mac_control_n0049_GROM : STD_LOGIC; 
  signal mac_control_N69420_FROM : STD_LOGIC; 
  signal mac_control_N69420_GROM : STD_LOGIC; 
  signal mac_control_n0081_FROM : STD_LOGIC; 
  signal mac_control_n0081_GROM : STD_LOGIC; 
  signal mac_control_n0085_FROM : STD_LOGIC; 
  signal mac_control_n0085_GROM : STD_LOGIC; 
  signal mac_control_txf_rst_FROM : STD_LOGIC; 
  signal mac_control_n0062 : STD_LOGIC; 
  signal mac_control_n0082_FROM : STD_LOGIC; 
  signal mac_control_n0082_GROM : STD_LOGIC; 
  signal mac_control_n0083_FROM : STD_LOGIC; 
  signal mac_control_n0083_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2453_FFY_SET : STD_LOGIC; 
  signal mac_control_n0076_FROM : STD_LOGIC; 
  signal mac_control_n0076_GROM : STD_LOGIC; 
  signal mac_control_n0084_FROM : STD_LOGIC; 
  signal mac_control_n0084_GROM : STD_LOGIC; 
  signal mac_control_n0077_FROM : STD_LOGIC; 
  signal mac_control_n0077_GROM : STD_LOGIC; 
  signal mac_control_n0087_FROM : STD_LOGIC; 
  signal mac_control_n0087_GROM : STD_LOGIC; 
  signal mac_control_n0079_FROM : STD_LOGIC; 
  signal mac_control_n0079_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2600_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2600_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2443_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_27_FROM : STD_LOGIC; 
  signal mac_control_N74720 : STD_LOGIC; 
  signal mac_control_dout_19_FROM : STD_LOGIC; 
  signal mac_control_N74424 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE1201_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE1201_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE1541_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE1541_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_30_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0030_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0031_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd7_In : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd7_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1424_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd5_In : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd5_GROM : STD_LOGIC; 
  signal tx_output_addrl_11_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0028_GROM : STD_LOGIC; 
  signal tx_output_addrl_13_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1431_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0029_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2473_FFX_SET : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_3_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_3_CEMUXNOT : STD_LOGIC; 
  signal tx_output_addrl_15_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1417_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_0_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_0_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_5_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_5_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1438_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_2_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_2_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1410_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_4_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_4_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_0_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_1_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_cs_FFd15_FROM : STD_LOGIC; 
  signal tx_output_cs_FFd16_In : STD_LOGIC; 
  signal rx_input_memio_crcl_1_FROM : STD_LOGIC; 
  signal tx_output_N81617_FROM : STD_LOGIC; 
  signal tx_output_N81617_GROM : STD_LOGIC; 
  signal tx_output_crcl_30_FROM : STD_LOGIC; 
  signal mac_control_N81817_FROM : STD_LOGIC; 
  signal mac_control_N81817_GROM : STD_LOGIC; 
  signal rx_input_memio_n0049 : STD_LOGIC; 
  signal rx_input_memio_crcen_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcen_GROM : STD_LOGIC; 
  signal rx_input_memio_cs_Out916_2_FROM : STD_LOGIC; 
  signal rx_input_memio_cs_Out916_2_GROM : STD_LOGIC; 
  signal rx_input_memio_n0031_GROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd8_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd8_GROM : STD_LOGIC; 
  signal rx_input_memio_n0033_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_5_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2453_FFX_SET : STD_LOGIC; 
  signal rx_input_memio_n0044_GROM : STD_LOGIC; 
  signal rx_input_memio_n0046_GROM : STD_LOGIC; 
  signal rx_input_memio_n0047_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE2913_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1821_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1821_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2486_FFY_RST : STD_LOGIC; 
  signal mac_control_CHOICE2662_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2662_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_n0011_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_n0011_GROM : STD_LOGIC; 
  signal tx_output_N81605_FROM : STD_LOGIC; 
  signal tx_output_N81605_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11_FFY_RST : STD_LOGIC; 
  signal mac_control_N81753_FROM : STD_LOGIC; 
  signal mac_control_N81753_GROM : STD_LOGIC; 
  signal tx_output_bcntl_12_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_14_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_14_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_15_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_15_CEMUXNOT : STD_LOGIC; 
  signal rx_output_bpl_11_CEMUXNOT : STD_LOGIC; 
  signal rx_output_bpl_13_FFY_RST : STD_LOGIC; 
  signal rx_output_bpl_13_CEMUXNOT : STD_LOGIC; 
  signal rx_output_bpl_15_FFY_RST : STD_LOGIC; 
  signal rx_output_bpl_15_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifo_N1546_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N2499 : STD_LOGIC; 
  signal rx_output_fifo_N1610_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N3427 : STD_LOGIC; 
  signal rx_output_fifo_N1563_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2486_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1567_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1627_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N19_FROM : STD_LOGIC; 
  signal rx_output_fifo_N19_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1565_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1629_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1633_FFY_RST : STD_LOGIC; 
  signal q2_21_FFY_RST : STD_LOGIC; 
  signal q2_13_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1631_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1573_FFY_RST : STD_LOGIC; 
  signal q2_31_FFY_RST : STD_LOGIC; 
  signal q2_15_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1577_FFY_SET : STD_LOGIC; 
  signal mac_control_phystat_11_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1575_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1517_GROM : STD_LOGIC; 
  signal q2_17_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd18_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd18_FROM : STD_LOGIC; 
  signal rx_output_cs_FFd18_In : STD_LOGIC; 
  signal rx_output_fifo_N1609_FFY_SET : STD_LOGIC; 
  signal mac_control_phystat_21_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_13_FFY_RST : STD_LOGIC; 
  signal q2_27_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2436_FFY_SET : STD_LOGIC; 
  signal q2_19_FFY_RST : STD_LOGIC; 
  signal q3_11_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1585_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_23_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_31_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1571_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2425_FFY_SET : STD_LOGIC; 
  signal q2_29_FFY_RST : STD_LOGIC; 
  signal q3_21_FFY_RST : STD_LOGIC; 
  signal q3_13_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1586_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N3974 : STD_LOGIC; 
  signal rx_output_fifo_N1591_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N3970 : STD_LOGIC; 
  signal rx_output_fifo_N1591_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1603_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1607_FFY_SET : STD_LOGIC; 
  signal mac_control_phystat_25_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_17_FFY_RST : STD_LOGIC; 
  signal q3_31_FFY_RST : STD_LOGIC; 
  signal q3_23_FFY_RST : STD_LOGIC; 
  signal q3_15_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1579_FFY_SET : STD_LOGIC; 
  signal mac_control_phystat_19_FFY_RST : STD_LOGIC; 
  signal q3_25_FFY_RST : STD_LOGIC; 
  signal q3_17_FFY_RST : STD_LOGIC; 
  signal memcontroller_wen : STD_LOGIC; 
  signal memcontroller_oe_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2425_FFX_RST : STD_LOGIC; 
  signal q3_27_FFY_RST : STD_LOGIC; 
  signal q3_19_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1581_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2445_FFY_RST : STD_LOGIC; 
  signal q3_29_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd17_FFY_SET : STD_LOGIC; 
  signal tx_output_cs_FFd17_FROM : STD_LOGIC; 
  signal tx_output_cs_FFd17_In : STD_LOGIC; 
  signal rx_output_ceinll_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0013_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0013_GROM : STD_LOGIC; 
  signal tx_output_crcl_10_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0016_GROM : STD_LOGIC; 
  signal tx_output_addrl_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_addrl_3_FFY_RST : STD_LOGIC; 
  signal tx_output_addrl_3_CEMUXNOT : STD_LOGIC; 
  signal tx_output_addrl_5_FFY_RST : STD_LOGIC; 
  signal tx_output_addrl_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_addrl_7_FFY_RST : STD_LOGIC; 
  signal tx_output_addrl_7_CEMUXNOT : STD_LOGIC; 
  signal rx_output_len_11_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2436_FFX_SET : STD_LOGIC; 
  signal rx_output_mdl_11_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_11_CEMUXNOT : STD_LOGIC; 
  signal tx_output_addrl_9_CEMUXNOT : STD_LOGIC; 
  signal rx_output_len_13_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_21_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_21_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_13_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_13_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_31_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_31_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_23_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_23_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_15_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_15_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2445_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_25_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_17_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_17_CEMUXNOT : STD_LOGIC; 
  signal mac_control_CHOICE2693_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2693_GROM : STD_LOGIC; 
  signal rx_output_mdl_27_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_19_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_19_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_29_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_29_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lmasell_FFY_RST : STD_LOGIC; 
  signal rx_output_lmasell_CEMUXNOT : STD_LOGIC; 
  signal tx_output_cs_FFd3_FROM : STD_LOGIC; 
  signal tx_output_cs_FFd4_In : STD_LOGIC; 
  signal tx_input_enable_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_crcl_3_FROM : STD_LOGIC; 
  signal mac_control_N82125_FROM : STD_LOGIC; 
  signal mac_control_N82125_GROM : STD_LOGIC; 
  signal txfifofull_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2475_FFX_SET : STD_LOGIC; 
  signal mac_control_CHOICE2631_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2631_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2455_FFY_SET : STD_LOGIC; 
  signal tx_output_bcntl_2_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_4_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_4_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_6_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_6_CEMUXNOT : STD_LOGIC; 
  signal rx_output_bpl_1_FFY_RST : STD_LOGIC; 
  signal rx_output_bpl_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_8_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_8_CEMUXNOT : STD_LOGIC; 
  signal rx_output_bpl_3_FFY_RST : STD_LOGIC; 
  signal rx_output_bpl_3_CEMUXNOT : STD_LOGIC; 
  signal tx_output_datal_1_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_10_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_10_CEMUXNOT : STD_LOGIC; 
  signal rx_output_bpl_5_FFY_RST : STD_LOGIC; 
  signal rx_output_bpl_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_datal_3_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_3_CEMUXNOT : STD_LOGIC; 
  signal rx_output_bpl_7_FFY_RST : STD_LOGIC; 
  signal rx_output_bpl_7_CEMUXNOT : STD_LOGIC; 
  signal tx_output_datal_5_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_11_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_11_FROM : STD_LOGIC; 
  signal rx_output_bpl_9_CEMUXNOT : STD_LOGIC; 
  signal tx_output_datal_7_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_dout_1_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_1_FROM : STD_LOGIC; 
  signal mac_control_N76543 : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_2_GROM : STD_LOGIC; 
  signal rx_output_mdl_1_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_1_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_3_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_3_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_5_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_5_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_7_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_7_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2455_FFX_SET : STD_LOGIC; 
  signal rx_output_mdl_9_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_9_CEMUXNOT : STD_LOGIC; 
  signal tx_output_N70584_FROM : STD_LOGIC; 
  signal tx_output_N70584_GROM : STD_LOGIC; 
  signal rx_input_GMII_ro_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_n00561_2_FROM : STD_LOGIC; 
  signal mac_control_n00561_2_GROM : STD_LOGIC; 
  signal tx_output_outselll_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_outselll_3_CEMUXNOT : STD_LOGIC; 
  signal tx_output_N70557_FROM : STD_LOGIC; 
  signal tx_output_N70557_GROM : STD_LOGIC; 
  signal tx_output_N70530_FROM : STD_LOGIC; 
  signal tx_output_N70530_GROM : STD_LOGIC; 
  signal rx_input_fifo_dout_9_FFY_RST : STD_LOGIC; 
  signal tx_output_data_0_FROM : STD_LOGIC; 
  signal tx_output_data_0_CEMUXNOT : STD_LOGIC; 
  signal tx_output_data_1_FROM : STD_LOGIC; 
  signal tx_output_data_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_12_FROM : STD_LOGIC; 
  signal tx_output_data_2_FROM : STD_LOGIC; 
  signal tx_output_data_2_CEMUXNOT : STD_LOGIC; 
  signal tx_output_data_3_FROM : STD_LOGIC; 
  signal tx_output_data_3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_dout_2_FROM : STD_LOGIC; 
  signal mac_control_N76751 : STD_LOGIC; 
  signal tx_output_data_4_FROM : STD_LOGIC; 
  signal tx_output_data_4_CEMUXNOT : STD_LOGIC; 
  signal tx_output_N70503_FROM : STD_LOGIC; 
  signal tx_output_N70503_GROM : STD_LOGIC; 
  signal tx_output_data_5_FROM : STD_LOGIC; 
  signal tx_output_data_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_data_6_FROM : STD_LOGIC; 
  signal tx_output_data_6_CEMUXNOT : STD_LOGIC; 
  signal tx_output_data_7_FROM : STD_LOGIC; 
  signal tx_output_data_7_CEMUXNOT : STD_LOGIC; 
  signal tx_output_cs_Out1160_2_FROM : STD_LOGIC; 
  signal tx_output_cs_Out1160_2_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1229_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1229_GROM : STD_LOGIC; 
  signal tx_output_N69304_FROM : STD_LOGIC; 
  signal tx_output_N69304_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1265_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1265_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1205_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1205_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1217_GROM : STD_LOGIC; 
  signal RESET_IBUF_1_FROM : STD_LOGIC; 
  signal RESET_IBUF_1_GROM : STD_LOGIC; 
  signal RESET_IBUF_2_FROM : STD_LOGIC; 
  signal RESET_IBUF_2_GROM : STD_LOGIC; 
  signal MDIO_ENABLE : STD_LOGIC; 
  signal MDIO_TORGTS : STD_LOGIC; 
  signal MDIO_OUTMUX : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_sin : STD_LOGIC; 
  signal rx_input_fifo_fifo_empty_FFX_SET : STD_LOGIC; 
  signal DOUT_10_ENABLE : STD_LOGIC; 
  signal DOUT_10_TORGTS : STD_LOGIC; 
  signal DOUT_10_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_10_OBUF : STD_LOGIC; 
  signal DOUT_10_OD : STD_LOGIC; 
  signal DOUT_11_ENABLE : STD_LOGIC; 
  signal DOUT_11_TORGTS : STD_LOGIC; 
  signal DOUT_11_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_11_OBUF : STD_LOGIC; 
  signal DOUT_11_OD : STD_LOGIC; 
  signal DOUT_12_ENABLE : STD_LOGIC; 
  signal DOUT_12_TORGTS : STD_LOGIC; 
  signal DOUT_12_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_12_OBUF : STD_LOGIC; 
  signal DOUT_12_OD : STD_LOGIC; 
  signal DOUT_13_ENABLE : STD_LOGIC; 
  signal DOUT_13_TORGTS : STD_LOGIC; 
  signal DOUT_13_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_13_OBUF : STD_LOGIC; 
  signal DOUT_13_OD : STD_LOGIC; 
  signal DOUT_14_ENABLE : STD_LOGIC; 
  signal DOUT_14_TORGTS : STD_LOGIC; 
  signal DOUT_14_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_14_OBUF : STD_LOGIC; 
  signal DOUT_14_OD : STD_LOGIC; 
  signal DOUT_15_ENABLE : STD_LOGIC; 
  signal DOUT_15_TORGTS : STD_LOGIC; 
  signal DOUT_15_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_15_OBUF : STD_LOGIC; 
  signal DOUT_15_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2497_FFY_SET : STD_LOGIC; 
  signal MDC_ENABLE : STD_LOGIC; 
  signal MDC_TORGTS : STD_LOGIC; 
  signal MDC_OUTMUX : STD_LOGIC; 
  signal SCS_IBUF_1 : STD_LOGIC; 
  signal SIN_IBUF_2 : STD_LOGIC; 
  signal LED100_ENABLE : STD_LOGIC; 
  signal LED100_TORGTS : STD_LOGIC; 
  signal LED100_OUTMUX : STD_LOGIC; 
  signal mac_control_LED100_OBUF : STD_LOGIC; 
  signal LED100_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2397_FFY_RST : STD_LOGIC; 
  signal MCLK_ENABLE : STD_LOGIC; 
  signal MCLK_TORGTS : STD_LOGIC; 
  signal MCLK_OUTMUX : STD_LOGIC; 
  signal tx_input_NEWFRAME_IBUF : STD_LOGIC; 
  signal LED1000_ENABLE : STD_LOGIC; 
  signal LED1000_TORGTS : STD_LOGIC; 
  signal LED1000_OUTMUX : STD_LOGIC; 
  signal mac_control_LED1000_OBUF : STD_LOGIC; 
  signal LED1000_OD : STD_LOGIC; 
  signal TX_EN_ENABLE : STD_LOGIC; 
  signal TX_EN_TORGTS : STD_LOGIC; 
  signal TX_EN_OUTMUX : STD_LOGIC; 
  signal tx_output_TXEN : STD_LOGIC; 
  signal TX_EN_OCEMUXNOT : STD_LOGIC; 
  signal TX_EN_OD : STD_LOGIC; 
  signal DOUTEN_ENABLE : STD_LOGIC; 
  signal DOUTEN_TORGTS : STD_LOGIC; 
  signal DOUTEN_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUTEN_OBUF : STD_LOGIC; 
  signal DOUTEN_OD : STD_LOGIC; 
  signal MWE_ENABLE : STD_LOGIC; 
  signal MWE_TORGTS : STD_LOGIC; 
  signal MWE_OUTMUX : STD_LOGIC; 
  signal memcontroller_WEEXT : STD_LOGIC; 
  signal MWE_OCEMUXNOT : STD_LOGIC; 
  signal MWE_OD : STD_LOGIC; 
  signal RESET_IBUF_3 : STD_LOGIC; 
  signal rx_output_NEXTFRAME_IBUF : STD_LOGIC; 
  signal LEDACT_ENABLE : STD_LOGIC; 
  signal LEDACT_TORGTS : STD_LOGIC; 
  signal LEDACT_OUTMUX : STD_LOGIC; 
  signal mac_control_LEDACT_OBUF : STD_LOGIC; 
  signal LEDACT_OD : STD_LOGIC; 
  signal TXD_0_ENABLE : STD_LOGIC; 
  signal TXD_0_TORGTS : STD_LOGIC; 
  signal TXD_0_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_0_OBUF : STD_LOGIC; 
  signal TXD_0_OCEMUXNOT : STD_LOGIC; 
  signal TXD_0_OD : STD_LOGIC; 
  signal TXD_1_ENABLE : STD_LOGIC; 
  signal TXD_1_TORGTS : STD_LOGIC; 
  signal TXD_1_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_1_OBUF : STD_LOGIC; 
  signal TXD_1_OCEMUXNOT : STD_LOGIC; 
  signal TXD_1_OD : STD_LOGIC; 
  signal TXD_2_ENABLE : STD_LOGIC; 
  signal TXD_2_TORGTS : STD_LOGIC; 
  signal TXD_2_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_2_OBUF : STD_LOGIC; 
  signal TXD_2_OCEMUXNOT : STD_LOGIC; 
  signal TXD_2_OD : STD_LOGIC; 
  signal TXD_3_ENABLE : STD_LOGIC; 
  signal TXD_3_TORGTS : STD_LOGIC; 
  signal TXD_3_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_3_OBUF : STD_LOGIC; 
  signal TXD_3_OCEMUXNOT : STD_LOGIC; 
  signal TXD_3_OD : STD_LOGIC; 
  signal TXD_4_ENABLE : STD_LOGIC; 
  signal TXD_4_TORGTS : STD_LOGIC; 
  signal TXD_4_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_4_OBUF : STD_LOGIC; 
  signal TXD_4_OCEMUXNOT : STD_LOGIC; 
  signal TXD_4_OD : STD_LOGIC; 
  signal TXD_5_ENABLE : STD_LOGIC; 
  signal TXD_5_TORGTS : STD_LOGIC; 
  signal TXD_5_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_5_OBUF : STD_LOGIC; 
  signal TXD_5_OCEMUXNOT : STD_LOGIC; 
  signal TXD_5_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N13_FFY_RST : STD_LOGIC; 
  signal TXD_6_ENABLE : STD_LOGIC; 
  signal TXD_6_TORGTS : STD_LOGIC; 
  signal TXD_6_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_6_OBUF : STD_LOGIC; 
  signal TXD_6_OCEMUXNOT : STD_LOGIC; 
  signal TXD_6_OD : STD_LOGIC; 
  signal TXD_7_ENABLE : STD_LOGIC; 
  signal TXD_7_TORGTS : STD_LOGIC; 
  signal TXD_7_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_7_OBUF : STD_LOGIC; 
  signal TXD_7_OCEMUXNOT : STD_LOGIC; 
  signal TXD_7_OD : STD_LOGIC; 
  signal tx_output_crcl_23_FROM : STD_LOGIC; 
  signal tx_output_crcl_15_FROM : STD_LOGIC; 
  signal mac_control_dout_5_FROM : STD_LOGIC; 
  signal mac_control_N77167 : STD_LOGIC; 
  signal rx_input_memio_crcl_10_FROM : STD_LOGIC; 
  signal mac_control_lmacaddr_47_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_8_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2382_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2382_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2458_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2458_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2306_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2306_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2420_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2420_GROM : STD_LOGIC; 
  signal memcontroller_dnl2_11_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_21_CEMUXNOT : STD_LOGIC; 
  signal rxbp_11_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_13_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_31_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_23_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_15_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_25_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_17_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_27_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_19_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_29_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_datal_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_datal_3_CEMUXNOT : STD_LOGIC; 
  signal rxbp_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_datal_5_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_datal_7_CEMUXNOT : STD_LOGIC; 
  signal rxbp_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_0_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_0_rt : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_0_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_0_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_2_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_2_rt : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_2_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_2_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_4_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_4_rt : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_4_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_4_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_24_FROM : STD_LOGIC; 
  signal tx_output_crcl_16_FROM : STD_LOGIC; 
  signal mac_control_dout_6_FROM : STD_LOGIC; 
  signal mac_control_N76959 : STD_LOGIC; 
  signal rx_input_memio_crcl_11_FROM : STD_LOGIC; 
  signal mac_control_n0238_FROM : STD_LOGIC; 
  signal mac_control_n0238_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_9_FROM : STD_LOGIC; 
  signal MA_13_ENABLE : STD_LOGIC; 
  signal MA_13_TORGTS : STD_LOGIC; 
  signal MA_13_OUTMUX : STD_LOGIC; 
  signal MA_13_OCEMUXNOT : STD_LOGIC; 
  signal MA_13_OD : STD_LOGIC; 
  signal MA_14_ENABLE : STD_LOGIC; 
  signal MA_14_TORGTS : STD_LOGIC; 
  signal MA_14_OUTMUX : STD_LOGIC; 
  signal MA_14_OCEMUXNOT : STD_LOGIC; 
  signal MA_14_OD : STD_LOGIC; 
  signal MA_15_ENABLE : STD_LOGIC; 
  signal MA_15_TORGTS : STD_LOGIC; 
  signal MA_15_OUTMUX : STD_LOGIC; 
  signal MA_15_OCEMUXNOT : STD_LOGIC; 
  signal MA_15_OD : STD_LOGIC; 
  signal MA_16_ENABLE : STD_LOGIC; 
  signal MA_16_TORGTS : STD_LOGIC; 
  signal MA_16_OUTMUX : STD_LOGIC; 
  signal MA_16_OCEMUXNOT : STD_LOGIC; 
  signal MA_16_OD : STD_LOGIC; 
  signal MD_10_ENABLE : STD_LOGIC; 
  signal MD_10_TORGTS : STD_LOGIC; 
  signal MD_10_OUTMUX : STD_LOGIC; 
  signal MD_10_OD : STD_LOGIC; 
  signal MD_11_ENABLE : STD_LOGIC; 
  signal MD_11_TORGTS : STD_LOGIC; 
  signal MD_11_OUTMUX : STD_LOGIC; 
  signal MD_11_OD : STD_LOGIC; 
  signal MD_20_ENABLE : STD_LOGIC; 
  signal MD_20_TORGTS : STD_LOGIC; 
  signal MD_20_OUTMUX : STD_LOGIC; 
  signal MD_20_OD : STD_LOGIC; 
  signal MD_12_ENABLE : STD_LOGIC; 
  signal MD_12_TORGTS : STD_LOGIC; 
  signal MD_12_OUTMUX : STD_LOGIC; 
  signal MD_12_OD : STD_LOGIC; 
  signal MD_21_ENABLE : STD_LOGIC; 
  signal MD_21_TORGTS : STD_LOGIC; 
  signal MD_21_OUTMUX : STD_LOGIC; 
  signal MD_21_OD : STD_LOGIC; 
  signal MD_13_ENABLE : STD_LOGIC; 
  signal MD_13_TORGTS : STD_LOGIC; 
  signal MD_13_OUTMUX : STD_LOGIC; 
  signal MD_13_OD : STD_LOGIC; 
  signal MD_22_ENABLE : STD_LOGIC; 
  signal MD_22_TORGTS : STD_LOGIC; 
  signal MD_22_OUTMUX : STD_LOGIC; 
  signal MD_22_OD : STD_LOGIC; 
  signal MD_14_ENABLE : STD_LOGIC; 
  signal MD_14_TORGTS : STD_LOGIC; 
  signal MD_14_OUTMUX : STD_LOGIC; 
  signal MD_14_OD : STD_LOGIC; 
  signal MD_30_ENABLE : STD_LOGIC; 
  signal MD_30_TORGTS : STD_LOGIC; 
  signal MD_30_OUTMUX : STD_LOGIC; 
  signal MD_30_OD : STD_LOGIC; 
  signal MD_23_ENABLE : STD_LOGIC; 
  signal MD_23_TORGTS : STD_LOGIC; 
  signal MD_23_OUTMUX : STD_LOGIC; 
  signal MD_23_OD : STD_LOGIC; 
  signal MD_15_ENABLE : STD_LOGIC; 
  signal MD_15_TORGTS : STD_LOGIC; 
  signal MD_15_OUTMUX : STD_LOGIC; 
  signal MD_15_OD : STD_LOGIC; 
  signal MD_31_TFF_RST : STD_LOGIC; 
  signal MD_31_OFF_RST : STD_LOGIC; 
  signal MD_31_ENABLE : STD_LOGIC; 
  signal MD_31_TORGTS : STD_LOGIC; 
  signal MD_31_OUTMUX : STD_LOGIC; 
  signal MD_31_OD : STD_LOGIC; 
  signal MD_24_TFF_RST : STD_LOGIC; 
  signal MD_24_OFF_RST : STD_LOGIC; 
  signal MD_24_IFF_RST : STD_LOGIC; 
  signal MD_24_ENABLE : STD_LOGIC; 
  signal MD_24_TORGTS : STD_LOGIC; 
  signal MD_24_OUTMUX : STD_LOGIC; 
  signal MD_24_OD : STD_LOGIC; 
  signal MD_16_TFF_RST : STD_LOGIC; 
  signal MD_16_OFF_RST : STD_LOGIC; 
  signal MD_16_IFF_RST : STD_LOGIC; 
  signal MD_16_ENABLE : STD_LOGIC; 
  signal MD_16_TORGTS : STD_LOGIC; 
  signal MD_16_OUTMUX : STD_LOGIC; 
  signal MD_16_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2400_FFX_RST : STD_LOGIC; 
  signal MD_17_TFF_RST : STD_LOGIC; 
  signal MD_17_OFF_RST : STD_LOGIC; 
  signal MD_17_IFF_RST : STD_LOGIC; 
  signal MD_17_ENABLE : STD_LOGIC; 
  signal MD_17_TORGTS : STD_LOGIC; 
  signal MD_17_OUTMUX : STD_LOGIC; 
  signal MD_17_OD : STD_LOGIC; 
  signal MD_25_TFF_RST : STD_LOGIC; 
  signal MD_25_OFF_RST : STD_LOGIC; 
  signal MD_25_IFF_RST : STD_LOGIC; 
  signal MD_25_ENABLE : STD_LOGIC; 
  signal MD_25_TORGTS : STD_LOGIC; 
  signal MD_25_OUTMUX : STD_LOGIC; 
  signal MD_25_OD : STD_LOGIC; 
  signal MD_18_TFF_RST : STD_LOGIC; 
  signal MD_18_OFF_RST : STD_LOGIC; 
  signal MD_18_IFF_RST : STD_LOGIC; 
  signal MD_18_ENABLE : STD_LOGIC; 
  signal MD_18_TORGTS : STD_LOGIC; 
  signal MD_18_OUTMUX : STD_LOGIC; 
  signal MD_18_OD : STD_LOGIC; 
  signal MD_26_IFF_RST : STD_LOGIC; 
  signal MD_26_ENABLE : STD_LOGIC; 
  signal MD_26_TORGTS : STD_LOGIC; 
  signal MD_26_OUTMUX : STD_LOGIC; 
  signal MD_26_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2500_FFY_RST : STD_LOGIC; 
  signal MD_19_ENABLE : STD_LOGIC; 
  signal MD_19_TORGTS : STD_LOGIC; 
  signal MD_19_OUTMUX : STD_LOGIC; 
  signal MD_19_OD : STD_LOGIC; 
  signal MD_27_ENABLE : STD_LOGIC; 
  signal MD_27_TORGTS : STD_LOGIC; 
  signal MD_27_OUTMUX : STD_LOGIC; 
  signal MD_27_OD : STD_LOGIC; 
  signal MD_28_ENABLE : STD_LOGIC; 
  signal MD_28_TORGTS : STD_LOGIC; 
  signal MD_28_OUTMUX : STD_LOGIC; 
  signal MD_28_OD : STD_LOGIC; 
  signal MD_29_ENABLE : STD_LOGIC; 
  signal MD_29_TORGTS : STD_LOGIC; 
  signal MD_29_OUTMUX : STD_LOGIC; 
  signal MD_29_OD : STD_LOGIC; 
  signal LEDPOWER_ENABLE : STD_LOGIC; 
  signal LEDPOWER_TORGTS : STD_LOGIC; 
  signal LEDPOWER_OUTMUX : STD_LOGIC; 
  signal LEDPOWER_LOGIC_ONE : STD_LOGIC; 
  signal MA_0_ENABLE : STD_LOGIC; 
  signal MA_0_TORGTS : STD_LOGIC; 
  signal MA_0_OUTMUX : STD_LOGIC; 
  signal MA_0_OCEMUXNOT : STD_LOGIC; 
  signal MA_0_OD : STD_LOGIC; 
  signal MA_1_ENABLE : STD_LOGIC; 
  signal MA_1_TORGTS : STD_LOGIC; 
  signal MA_1_OUTMUX : STD_LOGIC; 
  signal MA_1_OCEMUXNOT : STD_LOGIC; 
  signal MA_1_OD : STD_LOGIC; 
  signal MA_2_ENABLE : STD_LOGIC; 
  signal MA_2_TORGTS : STD_LOGIC; 
  signal MA_2_OUTMUX : STD_LOGIC; 
  signal MA_2_OCEMUXNOT : STD_LOGIC; 
  signal MA_2_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2499_FFX_RST : STD_LOGIC; 
  signal MA_3_ENABLE : STD_LOGIC; 
  signal MA_3_TORGTS : STD_LOGIC; 
  signal MA_3_OUTMUX : STD_LOGIC; 
  signal MA_3_OCEMUXNOT : STD_LOGIC; 
  signal MA_3_OD : STD_LOGIC; 
  signal MA_4_ENABLE : STD_LOGIC; 
  signal MA_4_TORGTS : STD_LOGIC; 
  signal MA_4_OUTMUX : STD_LOGIC; 
  signal MA_4_OCEMUXNOT : STD_LOGIC; 
  signal MA_4_OD : STD_LOGIC; 
  signal MA_5_ENABLE : STD_LOGIC; 
  signal MA_5_TORGTS : STD_LOGIC; 
  signal MA_5_OUTMUX : STD_LOGIC; 
  signal MA_5_OCEMUXNOT : STD_LOGIC; 
  signal MA_5_OD : STD_LOGIC; 
  signal MA_6_ENABLE : STD_LOGIC; 
  signal MA_6_TORGTS : STD_LOGIC; 
  signal MA_6_OUTMUX : STD_LOGIC; 
  signal MA_6_OCEMUXNOT : STD_LOGIC; 
  signal MA_6_OD : STD_LOGIC; 
  signal MA_7_ENABLE : STD_LOGIC; 
  signal MA_7_TORGTS : STD_LOGIC; 
  signal MA_7_OUTMUX : STD_LOGIC; 
  signal MA_7_OCEMUXNOT : STD_LOGIC; 
  signal MA_7_OD : STD_LOGIC; 
  signal MA_8_ENABLE : STD_LOGIC; 
  signal MA_8_TORGTS : STD_LOGIC; 
  signal MA_8_OUTMUX : STD_LOGIC; 
  signal MA_8_OCEMUXNOT : STD_LOGIC; 
  signal MA_8_OD : STD_LOGIC; 
  signal MA_9_ENABLE : STD_LOGIC; 
  signal MA_9_TORGTS : STD_LOGIC; 
  signal MA_9_OUTMUX : STD_LOGIC; 
  signal MA_9_OCEMUXNOT : STD_LOGIC; 
  signal MA_9_OD : STD_LOGIC; 
  signal PHYRESET_ENABLE : STD_LOGIC; 
  signal PHYRESET_TORGTS : STD_LOGIC; 
  signal PHYRESET_OUTMUX : STD_LOGIC; 
  signal mac_control_PHYRESET_OBUF : STD_LOGIC; 
  signal PHYRESET_OD : STD_LOGIC; 
  signal MD_0_ENABLE : STD_LOGIC; 
  signal MD_0_TORGTS : STD_LOGIC; 
  signal MD_0_OUTMUX : STD_LOGIC; 
  signal MD_0_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15_FFY_RST : STD_LOGIC; 
  signal MD_1_ENABLE : STD_LOGIC; 
  signal MD_1_TORGTS : STD_LOGIC; 
  signal MD_1_OUTMUX : STD_LOGIC; 
  signal MD_1_OD : STD_LOGIC; 
  signal MD_2_ENABLE : STD_LOGIC; 
  signal MD_2_TORGTS : STD_LOGIC; 
  signal MD_2_OUTMUX : STD_LOGIC; 
  signal MD_2_OD : STD_LOGIC; 
  signal MD_3_ENABLE : STD_LOGIC; 
  signal MD_3_TORGTS : STD_LOGIC; 
  signal MD_3_OUTMUX : STD_LOGIC; 
  signal MD_3_OD : STD_LOGIC; 
  signal MD_4_ENABLE : STD_LOGIC; 
  signal MD_4_TORGTS : STD_LOGIC; 
  signal MD_4_OUTMUX : STD_LOGIC; 
  signal MD_4_OD : STD_LOGIC; 
  signal MD_5_ENABLE : STD_LOGIC; 
  signal MD_5_TORGTS : STD_LOGIC; 
  signal MD_5_OUTMUX : STD_LOGIC; 
  signal MD_5_OD : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd2_In : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd1_In : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4_In : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd3_In : STD_LOGIC; 
  signal rx_output_cs_FFd2_In : STD_LOGIC; 
  signal rx_output_cs_FFd1_In : STD_LOGIC; 
  signal mac_control_lmacaddr_23_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd4_In : STD_LOGIC; 
  signal rx_output_cs_FFd3_In : STD_LOGIC; 
  signal rx_output_cs_FFd8_In : STD_LOGIC; 
  signal rx_output_cs_FFd7_In : STD_LOGIC; 
  signal tx_input_cs_FFd2_In : STD_LOGIC; 
  signal tx_input_cs_FFd3_In : STD_LOGIC; 
  signal tx_input_cs_FFd8_In : STD_LOGIC; 
  signal tx_input_cs_FFd7_In : STD_LOGIC; 
  signal tx_input_cs_FFd9_In : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_10_59_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_10_net14 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_10_59_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_11_58_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_11_net12 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_11_58_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_12_57_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_12_net10 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_12_57_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_13_56_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_13_net8 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_13_56_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_14_55_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_14_net6 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_14_55_CEMUXNOT : STD_LOGIC; 
  signal mac_control_lmacaddr_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_15_54_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_15_net4 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_15_54_CEMUXNOT : STD_LOGIC; 
  signal mac_control_Mshreg_sinlll_net185 : STD_LOGIC; 
  signal mac_control_phyaddr_31_FROM : STD_LOGIC; 
  signal mac_control_phyaddr_31_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1551_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N2339 : STD_LOGIC; 
  signal rx_output_fifo_N2379 : STD_LOGIC; 
  signal rx_output_fifo_N2419 : STD_LOGIC; 
  signal rx_output_fifo_N2459 : STD_LOGIC; 
  signal rx_output_fifo_N3267 : STD_LOGIC; 
  signal rx_output_fifo_N3307 : STD_LOGIC; 
  signal rx_output_fifo_N3187 : STD_LOGIC; 
  signal rx_output_fifo_N3227 : STD_LOGIC; 
  signal rx_output_fifo_N3347 : STD_LOGIC; 
  signal rx_output_fifo_N3387 : STD_LOGIC; 
  signal rx_output_fifo_N1589_FROM : STD_LOGIC; 
  signal rx_output_fifo_N3971 : STD_LOGIC; 
  signal rx_output_fifo_N3973 : STD_LOGIC; 
  signal rx_output_fifo_N3968 : STD_LOGIC; 
  signal rx_output_fifo_N3969 : STD_LOGIC; 
  signal mac_control_lmacaddr_15_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd6_In : STD_LOGIC; 
  signal tx_output_cs_FFd5_In : STD_LOGIC; 
  signal tx_output_cs_FFd8_In : STD_LOGIC; 
  signal tx_output_cs_FFd7_In : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_0_69_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_0_net34 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_0_69_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_1_68_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_1_net32 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_1_68_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_2_67_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_2_net30 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_2_67_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_3_66_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_3_net28 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_3_66_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_4_65_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_4_net26 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_4_65_CEMUXNOT : STD_LOGIC; 
  signal MD_6_ENABLE : STD_LOGIC; 
  signal MD_6_TORGTS : STD_LOGIC; 
  signal MD_6_OUTMUX : STD_LOGIC; 
  signal MD_6_OD : STD_LOGIC; 
  signal MD_7_ENABLE : STD_LOGIC; 
  signal MD_7_TORGTS : STD_LOGIC; 
  signal MD_7_OUTMUX : STD_LOGIC; 
  signal MD_7_OD : STD_LOGIC; 
  signal MD_8_ENABLE : STD_LOGIC; 
  signal MD_8_TORGTS : STD_LOGIC; 
  signal MD_8_OUTMUX : STD_LOGIC; 
  signal MD_8_OD : STD_LOGIC; 
  signal MD_9_ENABLE : STD_LOGIC; 
  signal MD_9_TORGTS : STD_LOGIC; 
  signal MD_9_OUTMUX : STD_LOGIC; 
  signal MD_9_OD : STD_LOGIC; 
  signal GTX_CLK_ENABLE : STD_LOGIC; 
  signal GTX_CLK_TORGTS : STD_LOGIC; 
  signal GTX_CLK_OUTMUX : STD_LOGIC; 
  signal clkio_dll_LOCKED : STD_LOGIC; 
  signal clkio_dll_CLKDV : STD_LOGIC; 
  signal clkio_dll_CLK2X180 : STD_LOGIC; 
  signal clkio_dll_CLK2X : STD_LOGIC; 
  signal clkio_dll_CLK270 : STD_LOGIC; 
  signal clkio_dll_CLK180 : STD_LOGIC; 
  signal clkio_dll_CLK90 : STD_LOGIC; 
  signal clk_dll_LOCKED : STD_LOGIC; 
  signal clk_dll_CLKDV : STD_LOGIC; 
  signal clk_dll_CLK2X180 : STD_LOGIC; 
  signal clk_dll_CLK2X : STD_LOGIC; 
  signal clk_dll_CLK270 : STD_LOGIC; 
  signal clk_dll_CLK180 : STD_LOGIC; 
  signal clkrx_dll_LOCKED : STD_LOGIC; 
  signal clkrx_dll_CLKDV : STD_LOGIC; 
  signal clkrx_dll_CLK2X180 : STD_LOGIC; 
  signal clkrx_dll_CLK2X : STD_LOGIC; 
  signal clkrx_dll_CLK270 : STD_LOGIC; 
  signal clkrx_dll_CLK180 : STD_LOGIC; 
  signal clkrx_dll_CLK90 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOB4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA3 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA2 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DOA0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIB4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_DIA4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_ADDRB1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_ADDRB0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_ADDRA1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_ADDRA0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_B11_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB3 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB2 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOB1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA3 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA2 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DOA0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIB4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_DIA4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_ADDRB1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_ADDRB0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_ADDRA1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_ADDRA0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_B15_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA3 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA2 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIB4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DIA4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRB1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRB0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRA1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRA0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA15 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA14 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA13 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA12 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA11 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA10 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA9 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA8 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA7 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA6 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA5 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA4 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA3 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA2 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA1 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA0 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRB3 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRB2 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRB1 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRB0 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRA3 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRA2 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRA1 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRA0 : STD_LOGIC; 
  signal rx_output_fifo_B7_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_B7_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_N82511 : STD_LOGIC; 
  signal mac_control_N82509 : STD_LOGIC; 
  signal mac_control_CHOICE1813_F5MUX : STD_LOGIC; 
  signal mac_control_N82501 : STD_LOGIC; 
  signal mac_control_N82499 : STD_LOGIC; 
  signal mac_control_CHOICE1869_F5MUX : STD_LOGIC; 
  signal mac_control_N82506 : STD_LOGIC; 
  signal mac_control_N82504 : STD_LOGIC; 
  signal mac_control_CHOICE1841_F5MUX : STD_LOGIC; 
  signal mac_control_N82496 : STD_LOGIC; 
  signal mac_control_N82494 : STD_LOGIC; 
  signal mac_control_CHOICE1897_F5MUX : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N82491 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N82489 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2588_F5MUX : STD_LOGIC; 
  signal memcontroller_N82421 : STD_LOGIC; 
  signal memcontroller_N82419 : STD_LOGIC; 
  signal memcontroller_addrn_10_F5MUX : STD_LOGIC; 
  signal memcontroller_N82426 : STD_LOGIC; 
  signal memcontroller_N82424 : STD_LOGIC; 
  signal memcontroller_addrn_11_F5MUX : STD_LOGIC; 
  signal memcontroller_N82431 : STD_LOGIC; 
  signal memcontroller_N82429 : STD_LOGIC; 
  signal memcontroller_addrn_12_F5MUX : STD_LOGIC; 
  signal memcontroller_N82436 : STD_LOGIC; 
  signal memcontroller_N82434 : STD_LOGIC; 
  signal memcontroller_addrn_13_F5MUX : STD_LOGIC; 
  signal memcontroller_N82441 : STD_LOGIC; 
  signal memcontroller_N82439 : STD_LOGIC; 
  signal memcontroller_addrn_14_F5MUX : STD_LOGIC; 
  signal memcontroller_N82446 : STD_LOGIC; 
  signal memcontroller_N82444 : STD_LOGIC; 
  signal memcontroller_addrn_15_F5MUX : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2401_FFY_RST : STD_LOGIC; 
  signal memcontroller_addrn_16_FROM : STD_LOGIC; 
  signal memcontroller_addrn_16_GROM : STD_LOGIC; 
  signal memcontroller_addrn_16_F5MUX : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15_FFX_RST : STD_LOGIC; 
  signal memcontroller_N82471 : STD_LOGIC; 
  signal memcontroller_N82469 : STD_LOGIC; 
  signal memcontroller_dnl1_3_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82476 : STD_LOGIC; 
  signal memcontroller_N82474 : STD_LOGIC; 
  signal memcontroller_dnl1_4_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82481 : STD_LOGIC; 
  signal memcontroller_N82479 : STD_LOGIC; 
  signal memcontroller_dnl1_5_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82331 : STD_LOGIC; 
  signal memcontroller_N82329 : STD_LOGIC; 
  signal memcontroller_dnl1_13_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82326 : STD_LOGIC; 
  signal memcontroller_N82324 : STD_LOGIC; 
  signal memcontroller_dnl1_14_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82486 : STD_LOGIC; 
  signal memcontroller_N82484 : STD_LOGIC; 
  signal memcontroller_dnl1_6_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82361 : STD_LOGIC; 
  signal memcontroller_N82359 : STD_LOGIC; 
  signal memcontroller_dnl1_7_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82321 : STD_LOGIC; 
  signal memcontroller_N82319 : STD_LOGIC; 
  signal memcontroller_dnl1_15_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82281 : STD_LOGIC; 
  signal memcontroller_N82279 : STD_LOGIC; 
  signal memcontroller_dnl1_23_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82456 : STD_LOGIC; 
  signal memcontroller_N82454 : STD_LOGIC; 
  signal memcontroller_dnl1_0_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82356 : STD_LOGIC; 
  signal memcontroller_N82354 : STD_LOGIC; 
  signal memcontroller_dnl1_8_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82316 : STD_LOGIC; 
  signal memcontroller_N82314 : STD_LOGIC; 
  signal memcontroller_dnl1_16_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82276 : STD_LOGIC; 
  signal memcontroller_N82274 : STD_LOGIC; 
  signal memcontroller_dnl1_24_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82461 : STD_LOGIC; 
  signal memcontroller_N82459 : STD_LOGIC; 
  signal memcontroller_dnl1_1_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82351 : STD_LOGIC; 
  signal memcontroller_N82349 : STD_LOGIC; 
  signal memcontroller_dnl1_9_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82311 : STD_LOGIC; 
  signal memcontroller_N82309 : STD_LOGIC; 
  signal memcontroller_dnl1_17_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82271 : STD_LOGIC; 
  signal memcontroller_N82269 : STD_LOGIC; 
  signal memcontroller_dnl1_25_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82466 : STD_LOGIC; 
  signal memcontroller_N82464 : STD_LOGIC; 
  signal memcontroller_dnl1_2_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82346 : STD_LOGIC; 
  signal memcontroller_N82344 : STD_LOGIC; 
  signal memcontroller_dnl1_10_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82306 : STD_LOGIC; 
  signal memcontroller_N82304 : STD_LOGIC; 
  signal memcontroller_dnl1_18_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82266 : STD_LOGIC; 
  signal memcontroller_N82264 : STD_LOGIC; 
  signal memcontroller_dnl1_26_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N17_FFY_RST : STD_LOGIC; 
  signal memcontroller_N82341 : STD_LOGIC; 
  signal memcontroller_N82339 : STD_LOGIC; 
  signal memcontroller_dnl1_11_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82301 : STD_LOGIC; 
  signal memcontroller_N82299 : STD_LOGIC; 
  signal memcontroller_dnl1_19_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82261 : STD_LOGIC; 
  signal memcontroller_N82259 : STD_LOGIC; 
  signal memcontroller_dnl1_27_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82336 : STD_LOGIC; 
  signal memcontroller_N82334 : STD_LOGIC; 
  signal memcontroller_dnl1_12_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82296 : STD_LOGIC; 
  signal memcontroller_N82294 : STD_LOGIC; 
  signal memcontroller_dnl1_20_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82251 : STD_LOGIC; 
  signal memcontroller_N82249 : STD_LOGIC; 
  signal memcontroller_dnl1_28_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82291 : STD_LOGIC; 
  signal memcontroller_N82289 : STD_LOGIC; 
  signal memcontroller_dnl1_21_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82246 : STD_LOGIC; 
  signal memcontroller_N82244 : STD_LOGIC; 
  signal memcontroller_dnl1_29_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82286 : STD_LOGIC; 
  signal memcontroller_N82284 : STD_LOGIC; 
  signal memcontroller_dnl1_22_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82256 : STD_LOGIC; 
  signal memcontroller_N82254 : STD_LOGIC; 
  signal memcontroller_dnl1_30_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2500_FFX_RST : STD_LOGIC; 
  signal memcontroller_N82451 : STD_LOGIC; 
  signal memcontroller_N82449 : STD_LOGIC; 
  signal memcontroller_dnl1_31_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N82371 : STD_LOGIC; 
  signal memcontroller_N82369 : STD_LOGIC; 
  signal memcontroller_addrn_0_F5MUX : STD_LOGIC; 
  signal memcontroller_N82381 : STD_LOGIC; 
  signal memcontroller_N82379 : STD_LOGIC; 
  signal memcontroller_addrn_2_F5MUX : STD_LOGIC; 
  signal memcontroller_N82386 : STD_LOGIC; 
  signal memcontroller_N82384 : STD_LOGIC; 
  signal memcontroller_addrn_3_F5MUX : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2401_FFX_RST : STD_LOGIC; 
  signal memcontroller_N82391 : STD_LOGIC; 
  signal memcontroller_N82389 : STD_LOGIC; 
  signal memcontroller_addrn_4_F5MUX : STD_LOGIC; 
  signal memcontroller_N82376 : STD_LOGIC; 
  signal memcontroller_N82374 : STD_LOGIC; 
  signal memcontroller_addrn_1_F5MUX : STD_LOGIC; 
  signal memcontroller_N82396 : STD_LOGIC; 
  signal memcontroller_N82394 : STD_LOGIC; 
  signal memcontroller_addrn_5_F5MUX : STD_LOGIC; 
  signal memcontroller_N82401 : STD_LOGIC; 
  signal memcontroller_N82399 : STD_LOGIC; 
  signal memcontroller_addrn_6_F5MUX : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2502_FFY_RST : STD_LOGIC; 
  signal memcontroller_N82406 : STD_LOGIC; 
  signal memcontroller_N82404 : STD_LOGIC; 
  signal memcontroller_addrn_7_F5MUX : STD_LOGIC; 
  signal memcontroller_N82411 : STD_LOGIC; 
  signal memcontroller_N82409 : STD_LOGIC; 
  signal memcontroller_addrn_8_F5MUX : STD_LOGIC; 
  signal memcontroller_N82416 : STD_LOGIC; 
  signal memcontroller_N82414 : STD_LOGIC; 
  signal memcontroller_addrn_9_F5MUX : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_lut2_0 : STD_LOGIC; 
  signal addr2ext_0_CYMUXG : STD_LOGIC; 
  signal addr2ext_0_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_0 : STD_LOGIC; 
  signal addr2ext_0_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_2_FROM : STD_LOGIC; 
  signal addr2ext_2_CYMUXG : STD_LOGIC; 
  signal addr2ext_2_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_2_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_2 : STD_LOGIC; 
  signal addr2ext_2_CYINIT : STD_LOGIC; 
  signal addr2ext_4_FROM : STD_LOGIC; 
  signal addr2ext_4_CYMUXG : STD_LOGIC; 
  signal addr2ext_4_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_4_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_4 : STD_LOGIC; 
  signal addr2ext_4_CYINIT : STD_LOGIC; 
  signal addr2ext_6_FROM : STD_LOGIC; 
  signal addr2ext_6_CYMUXG : STD_LOGIC; 
  signal addr2ext_6_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_6_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_6 : STD_LOGIC; 
  signal addr2ext_6_CYINIT : STD_LOGIC; 
  signal addr2ext_8_FROM : STD_LOGIC; 
  signal addr2ext_8_CYMUXG : STD_LOGIC; 
  signal addr2ext_8_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_8_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_8 : STD_LOGIC; 
  signal addr2ext_8_CYINIT : STD_LOGIC; 
  signal addr2ext_10_FROM : STD_LOGIC; 
  signal addr2ext_10_CYMUXG : STD_LOGIC; 
  signal addr2ext_10_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_10_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_10 : STD_LOGIC; 
  signal addr2ext_10_CYINIT : STD_LOGIC; 
  signal addr2ext_12_FROM : STD_LOGIC; 
  signal addr2ext_12_CYMUXG : STD_LOGIC; 
  signal addr2ext_12_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_12_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_12 : STD_LOGIC; 
  signal addr2ext_12_CYINIT : STD_LOGIC; 
  signal addr2ext_14_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_14_FROM : STD_LOGIC; 
  signal addr2ext_15_rt : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_14 : STD_LOGIC; 
  signal addr2ext_14_CYINIT : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_rt : STD_LOGIC; 
  signal rx_input_memio_bcnt_86_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_72 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_270 : STD_LOGIC; 
  signal rx_input_memio_bcnt_86_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_235 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_73 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_236 : STD_LOGIC; 
  signal rx_input_memio_bcnt_87_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_87_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_74 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_272 : STD_LOGIC; 
  signal rx_input_memio_bcnt_87_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_237 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_75 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_238 : STD_LOGIC; 
  signal rx_input_memio_bcnt_89_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_89_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_76 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_274 : STD_LOGIC; 
  signal rx_input_memio_bcnt_89_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_239 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_77 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_240 : STD_LOGIC; 
  signal rx_input_memio_bcnt_91_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_91_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_78 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_276 : STD_LOGIC; 
  signal rx_input_memio_bcnt_91_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_241 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_79 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_242 : STD_LOGIC; 
  signal rx_input_memio_bcnt_93_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_93_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_80 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_278 : STD_LOGIC; 
  signal rx_input_memio_bcnt_93_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_243 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_81 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_244 : STD_LOGIC; 
  signal rx_input_memio_bcnt_95_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_95_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_82 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_280 : STD_LOGIC; 
  signal rx_input_memio_bcnt_95_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_245 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_83 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_246 : STD_LOGIC; 
  signal rx_input_memio_bcnt_97_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_97_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_84 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_282 : STD_LOGIC; 
  signal rx_input_memio_bcnt_97_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_247 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_85 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_248 : STD_LOGIC; 
  signal rx_input_memio_bcnt_99_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_99_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_86 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_284 : STD_LOGIC; 
  signal rx_input_memio_bcnt_99_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_249 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_87 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_250 : STD_LOGIC; 
  signal rx_input_memio_bcnt_101_GROM : STD_LOGIC; 
  signal rx_input_memio_bcnt_101_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_lut2_48 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_49_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_lut2_49 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_48 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_49_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_2_FROM : STD_LOGIC; 
  signal rx_output_n0060_2_XORF : STD_LOGIC; 
  signal rx_output_n0060_2_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_2_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_2_XORG : STD_LOGIC; 
  signal rx_output_n0060_2_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_50 : STD_LOGIC; 
  signal rx_output_n0060_2_CYINIT : STD_LOGIC; 
  signal rx_output_n0060_4_FROM : STD_LOGIC; 
  signal rx_output_n0060_4_XORF : STD_LOGIC; 
  signal rx_output_n0060_4_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_4_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_4_XORG : STD_LOGIC; 
  signal rx_output_n0060_4_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_52 : STD_LOGIC; 
  signal rx_output_n0060_4_CYINIT : STD_LOGIC; 
  signal rx_output_n0060_6_FROM : STD_LOGIC; 
  signal rx_output_n0060_6_XORF : STD_LOGIC; 
  signal rx_output_n0060_6_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_6_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_6_XORG : STD_LOGIC; 
  signal rx_output_n0060_6_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_54 : STD_LOGIC; 
  signal rx_output_n0060_6_CYINIT : STD_LOGIC; 
  signal rx_output_n0060_8_FROM : STD_LOGIC; 
  signal rx_output_n0060_8_XORF : STD_LOGIC; 
  signal rx_output_n0060_8_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_8_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_8_XORG : STD_LOGIC; 
  signal rx_output_n0060_8_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_56 : STD_LOGIC; 
  signal rx_output_n0060_8_CYINIT : STD_LOGIC; 
  signal rx_output_n0060_10_FROM : STD_LOGIC; 
  signal rx_output_n0060_10_XORF : STD_LOGIC; 
  signal rx_output_n0060_10_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_10_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_10_XORG : STD_LOGIC; 
  signal rx_output_n0060_10_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_58 : STD_LOGIC; 
  signal rx_output_n0060_10_CYINIT : STD_LOGIC; 
  signal rx_output_n0060_12_FROM : STD_LOGIC; 
  signal rx_output_n0060_12_XORF : STD_LOGIC; 
  signal rx_output_n0060_12_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_12_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_12_XORG : STD_LOGIC; 
  signal rx_output_n0060_12_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_60 : STD_LOGIC; 
  signal rx_output_n0060_12_CYINIT : STD_LOGIC; 
  signal rx_output_n0060_14_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_14_FROM : STD_LOGIC; 
  signal rx_output_n0060_14_XORF : STD_LOGIC; 
  signal rx_output_n0060_14_XORG : STD_LOGIC; 
  signal rx_output_len_15_rt : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_62 : STD_LOGIC; 
  signal rx_output_n0060_14_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_4_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_4_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_10_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N17_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_31_rt : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_30_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_0_FROM : STD_LOGIC; 
  signal rx_input_memio_bp_0_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_134 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_221 : STD_LOGIC; 
  signal rx_input_memio_bp_0_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_0_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_bp_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_135 : STD_LOGIC; 
  signal rx_input_memio_bp_2_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_136 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_223 : STD_LOGIC; 
  signal rx_input_memio_bp_2_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2404_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bp_4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_137 : STD_LOGIC; 
  signal rx_input_memio_bp_4_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_138 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_225 : STD_LOGIC; 
  signal rx_input_memio_bp_4_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_6_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_139 : STD_LOGIC; 
  signal rx_input_memio_bp_6_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_140 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_227 : STD_LOGIC; 
  signal rx_input_memio_bp_6_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_8_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_141 : STD_LOGIC; 
  signal rx_input_memio_bp_8_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_142 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_229 : STD_LOGIC; 
  signal rx_input_memio_bp_8_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_10_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_143 : STD_LOGIC; 
  signal rx_input_memio_bp_10_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_144 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_231 : STD_LOGIC; 
  signal rx_input_memio_bp_10_CYINIT : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_145 : STD_LOGIC; 
  signal rx_input_memio_bp_12_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_146 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_233 : STD_LOGIC; 
  signal rx_input_memio_bp_12_CYINIT : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_147 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_148 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_235 : STD_LOGIC; 
  signal rx_input_memio_bp_14_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_4_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N19_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_24_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2502_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_31_rt : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_30_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_rst_rt : STD_LOGIC; 
  signal mac_control_ledrx_cnt_154_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_236 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_340 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_154_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_301 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_237 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_302 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_238 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_342 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_303 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_239 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_304 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_240 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_344 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_305 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_241 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_306 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_242 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_346 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_307 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_243 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_308 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_244 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_348 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_309 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_245 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_310 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_246 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_350 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_311 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_247 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_312 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_165_CYINIT : STD_LOGIC; 
  signal tx_output_bcntl_1_rt : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_195_CYMUXG : STD_LOGIC; 
  signal tx_output_SIG_25 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_194 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut1_6 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_197_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut1_7 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_196 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_197_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_197_CYINIT : STD_LOGIC; 
  signal tx_output_bcntl_3_rt : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_199_CYMUXG : STD_LOGIC; 
  signal tx_output_SIG_26 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_198 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_199_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_199_CYINIT : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut4_16 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_201_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut4_17 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_200 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_201_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_201_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2404_FFX_RST : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut4_18 : STD_LOGIC; 
  signal tx_output_n0035_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut4_19 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_202 : STD_LOGIC; 
  signal tx_output_n0035_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_n0035_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2504_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_14_CYINIT : STD_LOGIC; 
  signal MD_30_OFF_RST : STD_LOGIC; 
  signal MD_30_TFF_RST : STD_LOGIC; 
  signal MD_23_IFF_RST : STD_LOGIC; 
  signal MD_23_OFF_RST : STD_LOGIC; 
  signal MD_23_TFF_RST : STD_LOGIC; 
  signal MD_15_IFF_RST : STD_LOGIC; 
  signal MD_31_IFF_RST : STD_LOGIC; 
  signal MD_15_OFF_RST : STD_LOGIC; 
  signal MD_15_TFF_RST : STD_LOGIC; 
  signal DIN_3_IFF_RST : STD_LOGIC; 
  signal DIN_4_IFF_RST : STD_LOGIC; 
  signal DIN_5_IFF_RST : STD_LOGIC; 
  signal DIN_6_IFF_RST : STD_LOGIC; 
  signal DIN_7_IFF_RST : STD_LOGIC; 
  signal DIN_8_IFF_RST : STD_LOGIC; 
  signal DIN_9_IFF_RST : STD_LOGIC; 
  signal RX_ER_IFF_RST : STD_LOGIC; 
  signal RX_DV_IFF_RST : STD_LOGIC; 
  signal MA_10_OFF_RST : STD_LOGIC; 
  signal MD_26_OFF_RST : STD_LOGIC; 
  signal MD_26_TFF_RST : STD_LOGIC; 
  signal MD_19_IFF_RST : STD_LOGIC; 
  signal MD_19_OFF_RST : STD_LOGIC; 
  signal MD_19_TFF_RST : STD_LOGIC; 
  signal MD_27_IFF_RST : STD_LOGIC; 
  signal MD_28_IFF_RST : STD_LOGIC; 
  signal MD_27_OFF_RST : STD_LOGIC; 
  signal MD_27_TFF_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_31_rt : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_30_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_24_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N19_FFX_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_31_rt : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_30_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_16_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2406_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_31_rt : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_30_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_2_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_2_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_2_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_79 : STD_LOGIC; 
  signal rx_output_bp_0_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_80 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_86 : STD_LOGIC; 
  signal rx_output_bp_0_CYINIT : STD_LOGIC; 
  signal rx_output_bp_0_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_81 : STD_LOGIC; 
  signal rx_output_bp_2_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_82 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_88 : STD_LOGIC; 
  signal rx_output_bp_2_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_83 : STD_LOGIC; 
  signal rx_output_bp_4_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_84 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_90 : STD_LOGIC; 
  signal rx_output_bp_4_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_85 : STD_LOGIC; 
  signal rx_output_bp_6_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_86 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_92 : STD_LOGIC; 
  signal rx_output_bp_6_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_87 : STD_LOGIC; 
  signal rx_output_bp_8_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_88 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_94 : STD_LOGIC; 
  signal rx_output_bp_8_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_89 : STD_LOGIC; 
  signal rx_output_bp_10_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_90 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_96 : STD_LOGIC; 
  signal rx_output_bp_10_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_91 : STD_LOGIC; 
  signal rx_output_bp_12_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_92 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_98 : STD_LOGIC; 
  signal rx_output_bp_12_CYINIT : STD_LOGIC; 
  signal rx_output_bp_14_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_bp_14_FROM : STD_LOGIC; 
  signal rx_output_bp_15_rt : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_100 : STD_LOGIC; 
  signal rx_output_bp_14_CYINIT : STD_LOGIC; 
  signal tx_output_cs_FFd12_rt : STD_LOGIC; 
  signal tx_output_bcnt_38_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_40 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_204 : STD_LOGIC; 
  signal tx_output_bcnt_38_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_171 : STD_LOGIC; 
  signal tx_output_bcnt_39_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_41 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_172 : STD_LOGIC; 
  signal tx_output_bcnt_39_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_39_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_42 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_206 : STD_LOGIC; 
  signal tx_output_bcnt_39_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_173 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_43 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_174 : STD_LOGIC; 
  signal tx_output_bcnt_41_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_41_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_44 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_208 : STD_LOGIC; 
  signal tx_output_bcnt_41_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_175 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_45 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_176 : STD_LOGIC; 
  signal tx_output_bcnt_43_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_43_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_46 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_210 : STD_LOGIC; 
  signal tx_output_bcnt_43_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_177 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_47 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_178 : STD_LOGIC; 
  signal tx_output_bcnt_45_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_45_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_48 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_212 : STD_LOGIC; 
  signal tx_output_bcnt_45_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_179 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_49 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_180 : STD_LOGIC; 
  signal tx_output_bcnt_47_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_47_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_50 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_214 : STD_LOGIC; 
  signal tx_output_bcnt_47_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_181 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_51 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_182 : STD_LOGIC; 
  signal tx_output_bcnt_49_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_49_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_52 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_216 : STD_LOGIC; 
  signal tx_output_bcnt_49_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_183 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_53 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_184 : STD_LOGIC; 
  signal tx_output_bcnt_51_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_51_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_54 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_218 : STD_LOGIC; 
  signal tx_output_bcnt_51_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_185 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_55 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_186 : STD_LOGIC; 
  signal tx_output_bcnt_53_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2406_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_3_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_3_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_3_CYINIT : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_0 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_79_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_1 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_78 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_2 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_81_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_3 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_80 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_81_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_81_CYINIT : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_4 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_83_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_5 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_82 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_83_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_83_CYINIT : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_6 : STD_LOGIC; 
  signal rx_output_n0017_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_7 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_84 : STD_LOGIC; 
  signal rx_output_n0017_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0017_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_111 : STD_LOGIC; 
  signal rx_fifocheck_diff_0_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_112 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_161 : STD_LOGIC; 
  signal rx_fifocheck_diff_0_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_diff_0_LOGIC_ONE : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_113 : STD_LOGIC; 
  signal rx_fifocheck_diff_2_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_114 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_163 : STD_LOGIC; 
  signal rx_fifocheck_diff_2_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_115 : STD_LOGIC; 
  signal rx_fifocheck_diff_4_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_116 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_165 : STD_LOGIC; 
  signal rx_fifocheck_diff_4_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_117 : STD_LOGIC; 
  signal rx_fifocheck_diff_6_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_118 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_167 : STD_LOGIC; 
  signal rx_fifocheck_diff_6_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_119 : STD_LOGIC; 
  signal rx_fifocheck_diff_8_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_120 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_169 : STD_LOGIC; 
  signal rx_fifocheck_diff_8_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_121 : STD_LOGIC; 
  signal rx_fifocheck_diff_10_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_122 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_171 : STD_LOGIC; 
  signal rx_fifocheck_diff_10_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2505_FFY_SET : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_123 : STD_LOGIC; 
  signal rx_fifocheck_diff_12_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_124 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_173 : STD_LOGIC; 
  signal rx_fifocheck_diff_12_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_125 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_126 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_175 : STD_LOGIC; 
  signal rx_fifocheck_diff_14_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_111 : STD_LOGIC; 
  signal tx_fifocheck_diff_0_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_112 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_161 : STD_LOGIC; 
  signal tx_fifocheck_diff_0_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_0_LOGIC_ONE : STD_LOGIC; 
  signal tx_fifocheck_diff_2_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_113 : STD_LOGIC; 
  signal tx_fifocheck_diff_2_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_114 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_163 : STD_LOGIC; 
  signal tx_fifocheck_diff_2_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_4_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_115 : STD_LOGIC; 
  signal tx_fifocheck_diff_4_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_116 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_165 : STD_LOGIC; 
  signal tx_fifocheck_diff_4_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_6_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_117 : STD_LOGIC; 
  signal tx_fifocheck_diff_6_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_118 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_167 : STD_LOGIC; 
  signal tx_fifocheck_diff_6_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_8_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_119 : STD_LOGIC; 
  signal tx_fifocheck_diff_8_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_120 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_169 : STD_LOGIC; 
  signal tx_fifocheck_diff_8_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_10_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_121 : STD_LOGIC; 
  signal tx_fifocheck_diff_10_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_122 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_171 : STD_LOGIC; 
  signal tx_fifocheck_diff_10_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_12_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_123 : STD_LOGIC; 
  signal tx_fifocheck_diff_12_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_124 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_173 : STD_LOGIC; 
  signal tx_fifocheck_diff_12_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_14_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_125 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_126 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_175 : STD_LOGIC; 
  signal tx_fifocheck_diff_14_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_142_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_rst_rt : STD_LOGIC; 
  signal mac_control_ledtx_cnt_142_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_224 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_327 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_142_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_289 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_225 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_290 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_226 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_329 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_291 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_227 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_292 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_228 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_331 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_293 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_229 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_294 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_230 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_333 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_295 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_231 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_296 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_232 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_335 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_297 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_233 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_298 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_234 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_337 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_299 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_235 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_300 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_153_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N1912 : STD_LOGIC; 
  signal rx_output_fifo_N1904 : STD_LOGIC; 
  signal rx_output_fifo_N17_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N17_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1914 : STD_LOGIC; 
  signal rx_output_fifo_N17_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N17_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N1905 : STD_LOGIC; 
  signal rx_output_fifo_N15_FROM : STD_LOGIC; 
  signal rx_output_fifo_N1906 : STD_LOGIC; 
  signal rx_output_fifo_N15_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N15_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1924 : STD_LOGIC; 
  signal rx_output_fifo_N15_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N1907 : STD_LOGIC; 
  signal rx_output_fifo_N13_FROM : STD_LOGIC; 
  signal rx_output_fifo_N1908 : STD_LOGIC; 
  signal rx_output_fifo_N13_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N13_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1934 : STD_LOGIC; 
  signal rx_output_fifo_N13_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N1909 : STD_LOGIC; 
  signal rx_output_fifo_N11_FROM : STD_LOGIC; 
  signal rx_output_fifo_N1910 : STD_LOGIC; 
  signal rx_output_fifo_N10_rt : STD_LOGIC; 
  signal rx_output_fifo_N1944 : STD_LOGIC; 
  signal rx_output_fifo_N11_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N1911 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_95 : STD_LOGIC; 
  signal tx_input_n0074_0_XORF : STD_LOGIC; 
  signal tx_input_n0074_0_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_0_XORG : STD_LOGIC; 
  signal tx_input_n0074_0_GROM : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_118 : STD_LOGIC; 
  signal tx_input_n0074_0_CYINIT : STD_LOGIC; 
  signal tx_input_n0074_0_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_N21_FFX_RST : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_97 : STD_LOGIC; 
  signal tx_input_n0074_2_XORF : STD_LOGIC; 
  signal tx_input_n0074_2_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_2_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_98 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_120 : STD_LOGIC; 
  signal tx_input_n0074_2_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_99 : STD_LOGIC; 
  signal tx_input_n0074_4_XORF : STD_LOGIC; 
  signal tx_input_n0074_4_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_4_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_100 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_122 : STD_LOGIC; 
  signal tx_input_n0074_4_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_101 : STD_LOGIC; 
  signal tx_input_n0074_6_XORF : STD_LOGIC; 
  signal tx_input_n0074_6_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_6_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_102 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_124 : STD_LOGIC; 
  signal tx_input_n0074_6_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_103 : STD_LOGIC; 
  signal tx_input_n0074_8_XORF : STD_LOGIC; 
  signal tx_input_n0074_8_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_8_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_104 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_126 : STD_LOGIC; 
  signal tx_input_n0074_8_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_105 : STD_LOGIC; 
  signal tx_input_n0074_10_XORF : STD_LOGIC; 
  signal tx_input_n0074_10_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_10_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_106 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_128 : STD_LOGIC; 
  signal tx_input_n0074_10_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_107 : STD_LOGIC; 
  signal tx_input_n0074_12_XORF : STD_LOGIC; 
  signal tx_input_n0074_12_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_12_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_108 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_130 : STD_LOGIC; 
  signal tx_input_n0074_12_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_109 : STD_LOGIC; 
  signal tx_input_n0074_14_XORF : STD_LOGIC; 
  signal tx_input_n0074_14_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_110 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_132 : STD_LOGIC; 
  signal tx_input_n0074_14_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_1_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_1_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_1_CYINIT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd5_rt : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_32_CYMUXG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_34 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_187 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_32_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_165 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_35 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_166 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33_CYMUXG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_36 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_189 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33_CYINIT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_167 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_37 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_168 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35_CYMUXG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_38 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_191 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35_CYINIT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_169 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_39 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_170 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_37_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_37_CYINIT : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_0 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_79_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_1 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_78 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_2 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_81_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_3 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_80 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_81_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_81_CYINIT : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_4 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_83_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_5 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_82 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_83_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_83_CYINIT : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_6 : STD_LOGIC; 
  signal rx_output_n0018_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_7 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_84 : STD_LOGIC; 
  signal rx_output_n0018_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0018_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_txf_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_txf_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_txf_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_txf_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_txf_cnt_6_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_txf_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_txf_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_txf_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_txf_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_txf_cnt_16_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2505_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_txf_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_txf_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_txf_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_txf_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_txf_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_txf_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_31_rt : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_txf_cnt_30_CYINIT : STD_LOGIC; 
  signal rx_output_cs_FFd19_rt : STD_LOGIC; 
  signal addr3ext_0_CYMUXG : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_0 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_101 : STD_LOGIC; 
  signal addr3ext_0_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_95 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_1 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_96 : STD_LOGIC; 
  signal addr3ext_1_CYMUXG : STD_LOGIC; 
  signal addr3ext_1_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_2 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_103 : STD_LOGIC; 
  signal addr3ext_1_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_97 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_3 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_98 : STD_LOGIC; 
  signal addr3ext_3_CYMUXG : STD_LOGIC; 
  signal addr3ext_3_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_4 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_105 : STD_LOGIC; 
  signal addr3ext_3_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_99 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_5 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_100 : STD_LOGIC; 
  signal addr3ext_5_CYMUXG : STD_LOGIC; 
  signal addr3ext_5_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_6 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_107 : STD_LOGIC; 
  signal addr3ext_5_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_101 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_7 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_102 : STD_LOGIC; 
  signal addr3ext_7_CYMUXG : STD_LOGIC; 
  signal addr3ext_7_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_8 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_109 : STD_LOGIC; 
  signal addr3ext_7_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_103 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_9 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_104 : STD_LOGIC; 
  signal addr3ext_9_CYMUXG : STD_LOGIC; 
  signal addr3ext_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_10 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_111 : STD_LOGIC; 
  signal addr3ext_9_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_105 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_11 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_106 : STD_LOGIC; 
  signal addr3ext_11_CYMUXG : STD_LOGIC; 
  signal addr3ext_11_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_12 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_113 : STD_LOGIC; 
  signal addr3ext_11_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_107 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_13 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_108 : STD_LOGIC; 
  signal addr3ext_13_CYMUXG : STD_LOGIC; 
  signal addr3ext_13_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_14 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_115 : STD_LOGIC; 
  signal addr3ext_13_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_109 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_15 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_110 : STD_LOGIC; 
  signal addr3ext_15_GROM : STD_LOGIC; 
  signal addr3ext_15_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_diff_0_rt : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_SIG_27 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_151 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut4_8 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut4_9 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_153 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT : STD_LOGIC; 
  signal tx_input_dh_11_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut4_10 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut4_11 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_155 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_diff_13_rt : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_SIG_28 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_157 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_9_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut3_32 : STD_LOGIC; 
  signal rx_fifocheck_n0003_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut3_33 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_159 : STD_LOGIC; 
  signal rx_fifocheck_n0003_LOGIC_ONE : STD_LOGIC; 
  signal rx_fifocheck_n0003_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_0_rt : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_SIG_29 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_151 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut4_8 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut4_9 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_153 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut4_10 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut4_11 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_155 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_13_rt : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_SIG_30 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_157 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut3_32 : STD_LOGIC; 
  signal tx_fifocheck_n0003_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut3_33 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_159 : STD_LOGIC; 
  signal tx_fifocheck_n0003_LOGIC_ONE : STD_LOGIC; 
  signal tx_fifocheck_n0003_CYINIT : STD_LOGIC; 
  signal mac_control_N52153_rt : STD_LOGIC; 
  signal mac_control_phyrstcnt_110_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_192 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_294 : STD_LOGIC; 
  signal mac_control_phyrstcnt_110_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_257 : STD_LOGIC; 
  signal mac_control_phyrstcnt_111_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_193 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_258 : STD_LOGIC; 
  signal mac_control_phyrstcnt_111_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_111_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_194 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_296 : STD_LOGIC; 
  signal mac_control_phyrstcnt_111_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_259 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_195 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_260 : STD_LOGIC; 
  signal mac_control_phyrstcnt_113_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_113_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_196 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_298 : STD_LOGIC; 
  signal mac_control_phyrstcnt_113_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_261 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_197 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_262 : STD_LOGIC; 
  signal mac_control_phyrstcnt_115_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_115_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_198 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_300 : STD_LOGIC; 
  signal mac_control_phyrstcnt_115_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_263 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_199 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_264 : STD_LOGIC; 
  signal mac_control_phyrstcnt_117_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_117_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_200 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_302 : STD_LOGIC; 
  signal mac_control_phyrstcnt_117_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_265 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_201 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_266 : STD_LOGIC; 
  signal mac_control_phyrstcnt_119_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_119_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_202 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_304 : STD_LOGIC; 
  signal mac_control_phyrstcnt_119_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_267 : STD_LOGIC; 
  signal mac_control_phyrstcnt_121_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_203 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_268 : STD_LOGIC; 
  signal mac_control_phyrstcnt_121_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_121_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_204 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_306 : STD_LOGIC; 
  signal mac_control_phyrstcnt_121_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_269 : STD_LOGIC; 
  signal tx_input_dh_11_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_123_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_123_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_205 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_270 : STD_LOGIC; 
  signal mac_control_phyrstcnt_123_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_123_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_206 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_308 : STD_LOGIC; 
  signal mac_control_phyrstcnt_123_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_271 : STD_LOGIC; 
  signal mac_control_phyrstcnt_125_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_125_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_207 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_272 : STD_LOGIC; 
  signal mac_control_phyrstcnt_125_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_125_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_208 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_310 : STD_LOGIC; 
  signal mac_control_phyrstcnt_125_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_273 : STD_LOGIC; 
  signal mac_control_phyrstcnt_127_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_209 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_274 : STD_LOGIC; 
  signal mac_control_phyrstcnt_127_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_127_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_210 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_312 : STD_LOGIC; 
  signal mac_control_phyrstcnt_127_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_275 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_211 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_276 : STD_LOGIC; 
  signal mac_control_phyrstcnt_129_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_129_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_212 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_314 : STD_LOGIC; 
  signal mac_control_phyrstcnt_129_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_277 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_213 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_278 : STD_LOGIC; 
  signal mac_control_phyrstcnt_131_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_131_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_214 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_316 : STD_LOGIC; 
  signal mac_control_phyrstcnt_131_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_279 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_215 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_280 : STD_LOGIC; 
  signal mac_control_phyrstcnt_133_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_133_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_216 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_318 : STD_LOGIC; 
  signal mac_control_phyrstcnt_133_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_281 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_217 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_282 : STD_LOGIC; 
  signal mac_control_phyrstcnt_135_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_135_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_218 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_320 : STD_LOGIC; 
  signal mac_control_phyrstcnt_135_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_283 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_219 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_284 : STD_LOGIC; 
  signal mac_control_phyrstcnt_137_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_137_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_220 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_322 : STD_LOGIC; 
  signal mac_control_phyrstcnt_137_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_285 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_221 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_286 : STD_LOGIC; 
  signal mac_control_phyrstcnt_139_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_139_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_222 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_324 : STD_LOGIC; 
  signal mac_control_phyrstcnt_139_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_287 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_223 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_288 : STD_LOGIC; 
  signal mac_control_phyrstcnt_141_CYINIT : STD_LOGIC; 
  signal rx_input_memio_SIG_31 : STD_LOGIC; 
  signal rx_input_memio_macnt_70_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_56 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_253 : STD_LOGIC; 
  signal rx_input_memio_macnt_70_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_219 : STD_LOGIC; 
  signal tx_input_dh_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_57 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_220 : STD_LOGIC; 
  signal rx_input_memio_macnt_71_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_71_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_58 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_255 : STD_LOGIC; 
  signal rx_input_memio_macnt_71_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_221 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_59 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_222 : STD_LOGIC; 
  signal rx_input_memio_macnt_73_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_73_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_60 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_257 : STD_LOGIC; 
  signal rx_input_memio_macnt_73_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_223 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_61 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_224 : STD_LOGIC; 
  signal rx_input_memio_macnt_75_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_75_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_62 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_259 : STD_LOGIC; 
  signal rx_input_memio_macnt_75_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_225 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_63 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_226 : STD_LOGIC; 
  signal rx_input_memio_macnt_77_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_77_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_64 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_261 : STD_LOGIC; 
  signal rx_input_memio_macnt_77_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_227 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_65 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_228 : STD_LOGIC; 
  signal rx_input_memio_macnt_79_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_79_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_66 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_263 : STD_LOGIC; 
  signal rx_input_memio_macnt_79_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_229 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_67 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_230 : STD_LOGIC; 
  signal rx_input_memio_macnt_81_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_81_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_68 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_265 : STD_LOGIC; 
  signal rx_input_memio_macnt_81_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_231 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_69 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_232 : STD_LOGIC; 
  signal rx_input_memio_macnt_83_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_83_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_70 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_267 : STD_LOGIC; 
  signal rx_input_memio_macnt_83_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_233 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_71 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_234 : STD_LOGIC; 
  signal rx_input_memio_macnt_85_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_lut2_64 : STD_LOGIC; 
  signal rx_output_n0070_2_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_2_XORG : STD_LOGIC; 
  signal rx_output_n0070_2_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_63 : STD_LOGIC; 
  signal rx_output_n0070_2_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_3_FROM : STD_LOGIC; 
  signal rx_output_n0070_3_XORF : STD_LOGIC; 
  signal rx_output_n0070_3_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_3_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_3_XORG : STD_LOGIC; 
  signal rx_output_n0070_3_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_65 : STD_LOGIC; 
  signal rx_output_n0070_3_CYINIT : STD_LOGIC; 
  signal rx_output_n0070_5_FROM : STD_LOGIC; 
  signal rx_output_n0070_5_XORF : STD_LOGIC; 
  signal rx_output_n0070_5_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_5_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_5_XORG : STD_LOGIC; 
  signal rx_output_n0070_5_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_67 : STD_LOGIC; 
  signal rx_output_n0070_5_CYINIT : STD_LOGIC; 
  signal tx_input_dh_15_FFX_RST : STD_LOGIC; 
  signal rx_output_n0070_7_FROM : STD_LOGIC; 
  signal rx_output_n0070_7_XORF : STD_LOGIC; 
  signal rx_output_n0070_7_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_7_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_7_XORG : STD_LOGIC; 
  signal rx_output_n0070_7_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_69 : STD_LOGIC; 
  signal rx_output_n0070_7_CYINIT : STD_LOGIC; 
  signal rx_output_n0070_9_FROM : STD_LOGIC; 
  signal rx_output_n0070_9_XORF : STD_LOGIC; 
  signal rx_output_n0070_9_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_9_XORG : STD_LOGIC; 
  signal rx_output_n0070_9_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_71 : STD_LOGIC; 
  signal rx_output_n0070_9_CYINIT : STD_LOGIC; 
  signal rx_output_n0070_11_FROM : STD_LOGIC; 
  signal rx_output_n0070_11_XORF : STD_LOGIC; 
  signal rx_output_n0070_11_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_11_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_11_XORG : STD_LOGIC; 
  signal rx_output_n0070_11_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_73 : STD_LOGIC; 
  signal rx_output_n0070_11_CYINIT : STD_LOGIC; 
  signal rx_output_n0070_13_FROM : STD_LOGIC; 
  signal rx_output_n0070_13_XORF : STD_LOGIC; 
  signal rx_output_n0070_13_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_13_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_13_XORG : STD_LOGIC; 
  signal rx_output_n0070_13_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_75 : STD_LOGIC; 
  signal rx_output_n0070_13_CYINIT : STD_LOGIC; 
  signal rx_output_SIG_45 : STD_LOGIC; 
  signal rx_output_n0070_15_XORF : STD_LOGIC; 
  signal rx_output_n0070_15_CYINIT : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_0 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_79_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_1 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_78 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_2 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_81_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_3 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_80 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_81_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_81_CYINIT : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_4 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_83_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_5 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_82 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_83_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_83_CYINIT : STD_LOGIC; 
  signal rx_input_ince_FFX_RST : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_6 : STD_LOGIC; 
  signal tx_output_n0006_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_7 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_84 : STD_LOGIC; 
  signal tx_output_n0006_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_n0006_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_0_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_0_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_0_CYINIT : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_149 : STD_LOGIC; 
  signal rx_input_memio_bcntl_0_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_150 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_237 : STD_LOGIC; 
  signal rx_input_memio_bcntl_0_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_0_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_bcntl_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_2_FROM : STD_LOGIC; 
  signal rx_input_memio_bcntl_2_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_152 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_239 : STD_LOGIC; 
  signal rx_input_memio_bcntl_2_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_153 : STD_LOGIC; 
  signal rx_input_memio_bcntl_4_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_154 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_241 : STD_LOGIC; 
  signal rx_input_memio_bcntl_4_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_6_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_155 : STD_LOGIC; 
  signal rx_input_memio_bcntl_6_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_156 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_243 : STD_LOGIC; 
  signal rx_input_memio_bcntl_6_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_8_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_157 : STD_LOGIC; 
  signal rx_input_memio_bcntl_8_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_158 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_245 : STD_LOGIC; 
  signal rx_input_memio_bcntl_8_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_10_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_159 : STD_LOGIC; 
  signal rx_input_memio_bcntl_10_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_160 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_247 : STD_LOGIC; 
  signal rx_input_memio_bcntl_10_CYINIT : STD_LOGIC; 
  signal tx_input_dl_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_12_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_161 : STD_LOGIC; 
  signal rx_input_memio_bcntl_12_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_162 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_249 : STD_LOGIC; 
  signal rx_input_memio_bcntl_12_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_163 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_164 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_251 : STD_LOGIC; 
  signal rx_input_memio_bcntl_14_CYINIT : STD_LOGIC; 
  signal tx_input_addr_16_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd12_rt : STD_LOGIC; 
  signal tx_input_addr_16_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_16 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_134 : STD_LOGIC; 
  signal tx_input_addr_16_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_sum_127 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_17 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_128 : STD_LOGIC; 
  signal tx_input_addr_17_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_17_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_18 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_136 : STD_LOGIC; 
  signal tx_input_addr_17_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_129 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_19 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_130 : STD_LOGIC; 
  signal tx_input_addr_19_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_19_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_20 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_138 : STD_LOGIC; 
  signal tx_input_addr_19_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_131 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_21 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_132 : STD_LOGIC; 
  signal tx_input_addr_21_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_21_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_22 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_140 : STD_LOGIC; 
  signal tx_input_addr_21_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_133 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_23 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_134 : STD_LOGIC; 
  signal tx_input_addr_23_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_23_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_24 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_142 : STD_LOGIC; 
  signal tx_input_addr_23_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_135 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_25 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_136 : STD_LOGIC; 
  signal tx_input_addr_25_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_25_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_26 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_144 : STD_LOGIC; 
  signal tx_input_addr_25_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_137 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_27 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_138 : STD_LOGIC; 
  signal tx_input_addr_27_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_27_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_28 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_146 : STD_LOGIC; 
  signal tx_input_addr_27_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_139 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_29 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_140 : STD_LOGIC; 
  signal tx_input_addr_29_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_29_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_30 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_148 : STD_LOGIC; 
  signal tx_input_addr_29_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_141 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_31 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_142 : STD_LOGIC; 
  signal tx_input_addr_31_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_rxf_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_rxf_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_rxf_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_rxf_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_rxf_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_rxf_cnt_8_CYINIT : STD_LOGIC; 
  signal tx_input_dl_11_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_rxf_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_rxf_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_rxf_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_rxf_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_rxf_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_rxf_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_rxf_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_rxf_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_rxf_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_rxf_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_31_rt : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_rxf_cnt_30_CYINIT : STD_LOGIC; 
  signal txbp_11_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0078_inst_lut2_127 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_1_CYMUXG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_1_XORG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_1_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_181 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_1_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_2_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_2_XORF : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_2_CYMUXG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_2_XORG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_2_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_183 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_2_CYINIT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_4_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_4_XORF : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_4_XORG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_5_rt : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_185 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0078_4_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_5_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_5_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_5_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N2840 : STD_LOGIC; 
  signal rx_output_fifo_N2832 : STD_LOGIC; 
  signal rx_output_fifo_N9_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N9_GROM : STD_LOGIC; 
  signal rx_output_fifo_N2842 : STD_LOGIC; 
  signal rx_output_fifo_N9_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N2833 : STD_LOGIC; 
  signal rx_output_fifo_N7_FROM : STD_LOGIC; 
  signal rx_output_fifo_N2834 : STD_LOGIC; 
  signal rx_output_fifo_N7_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N7_GROM : STD_LOGIC; 
  signal rx_output_fifo_N2852 : STD_LOGIC; 
  signal rx_output_fifo_N7_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N2835 : STD_LOGIC; 
  signal rx_output_fifo_N5_FROM : STD_LOGIC; 
  signal rx_output_fifo_N2836 : STD_LOGIC; 
  signal rx_output_fifo_N5_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N5_GROM : STD_LOGIC; 
  signal rx_output_fifo_N2862 : STD_LOGIC; 
  signal rx_output_fifo_N5_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N2837 : STD_LOGIC; 
  signal rx_output_fifo_N3_FROM : STD_LOGIC; 
  signal rx_output_fifo_N2838 : STD_LOGIC; 
  signal rx_output_fifo_N2_rt : STD_LOGIC; 
  signal rx_output_fifo_N2872 : STD_LOGIC; 
  signal rx_output_fifo_N3_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N2839 : STD_LOGIC; 
  signal rx_output_fifo_N2569 : STD_LOGIC; 
  signal rx_output_fifo_N2576_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N2568 : STD_LOGIC; 
  signal rx_output_fifo_N2577 : STD_LOGIC; 
  signal rx_output_fifo_N2576_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N2576_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_fifo_N2567 : STD_LOGIC; 
  signal rx_output_fifo_N2574_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N2566 : STD_LOGIC; 
  signal rx_output_fifo_N2575 : STD_LOGIC; 
  signal rx_output_fifo_N2574_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N2574_CYINIT : STD_LOGIC; 
  signal tx_input_dl_13_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N2565 : STD_LOGIC; 
  signal rx_output_fifo_N2572_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N2564 : STD_LOGIC; 
  signal rx_output_fifo_N2573 : STD_LOGIC; 
  signal rx_output_fifo_N2572_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N2572_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N2563 : STD_LOGIC; 
  signal rx_output_fifo_BU172_O_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N2562 : STD_LOGIC; 
  signal rx_output_fifo_N2571 : STD_LOGIC; 
  signal rx_output_fifo_BU172_O_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_BU172_O_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_empty_FROM : STD_LOGIC; 
  signal rx_output_fifo_N2580 : STD_LOGIC; 
  signal rx_output_fifo_empty_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N3607 : STD_LOGIC; 
  signal rx_output_fifo_N3614_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N3606 : STD_LOGIC; 
  signal rx_output_fifo_N3615 : STD_LOGIC; 
  signal rx_output_fifo_N3614_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N3614_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_fifo_N3605 : STD_LOGIC; 
  signal rx_output_fifo_N3612_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N3604 : STD_LOGIC; 
  signal rx_output_fifo_N3613 : STD_LOGIC; 
  signal rx_output_fifo_N3612_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N3612_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N3603 : STD_LOGIC; 
  signal rx_output_fifo_N3610_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N3602 : STD_LOGIC; 
  signal rx_output_fifo_N3611 : STD_LOGIC; 
  signal rx_output_fifo_N3610_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N3610_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N3601 : STD_LOGIC; 
  signal rx_output_fifo_BU351_O_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N3600 : STD_LOGIC; 
  signal rx_output_fifo_N3609 : STD_LOGIC; 
  signal rx_output_fifo_BU351_O_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_BU351_O_CYINIT : STD_LOGIC; 
  signal tx_input_dl_15_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_full_FROM : STD_LOGIC; 
  signal rx_output_fifo_N3618 : STD_LOGIC; 
  signal rx_output_fifo_full_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N4756 : STD_LOGIC; 
  signal rx_output_fifo_N4763_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N4760 : STD_LOGIC; 
  signal rx_output_fifo_N4759 : STD_LOGIC; 
  signal rx_output_fifo_N4763_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_fifo_N4764 : STD_LOGIC; 
  signal rx_output_fifo_N4771_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N4768 : STD_LOGIC; 
  signal rx_output_fifo_N4767 : STD_LOGIC; 
  signal rx_output_fifo_N4771_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N4772 : STD_LOGIC; 
  signal rx_output_fifo_N4779_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N4776 : STD_LOGIC; 
  signal rx_output_fifo_N4775 : STD_LOGIC; 
  signal rx_output_fifo_N4779_CYINIT : STD_LOGIC; 
  signal txbp_13_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N4780 : STD_LOGIC; 
  signal rx_output_fifo_N4754 : STD_LOGIC; 
  signal rx_output_fifo_N4786 : STD_LOGIC; 
  signal rx_output_fifo_N4783 : STD_LOGIC; 
  signal rx_output_fifo_wrcount_0_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N4755 : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_103_rt : STD_LOGIC; 
  signal mac_control_bitcnt_104_CYMUXG : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_186 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_287 : STD_LOGIC; 
  signal mac_control_bitcnt_104_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_251 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_187 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_252 : STD_LOGIC; 
  signal mac_control_bitcnt_105_CYMUXG : STD_LOGIC; 
  signal mac_control_bitcnt_105_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_188 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_289 : STD_LOGIC; 
  signal mac_control_bitcnt_105_CYINIT : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_253 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_189 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_254 : STD_LOGIC; 
  signal mac_control_bitcnt_107_CYMUXG : STD_LOGIC; 
  signal mac_control_bitcnt_107_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_190 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_291 : STD_LOGIC; 
  signal mac_control_bitcnt_107_CYINIT : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_255 : STD_LOGIC; 
  signal tx_output_crcsell_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_n0063 : STD_LOGIC; 
  signal mac_control_n0064 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd4_In : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd3_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd10_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd9_In : STD_LOGIC; 
  signal tx_input_dl_15_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd3_In : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd5_In : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd4_In : STD_LOGIC; 
  signal txbp_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd12_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd11_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd14_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd13_In : STD_LOGIC; 
  signal mac_control_n0065 : STD_LOGIC; 
  signal mac_control_n0067 : STD_LOGIC; 
  signal rx_input_memio_menl_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_menl_FROM : STD_LOGIC; 
  signal rx_input_memio_menl_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxucastl_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_11_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_13_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_15_CEMUXNOT : STD_LOGIC; 
  signal tx_input_enableintl_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_enableintl_GSHIFT : STD_LOGIC; 
  signal tx_input_enableintl_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd2_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd1_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd4_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd3_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd6_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd5_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd8_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd7_In : STD_LOGIC; 
  signal tx_input_lden : STD_LOGIC; 
  signal tx_input_den_CEMUXNOT : STD_LOGIC; 
  signal rx_input_endfin_GROM : STD_LOGIC; 
  signal rx_output_fifo_N2259 : STD_LOGIC; 
  signal rx_output_fifo_N2299 : STD_LOGIC; 
  signal tx_output_crcenl_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcenl_FROM : STD_LOGIC; 
  signal tx_output_crcenl_GROM : STD_LOGIC; 
  signal mac_control_lsclkdelta : STD_LOGIC; 
  signal mac_control_lmacaddr_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_2_FROM : STD_LOGIC; 
  signal mac_control_n0068 : STD_LOGIC; 
  signal mac_control_n0066 : STD_LOGIC; 
  signal rx_output_fifodin_1_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_3_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_5_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_7_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_9_CEMUXNOT : STD_LOGIC; 
  signal rx_output_n0051 : STD_LOGIC; 
  signal rx_output_fifo_full_CEMUXNOT : STD_LOGIC; 
  signal rx_input_GMII_N80573 : STD_LOGIC; 
  signal rx_input_GMII_N80576 : STD_LOGIC; 
  signal rx_input_GMII_N80582 : STD_LOGIC; 
  signal rx_input_GMII_N80579 : STD_LOGIC; 
  signal mac_control_lmacaddr_21_FFX_RST : STD_LOGIC; 
  signal rx_input_GMII_N80561 : STD_LOGIC; 
  signal rx_input_GMII_N80570 : STD_LOGIC; 
  signal rx_input_GMII_N80567 : STD_LOGIC; 
  signal rx_input_GMII_N80564 : STD_LOGIC; 
  signal tx_input_dinint_11_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_11_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_13_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_13_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_15_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_15_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_n0061 : STD_LOGIC; 
  signal rx_input_memio_n0060 : STD_LOGIC; 
  signal rxfifowerr_CEMUXNOT : STD_LOGIC; 
  signal rx_output_cs_FFd17_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd17_In : STD_LOGIC; 
  signal rx_output_cs_FFd5_In : STD_LOGIC; 
  signal rx_output_cs_FFd19_In : STD_LOGIC; 
  signal rx_input_memio_n0058 : STD_LOGIC; 
  signal rx_input_memio_n0057 : STD_LOGIC; 
  signal rxoferr_CEMUXNOT : STD_LOGIC; 
  signal tx_input_cs_FFd11_FROM : STD_LOGIC; 
  signal tx_input_cs_FFd11_In : STD_LOGIC; 
  signal mac_control_lmacaddr_13_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_1_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_1_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_3_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_3_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_5_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_5_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_7_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_7_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_9_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_9_CEMUXNOT : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_net187 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_5_64_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_5_net24 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_5_64_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_6_63_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_6_net22 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_6_63_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_7_62_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_7_net20 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_7_62_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_8_61_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_8_net18 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_8_61_CEMUXNOT : STD_LOGIC; 
  signal mac_control_lmacaddr_33_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_9_60_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_9_net16 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_9_60_CEMUXNOT : STD_LOGIC; 
  signal tx_input_newfint_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_lnewfint : STD_LOGIC; 
  signal tx_input_newfint_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_22_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2197_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2197_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2277_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2277_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2021_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2021_GROM : STD_LOGIC; 
  signal mac_control_dout_11_FROM : STD_LOGIC; 
  signal mac_control_N79864 : STD_LOGIC; 
  signal mac_control_CHOICE2431_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2431_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2822_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2822_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2665_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2665_GROM : STD_LOGIC; 
  signal mac_control_lmacaddr_41_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE2869_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2869_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1942_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1942_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2322_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2322_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2366_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2366_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2673_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2673_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2833_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2833_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2606_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2606_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2290_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2290_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1939_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1939_GROM : STD_LOGIC; 
  signal mac_control_lmacaddr_17_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_20_FROM : STD_LOGIC; 
  signal mac_control_N74952 : STD_LOGIC; 
  signal mac_control_CHOICE2825_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2825_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2151_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2151_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2696_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2696_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2124_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2124_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2018_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2018_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2683_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2683_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2111_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2111_GROM : STD_LOGIC; 
  signal mac_control_lmacaddr_25_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE2704_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2704_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2618_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2618_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2637_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2637_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2385_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2385_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2057_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2057_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1965_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1965_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2114_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2114_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2614_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2614_GROM : STD_LOGIC; 
  signal mac_control_dout_12_FROM : STD_LOGIC; 
  signal mac_control_N78899 : STD_LOGIC; 
  signal mac_control_CHOICE2714_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2714_GROM : STD_LOGIC; 
  signal mac_control_dout_21_FROM : STD_LOGIC; 
  signal mac_control_N76020 : STD_LOGIC; 
  signal mac_control_lmacaddr_35_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE2391_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2391_GROM : STD_LOGIC; 
  signal mac_control_dout_30_FROM : STD_LOGIC; 
  signal mac_control_N75537 : STD_LOGIC; 
  signal mac_control_CHOICE1929_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1929_GROM : STD_LOGIC; 
  signal mac_control_dout_22_FROM : STD_LOGIC; 
  signal mac_control_N75069 : STD_LOGIC; 
  signal mac_control_CHOICE1998_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1998_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2044_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2044_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1926_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1926_GROM : STD_LOGIC; 
  signal mac_control_dout_15_FROM : STD_LOGIC; 
  signal mac_control_N80026 : STD_LOGIC; 
  signal mac_control_dout_13_FROM : STD_LOGIC; 
  signal mac_control_N79056 : STD_LOGIC; 
  signal mac_control_CHOICE2469_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2469_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1995_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1995_GROM : STD_LOGIC; 
  signal mac_control_lmacaddr_43_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_19_FROM : STD_LOGIC; 
  signal mac_control_dout_0_FROM : STD_LOGIC; 
  signal mac_control_N76337 : STD_LOGIC; 
  signal mac_control_CHOICE2309_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2309_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2103_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2103_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2233_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2233_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2901_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2901_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2175_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2175_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2347_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2347_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2216_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2216_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2135_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2135_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2649_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2649_GROM : STD_LOGIC; 
  signal mac_control_lmacaddr_19_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE1833_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1833_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1830_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1830_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2404_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2404_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2077_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2077_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1905_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1905_GROM : STD_LOGIC; 
  signal tx_output_crcl_13_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2127_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2127_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1988_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1988_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2138_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2138_GROM : STD_LOGIC; 
  signal mac_control_dout_16_FROM : STD_LOGIC; 
  signal mac_control_N75776 : STD_LOGIC; 
  signal mac_control_dout_24_FROM : STD_LOGIC; 
  signal mac_control_N76142 : STD_LOGIC; 
  signal mac_control_lmacaddr_27_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_25_FROM : STD_LOGIC; 
  signal mac_control_N75186 : STD_LOGIC; 
  signal mac_control_CHOICE2258_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2258_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2011_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2011_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1919_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1919_GROM : STD_LOGIC; 
  signal mac_control_dout_17_FROM : STD_LOGIC; 
  signal mac_control_N75898 : STD_LOGIC; 
  signal mac_control_dout_18_FROM : STD_LOGIC; 
  signal mac_control_N74835 : STD_LOGIC; 
  signal mac_control_dout_26_FROM : STD_LOGIC; 
  signal mac_control_N75303 : STD_LOGIC; 
  signal mac_control_CHOICE2296_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2296_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2246_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2246_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2034_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2034_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2360_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2360_GROM : STD_LOGIC; 
  signal mac_control_lmacaddr_37_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE1805_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1805_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1802_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1802_GROM : STD_LOGIC; 
  signal mac_control_dout_28_FROM : STD_LOGIC; 
  signal mac_control_N75420 : STD_LOGIC; 
  signal mac_control_CHOICE1889_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1889_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2080_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2080_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2087_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2087_GROM : STD_LOGIC; 
  signal mac_control_dout_29_FROM : STD_LOGIC; 
  signal mac_control_N75654 : STD_LOGIC; 
  signal mac_control_CHOICE2090_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2372_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2372_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_6_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2334_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2334_GROM : STD_LOGIC; 
  signal mac_control_lmacaddr_45_FFX_RST : STD_LOGIC; 
  signal tx_output_crcsell_3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_CHOICE2410_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2410_GROM : STD_LOGIC; 
  signal tx_input_cs_FFd5_FROM : STD_LOGIC; 
  signal tx_input_cs_FFd5_In : STD_LOGIC; 
  signal rx_input_RESET_1_FROM : STD_LOGIC; 
  signal rx_input_RESET_1_GROM : STD_LOGIC; 
  signal memcontroller_dnl2_1_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_3_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_5_CEMUXNOT : STD_LOGIC; 
  signal mac_control_lmacaddr_29_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_7_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_9_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcl_7_FROM : STD_LOGIC; 
  signal slowclock_rxcrcerrl_LOGIC_ZERO : STD_LOGIC; 
  signal slowclock_rxcrcerrl_GROM : STD_LOGIC; 
  signal mac_control_lmacaddr_39_FFX_RST : STD_LOGIC; 
  signal addr2ext_8_FFX_RST : STD_LOGIC; 
  signal addr2ext_10_FFX_RST : STD_LOGIC; 
  signal addr2ext_12_FFX_RST : STD_LOGIC; 
  signal addr2ext_14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_86_FFY_RST : STD_LOGIC; 
  signal addr2ext_4_FFX_RST : STD_LOGIC; 
  signal addr2ext_6_FFX_RST : STD_LOGIC; 
  signal addr2ext_8_FFY_RST : STD_LOGIC; 
  signal addr2ext_10_FFY_RST : STD_LOGIC; 
  signal addr2ext_12_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_95_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_97_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_99_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_101_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_99_FFX_RST : STD_LOGIC; 
  signal rxbp_15_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd10_In11_1_GROM : STD_LOGIC; 
  signal rx_output_invalid_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_3_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_5_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_7_CEMUXNOT : STD_LOGIC; 
  signal q2_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_9_CEMUXNOT : STD_LOGIC; 
  signal q2_1_FFX_RST : STD_LOGIC; 
  signal tx_output_ltxd_3_FROM : STD_LOGIC; 
  signal tx_output_ltxd_3_GROM : STD_LOGIC; 
  signal tx_output_ltxd_5_GROM : STD_LOGIC; 
  signal tx_output_crcl_17_FROM : STD_LOGIC; 
  signal rx_input_memio_crcl_12_FROM : STD_LOGIC; 
  signal rx_input_memio_dout_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_13_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_12_FFY_RST : STD_LOGIC; 
  signal q2_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_15_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_17_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_15_FFY_RST : STD_LOGIC; 
  signal q2_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_29_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpen_CEMUXNOT : STD_LOGIC; 
  signal q2_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_destok_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0053 : STD_LOGIC; 
  signal rx_input_memio_destok_CEMUXNOT : STD_LOGIC; 
  signal mac_control_n0033102_SW0_2_FROM : STD_LOGIC; 
  signal mac_control_n0033102_SW0_2_GROM : STD_LOGIC; 
  signal rx_output_cs_FFd10_FROM : STD_LOGIC; 
  signal rx_output_cs_FFd10_In : STD_LOGIC; 
  signal tx_output_crcl_18_FROM : STD_LOGIC; 
  signal tx_output_crcl_26_FROM : STD_LOGIC; 
  signal q3_1_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_8_FROM : STD_LOGIC; 
  signal mac_control_N77375 : STD_LOGIC; 
  signal rx_input_memio_crcl_19_FROM : STD_LOGIC; 
  signal slowclock_rxphyerrl_LOGIC_ZERO : STD_LOGIC; 
  signal slowclock_rxphyerrl_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_13_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2100_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2100_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2008_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2008_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1886_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1886_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2315_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2315_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2840_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2840_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1916_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1916_GROM : STD_LOGIC; 
  signal q2_7_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE2205_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2205_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2031_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2031_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2284_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2284_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2241_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2241_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2328_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2328_GROM : STD_LOGIC; 
  signal mac_control_dout_3_FROM : STD_LOGIC; 
  signal mac_control_N79540 : STD_LOGIC; 
  signal mac_control_CHOICE2279_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2279_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2603_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2603_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2805_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2805_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2611_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2611_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2808_GROM : STD_LOGIC; 
  signal q3_3_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE2621_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2621_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2398_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2398_GROM : STD_LOGIC; 
  signal mac_control_dout_4_FROM : STD_LOGIC; 
  signal mac_control_N78585 : STD_LOGIC; 
  signal mac_control_CHOICE2355_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2355_GROM : STD_LOGIC; 
  signal mac_control_dout_7_FROM : STD_LOGIC; 
  signal mac_control_N79702 : STD_LOGIC; 
  signal mac_control_CHOICE2317_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2317_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2837_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2837_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2842_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2634_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2634_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2393_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2393_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2642_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2642_GROM : STD_LOGIC; 
  signal q2_9_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE2652_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2652_GROM : STD_LOGIC; 
  signal mac_control_dout_9_FROM : STD_LOGIC; 
  signal mac_control_N78742 : STD_LOGIC; 
  signal tx_output_crcl_27_FROM : STD_LOGIC; 
  signal tx_input_cs_FFd12_FROM : STD_LOGIC; 
  signal tx_input_cs_FFd12_In : STD_LOGIC; 
  signal mac_control_N81741_GROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_18_42_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_18_42_1_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_11_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_21_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_13_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_13_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_31_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_23_CEMUXNOT : STD_LOGIC; 
  signal q3_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_15_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_41_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_41_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_33_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_33_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_25_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_17_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_43_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_43_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_35_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_27_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_19_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_45_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_45_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_37_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_37_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_29_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_47_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_47_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_39_CEMUXNOT : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_18_77_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_18_77_1_GROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_30_77_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_30_77_1_GROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_25_42_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_25_42_1_GROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_28_42_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_28_42_1_GROM : STD_LOGIC; 
  signal tx_output_crcl_28_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_25_77_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_25_77_1_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_23_FROM : STD_LOGIC; 
  signal rx_input_memio_crcl_15_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_16_80_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_16_80_1_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxallfl_CEMUXNOT : STD_LOGIC; 
  signal q3_7_FFX_RST : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_28_77_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_28_77_1_GROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_29_42_1_FROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_29_42_1_GROM : STD_LOGIC; 
  signal mac_control_n001220_SW0_1_GROM : STD_LOGIC; 
  signal mac_control_Mmux_n0017_Result_29_77_1_GROM : STD_LOGIC; 
  signal tx_output_crcl_29_FROM : STD_LOGIC; 
  signal rx_input_memio_crcll_11_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_13_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_21_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_15_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_31_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_23_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_17_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_25_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_27_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_19_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_29_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcl_24_FROM : STD_LOGIC; 
  signal rx_input_memio_crcl_16_FROM : STD_LOGIC; 
  signal mac_control_N52132_FROM : STD_LOGIC; 
  signal mac_control_N52132_GROM : STD_LOGIC; 
  signal q3_9_FFX_RST : STD_LOGIC; 
  signal mac_control_N52125_FROM : STD_LOGIC; 
  signal mac_control_N52125_GROM : STD_LOGIC; 
  signal mac_control_N52118_FROM : STD_LOGIC; 
  signal mac_control_N52118_GROM : STD_LOGIC; 
  signal mac_control_N52143_FROM : STD_LOGIC; 
  signal mac_control_N52143_GROM : STD_LOGIC; 
  signal mac_control_N52111_FROM : STD_LOGIC; 
  signal mac_control_N52111_GROM : STD_LOGIC; 
  signal mac_control_N52236_FROM : STD_LOGIC; 
  signal mac_control_N52236_GROM : STD_LOGIC; 
  signal mac_control_N52228_FROM : STD_LOGIC; 
  signal mac_control_N52228_GROM : STD_LOGIC; 
  signal mac_control_N52220_FROM : STD_LOGIC; 
  signal mac_control_N52220_GROM : STD_LOGIC; 
  signal mac_control_N52244_FROM : STD_LOGIC; 
  signal mac_control_N52244_GROM : STD_LOGIC; 
  signal mac_control_N52251_FROM : STD_LOGIC; 
  signal mac_control_N52251_GROM : STD_LOGIC; 
  signal mac_control_N52100_GROM : STD_LOGIC; 
  signal mac_control_N52268_FROM : STD_LOGIC; 
  signal mac_control_N52268_GROM : STD_LOGIC; 
  signal rxfbbp_15_FFX_RST : STD_LOGIC; 
  signal mac_control_N52198_GROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd3_FROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd3_In : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2564_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2564_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2574_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2574_GROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd4_FROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd4_In : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2591_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE2591_GROM : STD_LOGIC; 
  signal tx_output_bpl_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_3_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_7_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_9_CEMUXNOT : STD_LOGIC; 
  signal tx_output_N69282_FROM : STD_LOGIC; 
  signal tx_output_N69282_GROM : STD_LOGIC; 
  signal tx_output_bpl_11_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_13_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_addrl_3_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_addrl_4_FFY_RST : STD_LOGIC; 
  signal tx_input_CHOICE1722_FROM : STD_LOGIC; 
  signal tx_input_CHOICE1722_GROM : STD_LOGIC; 
  signal tx_input_CHOICE1702_GROM : STD_LOGIC; 
  signal tx_output_outsell_1_FROM : STD_LOGIC; 
  signal tx_output_outsel_1_Q : STD_LOGIC; 
  signal tx_output_outsell_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcl_17_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_n0019_SW0_2_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_n0019_SW0_2_GROM : STD_LOGIC; 
  signal tx_input_CHOICE1725_FROM : STD_LOGIC; 
  signal tx_input_CHOICE1725_GROM : STD_LOGIC; 
  signal tx_output_bpl_15_FFX_RST : STD_LOGIC; 
  signal memcontroller_oel_BYMUXNOT : STD_LOGIC; 
  signal memcontroller_oel_CEMUXNOT : STD_LOGIC; 
  signal slowclock_clkcnt_0_BXMUXNOT : STD_LOGIC; 
  signal rxoferrsr_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd6_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd6_In : STD_LOGIC; 
  signal rx_input_memio_crcl_18_FROM : STD_LOGIC; 
  signal rx_input_memio_crcl_26_FROM : STD_LOGIC; 
  signal memcontroller_clknum_0_BXMUXNOT : STD_LOGIC; 
  signal memcontroller_clknum_0_GROM : STD_LOGIC; 
  signal slowclock_rxfifowerrl_LOGIC_ZERO : STD_LOGIC; 
  signal slowclock_rxfifowerrl_GROM : STD_LOGIC; 
  signal txfbbp_1_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_3_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_5_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_7_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_9_CEMUXNOT : STD_LOGIC; 
  signal tx_output_outsell_2_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_9_rt : STD_LOGIC; 
  signal rx_input_fifo_control_d1_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_control_d0_9_rt : STD_LOGIC; 
  signal rx_input_fifo_control_d2_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_control_d1_9_rt : STD_LOGIC; 
  signal rx_input_memio_endbyte_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_control_d2_9_rt : STD_LOGIC; 
  signal rx_input_memio_crcl_27_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_miirw_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_miirw_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_cell_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcl_28_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_N41773_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_N41773_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_N41765_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_N41765_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_14_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_3_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_3_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_1_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_2_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_2_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_4_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_4_GROM : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1742_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_29_FROM : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1749_GROM : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1764_GROM : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1765_FROM : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1765_GROM : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1757_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_celll_CEMUXNOT : STD_LOGIC; 
  signal mac_control_addr_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_validmcast_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_CHOICE1570_GROM : STD_LOGIC; 
  signal mac_control_addr_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_rd_en_FROM : STD_LOGIC; 
  signal rx_input_fifo_rd_en_GROM : STD_LOGIC; 
  signal rx_input_fifo_rd_en_CEMUXNOT : STD_LOGIC; 
  signal rxfifofull_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxbcastl_CEMUXNOT : STD_LOGIC; 
  signal mac_control_addr_5_FFX_RST : STD_LOGIC; 
  signal rx_output_lenr_10_FROM : STD_LOGIC; 
  signal rx_output_lenr_10_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_11_FROM : STD_LOGIC; 
  signal rx_output_lenr_11_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_12_FROM : STD_LOGIC; 
  signal rx_output_lenr_12_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_13_FROM : STD_LOGIC; 
  signal rx_output_lenr_13_CEMUXNOT : STD_LOGIC; 
  signal mac_control_CHOICE2986_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2986_GROM : STD_LOGIC; 
  signal rx_output_lenr_14_FROM : STD_LOGIC; 
  signal rx_output_lenr_14_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_15_FROM : STD_LOGIC; 
  signal rx_output_lenr_15_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_14_FROM : STD_LOGIC; 
  signal mac_control_addr_7_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxmcastl_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_3_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_5_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_7_CEMUXNOT : STD_LOGIC; 
  signal tx_input_cs_FFd10_FFY_RST : STD_LOGIC; 
  signal mac_control_din_11_FFX_RST : STD_LOGIC; 
  signal mac_control_din_13_FFY_RST : STD_LOGIC; 
  signal mac_control_din_13_FFX_RST : STD_LOGIC; 
  signal mac_control_din_21_FFY_RST : STD_LOGIC; 
  signal mac_control_din_21_FFX_RST : STD_LOGIC; 
  signal mac_control_din_15_FFX_RST : STD_LOGIC; 
  signal mac_control_din_23_FFY_RST : STD_LOGIC; 
  signal mac_control_din_23_FFX_RST : STD_LOGIC; 
  signal mac_control_din_31_FFX_RST : STD_LOGIC; 
  signal mac_control_din_25_FFY_RST : STD_LOGIC; 
  signal mac_control_din_17_FFX_RST : STD_LOGIC; 
  signal rxfbbp_7_FFX_RST : STD_LOGIC; 
  signal rxfbbp_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_7_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_4_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_4_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_25_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_5_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_6_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_validbcast_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_7_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd12_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd14_FFX_RST : STD_LOGIC; 
  signal rx_output_ceinl_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd16_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cross_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd6_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_4_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_0_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_1_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd12_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd15_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd12_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd14_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd14_FFX_RST : STD_LOGIC; 
  signal mac_control_din_27_FFY_RST : STD_LOGIC; 
  signal mac_control_din_25_FFX_RST : STD_LOGIC; 
  signal mac_control_din_19_FFX_RST : STD_LOGIC; 
  signal mac_control_din_27_FFX_RST : STD_LOGIC; 
  signal mac_control_din_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd15_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_3_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_1_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_1_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_3_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_5_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_7_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_9_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_nearfull_FFY_RST : STD_LOGIC; 
  signal addr4ext_1_FFY_RST : STD_LOGIC; 
  signal addr4ext_1_FFX_RST : STD_LOGIC; 
  signal addr4ext_3_FFX_RST : STD_LOGIC; 
  signal addr4ext_5_FFX_RST : STD_LOGIC; 
  signal addr4ext_7_FFX_RST : STD_LOGIC; 
  signal d4_1_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_4_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_2_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_2_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_4_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_6_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_6_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_8_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_15_FFX_RST : STD_LOGIC; 
  signal rxf_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_1_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_1_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_3_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_5_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_7_FFX_RST : STD_LOGIC; 
  signal rxbp_3_FFX_RST : STD_LOGIC; 
  signal rxbp_5_FFX_RST : STD_LOGIC; 
  signal rxbp_7_FFX_RST : STD_LOGIC; 
  signal rxbp_9_FFX_RST : STD_LOGIC; 
  signal rxfbbp_1_FFX_RST : STD_LOGIC; 
  signal rxfbbp_3_FFX_RST : STD_LOGIC; 
  signal rxfbbp_7_FFY_RST : STD_LOGIC; 
  signal rxfbbp_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd8_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_5_FFX_RST : STD_LOGIC; 
  signal tx_input_dh_1_FFX_RST : STD_LOGIC; 
  signal tx_input_dh_3_FFX_RST : STD_LOGIC; 
  signal tx_input_dh_5_FFX_RST : STD_LOGIC; 
  signal tx_input_dh_7_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_7_FFX_RST : STD_LOGIC; 
  signal tx_input_dh_9_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_1_FFX_RST : STD_LOGIC; 
  signal txbp_1_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_1_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_1_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_3_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_5_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_7_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_13_FFX_RST : STD_LOGIC; 
  signal txbp_1_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_3_FFX_RST : STD_LOGIC; 
  signal txbp_3_FFY_RST : STD_LOGIC; 
  signal txbp_3_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_5_FFX_RST : STD_LOGIC; 
  signal txbp_5_FFY_RST : STD_LOGIC; 
  signal txbp_5_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_7_FFX_RST : STD_LOGIC; 
  signal txbp_7_FFY_RST : STD_LOGIC; 
  signal txbp_7_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_9_FFX_RST : STD_LOGIC; 
  signal txbp_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_5_FFX_RST : STD_LOGIC; 
  signal txfbbp_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_7_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_9_FFX_RST : STD_LOGIC; 
  signal rx_input_data_0_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd9_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_5_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_4_FFY_RST : STD_LOGIC; 
  signal tx_output_outsell_0_FFY_SET : STD_LOGIC; 
  signal mac_control_PHY_status_rwl_FFY_RST : STD_LOGIC; 
  signal rx_input_GMII_rx_of_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcrst_FFY_RST : STD_LOGIC; 
  signal mac_control_sclkll_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_1_FFX_RST : STD_LOGIC; 
  signal txfbbp_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_5_FFY_RST : STD_LOGIC; 
  signal txfbbp_13_FFX_RST : STD_LOGIC; 
  signal rx_input_data_1_FFY_RST : STD_LOGIC; 
  signal rx_input_data_2_FFY_RST : STD_LOGIC; 
  signal rx_input_data_3_FFY_RST : STD_LOGIC; 
  signal rx_input_data_4_FFY_RST : STD_LOGIC; 
  signal rx_input_data_5_FFY_RST : STD_LOGIC; 
  signal rx_input_data_6_FFY_RST : STD_LOGIC; 
  signal rx_input_data_7_FFY_RST : STD_LOGIC; 
  signal rx_input_endf_FFY_RST : STD_LOGIC; 
  signal rx_input_invalid_FFY_RST : STD_LOGIC; 
  signal tx_input_fifofulll_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcequal_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_10_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_phyaddrws_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_9_FFX_RST : STD_LOGIC; 
  signal rx_output_lenr_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_25_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cross_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_3_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1585_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_23_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_31_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_15_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_15_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1571_FFX_RST : STD_LOGIC; 
  signal q2_29_FFX_RST : STD_LOGIC; 
  signal q3_21_FFX_RST : STD_LOGIC; 
  signal q3_13_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1586_FFX_SET : STD_LOGIC; 
  signal addr4ext_9_FFX_RST : STD_LOGIC; 
  signal d4_1_FFX_RST : STD_LOGIC; 
  signal d4_3_FFX_RST : STD_LOGIC; 
  signal d4_5_FFX_RST : STD_LOGIC; 
  signal d4_7_FFX_RST : STD_LOGIC; 
  signal d4_9_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_11_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_13_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_15_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1605_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N1609_FFX_SET : STD_LOGIC; 
  signal mac_control_phystat_21_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_13_FFX_RST : STD_LOGIC; 
  signal q2_27_FFX_RST : STD_LOGIC; 
  signal q2_19_FFX_RST : STD_LOGIC; 
  signal q3_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_6_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_1_FFY_RST : STD_LOGIC; 
  signal macaddr_1_FFY_RST : STD_LOGIC; 
  signal macaddr_1_FFX_RST : STD_LOGIC; 
  signal macaddr_3_FFX_RST : STD_LOGIC; 
  signal macaddr_5_FFX_RST : STD_LOGIC; 
  signal macaddr_7_FFX_RST : STD_LOGIC; 
  signal macaddr_9_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_7_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_25_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_17_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_27_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_27_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_19_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_29_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd3_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_5_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_13_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_14_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_6_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_7_FFX_RST : STD_LOGIC; 
  signal MD_5_OFF_RST : STD_LOGIC; 
  signal MD_5_TFF_RST : STD_LOGIC; 
  signal MD_6_OFF_RST : STD_LOGIC; 
  signal MD_6_TFF_RST : STD_LOGIC; 
  signal MD_7_IFF_RST : STD_LOGIC; 
  signal MD_7_OFF_RST : STD_LOGIC; 
  signal MD_7_TFF_RST : STD_LOGIC; 
  signal MD_8_IFF_RST : STD_LOGIC; 
  signal MD_9_IFF_RST : STD_LOGIC; 
  signal MD_8_OFF_RST : STD_LOGIC; 
  signal MD_8_TFF_RST : STD_LOGIC; 
  signal MD_9_OFF_RST : STD_LOGIC; 
  signal MD_9_TFF_RST : STD_LOGIC; 
  signal addr2ext_0_FFY_RST : STD_LOGIC; 
  signal addr2ext_2_FFY_RST : STD_LOGIC; 
  signal addr2ext_6_FFY_RST : STD_LOGIC; 
  signal addr2ext_0_FFX_RST : STD_LOGIC; 
  signal addr2ext_2_FFX_RST : STD_LOGIC; 
  signal addr2ext_4_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_15_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_23_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_0_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_8_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_16_FFX_RST : STD_LOGIC; 
  signal rx_output_lenr_4_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_5_FFY_RST : STD_LOGIC; 
  signal rxbcast_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_14_FFY_RST : STD_LOGIC; 
  signal rx_output_bpl_5_FFX_RST : STD_LOGIC; 
  signal tx_output_datal_3_FFX_RST : STD_LOGIC; 
  signal rx_output_bpl_7_FFX_RST : STD_LOGIC; 
  signal tx_output_datal_5_FFX_RST : STD_LOGIC; 
  signal rx_output_bpl_9_FFX_RST : STD_LOGIC; 
  signal rx_output_bpl_9_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_7_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_8_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_10_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_10_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_0_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_1_FFY_RST : STD_LOGIC; 
  signal mac_control_bitcnt_109_FFX_RST : STD_LOGIC; 
  signal tx_input_DONE_FFY_RST : STD_LOGIC; 
  signal SOUT_OFF_RST : STD_LOGIC; 
  signal SCLK_IFF_RST : STD_LOGIC; 
  signal LEDRX_OFF_RST : STD_LOGIC; 
  signal LEDTX_OFF_RST : STD_LOGIC; 
  signal DIN_0_IFF_RST : STD_LOGIC; 
  signal DIN_1_IFF_RST : STD_LOGIC; 
  signal DIN_2_IFF_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_validucast_FFY_RST : STD_LOGIC; 
  signal rxmcast_FFY_RST : STD_LOGIC; 
  signal rxucast_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_30_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd7_FFX_SET : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd5_FFX_RST : STD_LOGIC; 
  signal tx_output_addrl_11_FFY_RST : STD_LOGIC; 
  signal tx_output_addrl_11_FFX_RST : STD_LOGIC; 
  signal tx_output_addrl_13_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_13_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_15_FFX_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_1_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_2_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_3_FFY_RST : STD_LOGIC; 
  signal tx_output_addrl_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_3_FFY_RST : STD_LOGIC; 
  signal txfifowerrsr_FFY_RST : STD_LOGIC; 
  signal tx_output_addrl_15_FFY_RST : STD_LOGIC; 
  signal tx_output_addrl_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_0_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_5_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_mcast_0_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_0_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_11_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_11_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_13_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_1_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_7_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_31_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_23_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_8_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_12_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_12_FFX_RST : STD_LOGIC; 
  signal tx_output_bcntl_14_FFX_RST : STD_LOGIC; 
  signal rx_output_bpl_11_FFY_RST : STD_LOGIC; 
  signal rx_output_bpl_11_FFX_RST : STD_LOGIC; 
  signal rx_output_bpl_13_FFX_RST : STD_LOGIC; 
  signal rx_output_bpl_15_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_1_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_30_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcen_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_7_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_11_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_13_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_15_FFX_RST : STD_LOGIC; 
  signal tx_output_ltxen3_FFY_RST : STD_LOGIC; 
  signal tx_output_ltxen3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_0_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_1_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_1_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_3_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_5_FFX_RST : STD_LOGIC; 
  signal q3_15_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1579_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1583_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1583_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_27_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_27_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_19_FFX_RST : STD_LOGIC; 
  signal q3_25_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_29_FFY_RST : STD_LOGIC; 
  signal q3_17_FFX_RST : STD_LOGIC; 
  signal memcontroller_oe_FFX_RST : STD_LOGIC; 
  signal MDIO_IFF_RST : STD_LOGIC; 
  signal DOUT_10_OFF_RST : STD_LOGIC; 
  signal rxcrcerrsr_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_27_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_19_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_rst_FFY_RST : STD_LOGIC; 
  signal q2_23_FFX_RST : STD_LOGIC; 
  signal q2_15_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1577_FFX_SET : STD_LOGIC; 
  signal mac_control_phystat_11_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1575_FFX_RST : STD_LOGIC; 
  signal q2_25_FFY_RST : STD_LOGIC; 
  signal q2_25_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1605_FFY_SET : STD_LOGIC; 
  signal q2_17_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1603_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N1607_FFX_SET : STD_LOGIC; 
  signal mac_control_phystat_25_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_17_FFX_RST : STD_LOGIC; 
  signal q3_31_FFX_RST : STD_LOGIC; 
  signal q3_23_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1546_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N1610_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N1563_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1567_FFX_RST : STD_LOGIC; 
  signal q2_11_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1627_FFX_RST : STD_LOGIC; 
  signal q2_11_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1569_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1565_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1569_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N1629_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1633_FFX_SET : STD_LOGIC; 
  signal q2_21_FFX_RST : STD_LOGIC; 
  signal q2_13_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1631_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1573_FFX_RST : STD_LOGIC; 
  signal q2_31_FFX_RST : STD_LOGIC; 
  signal q2_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_2_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_4_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_done_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_24_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_16_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_6_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_11_FFY_RST : STD_LOGIC; 
  signal tx_output_addrl_1_FFY_RST : STD_LOGIC; 
  signal tx_output_addrl_1_FFX_RST : STD_LOGIC; 
  signal tx_output_addrl_3_FFX_RST : STD_LOGIC; 
  signal tx_output_addrl_5_FFX_RST : STD_LOGIC; 
  signal tx_output_addrl_7_FFX_RST : STD_LOGIC; 
  signal rx_output_len_11_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_11_FFX_RST : STD_LOGIC; 
  signal tx_output_addrl_9_FFY_RST : STD_LOGIC; 
  signal DOUT_5_OFF_RST : STD_LOGIC; 
  signal DOUT_6_OFF_RST : STD_LOGIC; 
  signal DOUT_7_OFF_RST : STD_LOGIC; 
  signal DOUT_8_OFF_RST : STD_LOGIC; 
  signal DOUT_9_OFF_RST : STD_LOGIC; 
  signal rx_output_len_7_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_7_FFX_RST : STD_LOGIC; 
  signal rx_output_len_9_FFY_RST : STD_LOGIC; 
  signal rx_output_len_9_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_9_FFX_RST : STD_LOGIC; 
  signal tx_output_outselll_1_FFY_SET : STD_LOGIC; 
  signal tx_output_outselll_1_FFX_RST : STD_LOGIC; 
  signal tx_output_outselll_3_FFY_RST : STD_LOGIC; 
  signal tx_output_outselll_3_FFX_RST : STD_LOGIC; 
  signal tx_output_data_0_FFY_RST : STD_LOGIC; 
  signal tx_output_data_1_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_12_FFY_RST : STD_LOGIC; 
  signal tx_output_data_2_FFY_RST : STD_LOGIC; 
  signal tx_output_data_3_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_2_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd3_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd10_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd10_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_3_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_2_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_2_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_29_FFX_RST : STD_LOGIC; 
  signal q3_27_FFX_RST : STD_LOGIC; 
  signal q3_19_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1581_FFX_RST : STD_LOGIC; 
  signal q3_29_FFX_RST : STD_LOGIC; 
  signal rx_output_ceinll_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_10_FFY_RST : STD_LOGIC; 
  signal MD_28_OFF_RST : STD_LOGIC; 
  signal MD_28_TFF_RST : STD_LOGIC; 
  signal MD_29_IFF_RST : STD_LOGIC; 
  signal MD_29_OFF_RST : STD_LOGIC; 
  signal MD_29_TFF_RST : STD_LOGIC; 
  signal MA_0_OFF_RST : STD_LOGIC; 
  signal RXD_3_IFF_RST : STD_LOGIC; 
  signal RXD_4_IFF_RST : STD_LOGIC; 
  signal RXD_5_IFF_RST : STD_LOGIC; 
  signal RXD_6_IFF_RST : STD_LOGIC; 
  signal RXD_7_IFF_RST : STD_LOGIC; 
  signal DIN_10_IFF_RST : STD_LOGIC; 
  signal DIN_11_IFF_RST : STD_LOGIC; 
  signal DIN_12_IFF_RST : STD_LOGIC; 
  signal DIN_13_IFF_RST : STD_LOGIC; 
  signal DIN_14_IFF_RST : STD_LOGIC; 
  signal tx_output_data_4_FFY_RST : STD_LOGIC; 
  signal tx_output_data_5_FFY_RST : STD_LOGIC; 
  signal tx_output_data_6_FFY_RST : STD_LOGIC; 
  signal tx_output_data_7_FFY_RST : STD_LOGIC; 
  signal rx_output_denll_FFY_RST : STD_LOGIC; 
  signal rx_output_len_1_FFY_RST : STD_LOGIC; 
  signal rx_output_len_1_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_1_FFX_RST : STD_LOGIC; 
  signal rx_output_len_3_FFY_RST : STD_LOGIC; 
  signal rx_output_len_3_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_3_FFX_RST : STD_LOGIC; 
  signal rx_output_len_5_FFY_RST : STD_LOGIC; 
  signal rx_output_len_5_FFX_RST : STD_LOGIC; 
  signal rx_output_len_7_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_5_FFX_RST : STD_LOGIC; 
  signal tx_output_addrl_9_FFX_RST : STD_LOGIC; 
  signal rx_output_len_13_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_21_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_13_FFX_RST : STD_LOGIC; 
  signal rx_output_len_15_FFY_RST : STD_LOGIC; 
  signal rx_output_len_15_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_31_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_23_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_25_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_15_FFX_RST : STD_LOGIC; 
  signal DOUTEN_OFF_RST : STD_LOGIC; 
  signal MWE_OFF_SET : STD_LOGIC; 
  signal NEXTFRAME_IFF_RST : STD_LOGIC; 
  signal LEDACT_OFF_RST : STD_LOGIC; 
  signal TXD_0_OFF_RST : STD_LOGIC; 
  signal tx_output_bcntl_4_FFX_RST : STD_LOGIC; 
  signal tx_output_bcntl_6_FFX_RST : STD_LOGIC; 
  signal rx_output_bpl_1_FFX_RST : STD_LOGIC; 
  signal tx_output_bcntl_8_FFX_RST : STD_LOGIC; 
  signal rx_output_bpl_3_FFX_RST : STD_LOGIC; 
  signal tx_output_datal_1_FFX_RST : STD_LOGIC; 
  signal tx_output_bcntl_10_FFX_RST : STD_LOGIC; 
  signal LED100_OFF_RST : STD_LOGIC; 
  signal NEWFRAME_IFF_RST : STD_LOGIC; 
  signal LED1000_OFF_RST : STD_LOGIC; 
  signal TX_EN_OFF_RST : STD_LOGIC; 
  signal MD_13_OFF_RST : STD_LOGIC; 
  signal MD_13_TFF_RST : STD_LOGIC; 
  signal MD_22_IFF_RST : STD_LOGIC; 
  signal MD_22_OFF_RST : STD_LOGIC; 
  signal MD_22_TFF_RST : STD_LOGIC; 
  signal MD_14_IFF_RST : STD_LOGIC; 
  signal MD_30_IFF_RST : STD_LOGIC; 
  signal MD_14_OFF_RST : STD_LOGIC; 
  signal MD_14_TFF_RST : STD_LOGIC; 
  signal DOUT_11_OFF_RST : STD_LOGIC; 
  signal DOUT_12_OFF_RST : STD_LOGIC; 
  signal DOUT_13_OFF_RST : STD_LOGIC; 
  signal DOUT_14_OFF_RST : STD_LOGIC; 
  signal DOUT_15_OFF_RST : STD_LOGIC; 
  signal DIN_15_IFF_RST : STD_LOGIC; 
  signal DOUT_0_OFF_RST : STD_LOGIC; 
  signal DOUT_1_OFF_RST : STD_LOGIC; 
  signal DOUT_2_OFF_RST : STD_LOGIC; 
  signal DOUT_3_OFF_RST : STD_LOGIC; 
  signal DOUT_4_OFF_RST : STD_LOGIC; 
  signal MA_15_OFF_RST : STD_LOGIC; 
  signal MA_16_OFF_RST : STD_LOGIC; 
  signal MD_10_IFF_RST : STD_LOGIC; 
  signal MD_10_OFF_RST : STD_LOGIC; 
  signal MD_10_TFF_RST : STD_LOGIC; 
  signal MD_11_IFF_RST : STD_LOGIC; 
  signal MD_20_IFF_RST : STD_LOGIC; 
  signal MD_11_OFF_RST : STD_LOGIC; 
  signal MD_11_TFF_RST : STD_LOGIC; 
  signal TXD_1_OFF_RST : STD_LOGIC; 
  signal TXD_2_OFF_RST : STD_LOGIC; 
  signal TXD_3_OFF_RST : STD_LOGIC; 
  signal TXD_4_OFF_RST : STD_LOGIC; 
  signal TXD_5_OFF_RST : STD_LOGIC; 
  signal TXD_6_OFF_RST : STD_LOGIC; 
  signal TXD_7_OFF_RST : STD_LOGIC; 
  signal LEDDPX_OFF_RST : STD_LOGIC; 
  signal RXD_0_IFF_RST : STD_LOGIC; 
  signal RXD_1_IFF_RST : STD_LOGIC; 
  signal RXD_2_IFF_RST : STD_LOGIC; 
  signal MA_11_OFF_RST : STD_LOGIC; 
  signal MA_12_OFF_RST : STD_LOGIC; 
  signal MA_13_OFF_RST : STD_LOGIC; 
  signal MA_14_OFF_RST : STD_LOGIC; 
  signal MA_5_OFF_RST : STD_LOGIC; 
  signal MA_6_OFF_RST : STD_LOGIC; 
  signal MA_7_OFF_RST : STD_LOGIC; 
  signal MA_8_OFF_RST : STD_LOGIC; 
  signal MA_9_OFF_RST : STD_LOGIC; 
  signal PHYRESET_OFF_RST : STD_LOGIC; 
  signal memcontroller_dnl1_3_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_4_FFX_RST : STD_LOGIC; 
  signal MD_0_IFF_RST : STD_LOGIC; 
  signal MD_0_OFF_RST : STD_LOGIC; 
  signal MD_0_TFF_RST : STD_LOGIC; 
  signal MD_1_IFF_RST : STD_LOGIC; 
  signal MD_1_OFF_RST : STD_LOGIC; 
  signal MD_1_TFF_RST : STD_LOGIC; 
  signal MD_2_IFF_RST : STD_LOGIC; 
  signal MD_3_IFF_RST : STD_LOGIC; 
  signal MD_2_OFF_RST : STD_LOGIC; 
  signal MD_2_TFF_RST : STD_LOGIC; 
  signal MD_3_OFF_RST : STD_LOGIC; 
  signal MD_3_TFF_RST : STD_LOGIC; 
  signal MD_4_IFF_RST : STD_LOGIC; 
  signal MD_4_OFF_RST : STD_LOGIC; 
  signal MD_4_TFF_RST : STD_LOGIC; 
  signal MD_5_IFF_RST : STD_LOGIC; 
  signal MD_6_IFF_RST : STD_LOGIC; 
  signal MD_20_OFF_RST : STD_LOGIC; 
  signal MD_20_TFF_RST : STD_LOGIC; 
  signal MD_12_IFF_RST : STD_LOGIC; 
  signal MD_12_OFF_RST : STD_LOGIC; 
  signal MD_12_TFF_RST : STD_LOGIC; 
  signal MD_21_IFF_RST : STD_LOGIC; 
  signal MD_13_IFF_RST : STD_LOGIC; 
  signal MD_21_OFF_RST : STD_LOGIC; 
  signal MD_21_TFF_RST : STD_LOGIC; 
  signal MA_1_OFF_RST : STD_LOGIC; 
  signal MA_2_OFF_RST : STD_LOGIC; 
  signal MA_3_OFF_RST : STD_LOGIC; 
  signal MA_4_OFF_RST : STD_LOGIC; 
  signal mac_control_dout_28_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_29_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_31_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_23_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_15_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_15_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_25_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_25_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_17_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_17_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_27_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_27_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_19_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_19_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_datal_1_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_1_FFY_RST : STD_LOGIC; 
  signal rxphyerrsr_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_1_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_3_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_3_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_5_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_5_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_7_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_7_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_9_FFY_RST : STD_LOGIC; 
  signal mac_control_sclkdeltal_FFY_RST : STD_LOGIC; 
  signal addr2ext_14_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_87_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_87_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_89_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_91_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_2_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_10_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_18_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_26_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_11_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_24_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_1_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_9_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_17_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_89_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_91_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_93_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_93_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_95_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_97_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_21_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_29_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_22_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_30_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_0_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_2_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_4_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_19_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_27_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_12_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_20_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_28_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_0_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bp_10_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_12_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bp_14_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_165_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_6_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_12_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bp_8_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_154_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_8_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_10_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_12_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_12_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_14_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_14_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_38_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_2_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_4_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_6_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N13_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N11_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_0_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_2_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_0_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_4_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_49_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_51_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_51_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_53_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_14_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N17_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N17_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N15_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N11_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N15_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N13_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_0_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_2_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_4_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_8_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_4_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_6_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_2_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_4_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_6_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_10_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_6_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_8_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_111_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_113_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_117_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_113_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_115_FFY_RST : STD_LOGIC; 
  signal addr3ext_0_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_39_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_41_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_41_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_43_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_43_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_45_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_45_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_47_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_47_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_49_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_0_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_2_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_12_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_14_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_0_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_0_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_153_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_127_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_129_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_133_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_129_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_131_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_32_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_110_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_6_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_8_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_10_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_14_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_10_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_12_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_137_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_71_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_70_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_139_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_141_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_73_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_8_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_10_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_12_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_37_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_19_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_21_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_23_FFY_RST : STD_LOGIC; 
  signal tx_input_addr_27_FFY_RST : STD_LOGIC; 
  signal tx_input_addr_23_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_25_FFY_RST : STD_LOGIC; 
  signal addr3ext_3_FFX_RST : STD_LOGIC; 
  signal addr3ext_5_FFX_RST : STD_LOGIC; 
  signal addr3ext_7_FFY_RST : STD_LOGIC; 
  signal addr3ext_7_FFX_RST : STD_LOGIC; 
  signal addr3ext_9_FFY_RST : STD_LOGIC; 
  signal addr3ext_11_FFY_RST : STD_LOGIC; 
  signal addr3ext_1_FFY_RST : STD_LOGIC; 
  signal addr3ext_1_FFX_RST : STD_LOGIC; 
  signal addr3ext_3_FFY_RST : STD_LOGIC; 
  signal addr3ext_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_6_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_11_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_11_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_13_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_13_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_15_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_15_FFX_RST : STD_LOGIC; 
  signal tx_output_crcsell_3_FFY_RST : STD_LOGIC; 
  signal tx_output_crcsell_3_FFX_RST : STD_LOGIC; 
  signal tx_input_cs_FFd5_FFY_RST : STD_LOGIC; 
  signal addr3ext_9_FFX_RST : STD_LOGIC; 
  signal addr3ext_11_FFX_RST : STD_LOGIC; 
  signal addr3ext_13_FFY_RST : STD_LOGIC; 
  signal addr3ext_13_FFX_RST : STD_LOGIC; 
  signal addr3ext_15_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N7_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N5_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N3_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_7_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_9_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_115_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_117_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_119_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_119_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_121_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_131_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_133_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_135_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_139_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_135_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_137_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_0_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_0_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_71_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_73_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_75_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_79_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_75_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_77_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_2_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_4_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_6_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_83_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_85_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_25_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_27_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_29_FFY_RST : STD_LOGIC; 
  signal tx_input_addr_29_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_77_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_79_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_81_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_81_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_83_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_8_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_10_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_12_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_9_FFX_RST : STD_LOGIC; 
  signal rx_input_endfin_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1553_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1553_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_31_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_31_FFX_RST : STD_LOGIC; 
  signal mac_control_sclkdelta_FFY_RST : STD_LOGIC; 
  signal tx_output_crcenl_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_2_FFY_RST : STD_LOGIC; 
  signal tx_input_addr_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_14_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_21_FFY_RST : STD_LOGIC; 
  signal tx_input_addr_17_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_19_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_empty_FFX_SET : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd5_FFX_RST : STD_LOGIC; 
  signal addr1ext_7_FFX_RST : STD_LOGIC; 
  signal addr1ext_5_FFX_RST : STD_LOGIC; 
  signal addr1ext_7_FFY_RST : STD_LOGIC; 
  signal addr1ext_9_FFX_RST : STD_LOGIC; 
  signal addr1ext_9_FFY_RST : STD_LOGIC; 
  signal d1_1_FFX_RST : STD_LOGIC; 
  signal d1_1_FFY_RST : STD_LOGIC; 
  signal d1_3_FFX_RST : STD_LOGIC; 
  signal d1_3_FFY_RST : STD_LOGIC; 
  signal d1_5_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N9_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N9_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N7_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N5_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N3_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_3_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_5_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_5_FFX_RST : STD_LOGIC; 
  signal addr1ext_1_FFY_RST : STD_LOGIC; 
  signal addr1ext_1_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd3_FFY_RST : STD_LOGIC; 
  signal addr1ext_3_FFY_RST : STD_LOGIC; 
  signal addr1ext_3_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd5_FFY_RST : STD_LOGIC; 
  signal addr1ext_5_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_full_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_wrcount_0_FFY_RST : STD_LOGIC; 
  signal mac_control_bitcnt_104_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_wrcount_0_FFX_RST : STD_LOGIC; 
  signal mac_control_bitcnt_105_FFY_RST : STD_LOGIC; 
  signal tx_output_crcsell_1_FFY_SET : STD_LOGIC; 
  signal mac_control_bitcnt_105_FFX_RST : STD_LOGIC; 
  signal mac_control_bitcnt_107_FFY_RST : STD_LOGIC; 
  signal d1_23_FFX_RST : STD_LOGIC; 
  signal d1_15_FFX_RST : STD_LOGIC; 
  signal d1_25_FFX_RST : STD_LOGIC; 
  signal d1_25_FFY_RST : STD_LOGIC; 
  signal d1_17_FFY_RST : STD_LOGIC; 
  signal d1_17_FFX_RST : STD_LOGIC; 
  signal d1_27_FFY_RST : STD_LOGIC; 
  signal d1_27_FFX_RST : STD_LOGIC; 
  signal d1_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd12_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd14_FFX_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_rst_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_rst_FFX_RST : STD_LOGIC; 
  signal addr1ext_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_menl_FFX_RST : STD_LOGIC; 
  signal addr1ext_11_FFX_RST : STD_LOGIC; 
  signal addr1ext_13_FFX_RST : STD_LOGIC; 
  signal addr1ext_13_FFY_RST : STD_LOGIC; 
  signal addr1ext_15_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd4_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd6_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd8_FFX_SET : STD_LOGIC; 
  signal tx_output_crcsell_1_FFX_RST : STD_LOGIC; 
  signal mac_control_bitcnt_107_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_rst_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_rst_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd4_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd10_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd10_FFX_RST : STD_LOGIC; 
  signal tx_input_den_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_1_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_1_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_3_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_3_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_5_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_5_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_7_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_7_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_9_FFY_RST : STD_LOGIC; 
  signal d1_5_FFX_RST : STD_LOGIC; 
  signal d1_7_FFX_RST : STD_LOGIC; 
  signal d1_7_FFY_RST : STD_LOGIC; 
  signal d1_9_FFX_RST : STD_LOGIC; 
  signal d1_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd12_FFY_RST : STD_LOGIC; 
  signal d1_19_FFX_RST : STD_LOGIC; 
  signal d1_29_FFY_RST : STD_LOGIC; 
  signal d1_29_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_11_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_11_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_13_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_13_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_15_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_15_FFX_RST : STD_LOGIC; 
  signal tx_input_enableintl_FFY_RST : STD_LOGIC; 
  signal addr1ext_15_FFX_RST : STD_LOGIC; 
  signal d1_11_FFX_RST : STD_LOGIC; 
  signal d1_11_FFY_RST : STD_LOGIC; 
  signal d1_21_FFX_RST : STD_LOGIC; 
  signal d1_21_FFY_RST : STD_LOGIC; 
  signal d1_13_FFY_RST : STD_LOGIC; 
  signal d1_13_FFX_RST : STD_LOGIC; 
  signal d1_31_FFX_RST : STD_LOGIC; 
  signal d1_31_FFY_RST : STD_LOGIC; 
  signal d1_15_FFY_RST : STD_LOGIC; 
  signal d1_23_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_rst_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_rst_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_1_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_1_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_3_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_3_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_5_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_5_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_7_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_7_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_9_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_11_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_13_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_13_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_15_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_15_FFX_RST : STD_LOGIC; 
  signal rxfifowerr_FFY_RST : STD_LOGIC; 
  signal rxfifowerr_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd5_FFY_SET : STD_LOGIC; 
  signal tx_input_dinint_1_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_3_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_3_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_5_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_5_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_7_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_7_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_9_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_9_FFX_RST : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_103_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_11_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_11_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_21_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_21_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_13_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_13_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_31_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_23_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_9_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_full_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_11_FFY_RST : STD_LOGIC; 
  signal rxoferr_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd5_FFX_RST : STD_LOGIC; 
  signal rxoferr_FFX_RST : STD_LOGIC; 
  signal tx_input_cs_FFd11_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_11_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_11_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_13_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_13_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_15_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_15_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_1_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_19_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_0_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4_FFX_SET : STD_LOGIC; 
  signal rx_output_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd4_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1593_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1593_FFX_SET : STD_LOGIC; 
  signal tx_output_cs_FFd6_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd8_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_0_69_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_1_68_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_2_67_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_sclkdeltall_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_11_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_11_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_13_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_13_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_21_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_21_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_15_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_15_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_23_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_23_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_30_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_17_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd8_FFX_RST : STD_LOGIC; 
  signal tx_input_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal txfifowerr_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd4_FFX_RST : STD_LOGIC; 
  signal tx_input_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd8_FFX_RST : STD_LOGIC; 
  signal tx_input_cs_FFd9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_10_59_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_12_57_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_11_58_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_13_56_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_14_55_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_15_54_FFY_RST : STD_LOGIC; 
  signal mac_control_Mshreg_sinlll_102_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_31_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1551_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1615_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1549_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_3_66_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_4_65_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_5_64_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_6_63_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_7_62_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_8_61_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_9_60_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1549_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1615_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1617_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1617_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1613_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1613_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1589_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1588_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1589_FFX_SET : STD_LOGIC; 
  signal tx_output_crcl_21_FFY_RST : STD_LOGIC; 
  signal tx_input_newfint_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_21_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_22_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_11_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_17_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_25_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_25_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_19_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_19_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_27_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_27_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_29_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_13_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_31_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_13_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_12_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_23_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_15_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_12_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_1_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_1_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_3_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_3_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_1_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_5_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_3_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_7_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_5_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_9_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_16_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_24_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_25_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_17_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_18_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_26_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_20_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_5_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_5_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_7_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_7_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_21_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_30_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_22_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_15_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_13_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_13_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_19_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_27_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_27_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_29_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_7_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_11_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd6_FFY_SET : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_3_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_3_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_5_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_5_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_7_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_7_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd6_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_15_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_5_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_10_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_1_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_3_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_7_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_5_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_5_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_7_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_8_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_9_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_datal_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_datal_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_datal_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_datal_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_datal_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_datal_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_datal_7_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_0_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_0_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_23_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_41_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_33_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_33_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_41_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_17_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_35_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_27_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_9_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_7_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_9_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_7_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_9_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_12_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_11_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_11_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_13_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_13_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_15_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_7_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_9_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_23_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_41_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_33_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_17_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_43_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_35_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_35_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_43_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_43_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_37_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_37_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_45_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_45_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_39_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_39_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_47_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_47_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_7_FFY_RST : STD_LOGIC; 
  signal mac_control_lrxallf_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_doutl_7_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_8_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_wbpl_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_19_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_14_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_17_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_27_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_29_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_3_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_1_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_5_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_3_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_5_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_7_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_7_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_9_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpen_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_destok_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd10_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_18_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_26_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_3_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_35_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_27_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_45_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_37_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_39_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_47_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_13_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd12_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_23_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_17_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_27_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_39_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_28_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_24_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_16_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxallfl_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_1_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_1_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_3_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_3_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_5_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_7_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_5_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_7_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_9_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_9_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_13_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_29_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_5_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_7_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_8_FFY_RST : STD_LOGIC; 
  signal rxfsr_FFY_RST : STD_LOGIC; 
  signal txfsr_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_29_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_celll_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_rst_FFY_RST : STD_LOGIC; 
  signal macaddr_17_FFX_RST : STD_LOGIC; 
  signal macaddr_43_FFY_RST : STD_LOGIC; 
  signal macaddr_43_FFX_RST : STD_LOGIC; 
  signal macaddr_35_FFY_RST : STD_LOGIC; 
  signal macaddr_35_FFX_RST : STD_LOGIC; 
  signal macaddr_27_FFY_RST : STD_LOGIC; 
  signal macaddr_27_FFX_RST : STD_LOGIC; 
  signal macaddr_19_FFY_RST : STD_LOGIC; 
  signal macaddr_19_FFX_RST : STD_LOGIC; 
  signal macaddr_45_FFY_RST : STD_LOGIC; 
  signal macaddr_45_FFX_RST : STD_LOGIC; 
  signal macaddr_37_FFY_RST : STD_LOGIC; 
  signal macaddr_37_FFX_RST : STD_LOGIC; 
  signal macaddr_29_FFY_RST : STD_LOGIC; 
  signal macaddr_47_FFY_RST : STD_LOGIC; 
  signal macaddr_29_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_1_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_1_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_3_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_3_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_5_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_5_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_7_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_7_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_9_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_9_FFX_RST : STD_LOGIC; 
  signal macaddr_11_FFY_RST : STD_LOGIC; 
  signal macaddr_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal macaddr_11_FFX_RST : STD_LOGIC; 
  signal macaddr_21_FFX_RST : STD_LOGIC; 
  signal macaddr_13_FFY_RST : STD_LOGIC; 
  signal macaddr_13_FFX_RST : STD_LOGIC; 
  signal macaddr_31_FFY_RST : STD_LOGIC; 
  signal macaddr_31_FFX_RST : STD_LOGIC; 
  signal macaddr_23_FFY_RST : STD_LOGIC; 
  signal macaddr_23_FFX_RST : STD_LOGIC; 
  signal macaddr_15_FFY_RST : STD_LOGIC; 
  signal macaddr_15_FFX_RST : STD_LOGIC; 
  signal macaddr_41_FFY_RST : STD_LOGIC; 
  signal macaddr_41_FFX_RST : STD_LOGIC; 
  signal macaddr_33_FFY_RST : STD_LOGIC; 
  signal macaddr_33_FFX_RST : STD_LOGIC; 
  signal macaddr_25_FFY_RST : STD_LOGIC; 
  signal macaddr_17_FFY_RST : STD_LOGIC; 
  signal macaddr_25_FFX_RST : STD_LOGIC; 
  signal macaddr_47_FFX_RST : STD_LOGIC; 
  signal macaddr_39_FFY_RST : STD_LOGIC; 
  signal macaddr_39_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_addrl_1_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_addrl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_addrl_3_FFX_RST : STD_LOGIC; 
  signal tx_output_outsell_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_17_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_21_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_21_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_13_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_13_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_31_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_31_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_15_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_15_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_23_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_23_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_17_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_17_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_25_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_25_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_19_FFY_RST : STD_LOGIC; 
  signal mac_control_din_1_FFY_RST : STD_LOGIC; 
  signal mac_control_din_1_FFX_RST : STD_LOGIC; 
  signal mac_control_din_3_FFY_RST : STD_LOGIC; 
  signal mac_control_din_3_FFX_RST : STD_LOGIC; 
  signal mac_control_din_5_FFY_RST : STD_LOGIC; 
  signal mac_control_din_5_FFX_RST : STD_LOGIC; 
  signal mac_control_din_7_FFY_RST : STD_LOGIC; 
  signal mac_control_din_7_FFX_RST : STD_LOGIC; 
  signal mac_control_din_9_FFY_RST : STD_LOGIC; 
  signal mac_control_din_9_FFX_RST : STD_LOGIC; 
  signal memcontroller_oel_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_11_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_11_FFX_RST : STD_LOGIC; 
  signal txfbbp_1_FFX_RST : STD_LOGIC; 
  signal txfbbp_3_FFY_RST : STD_LOGIC; 
  signal txfbbp_3_FFX_RST : STD_LOGIC; 
  signal txfbbp_5_FFY_RST : STD_LOGIC; 
  signal txfbbp_5_FFX_RST : STD_LOGIC; 
  signal txfbbp_7_FFY_RST : STD_LOGIC; 
  signal txfbbp_7_FFX_RST : STD_LOGIC; 
  signal txfbbp_9_FFY_RST : STD_LOGIC; 
  signal txfbbp_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_11_FFX_RST : STD_LOGIC; 
  signal mac_control_lrxbcast_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_21_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_11_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_13_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_13_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_15_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_15_FFX_RST : STD_LOGIC; 
  signal rx_output_lenr_14_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_15_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxmcastl_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_13_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_23_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_17_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_27_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_19_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_11_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_13_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_13_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_15_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_18_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_26_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_0_FFY_RST : STD_LOGIC; 
  signal txfbbp_1_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_0_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_7_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_8_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_5_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_9_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_control_d2_9_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_7_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_9_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_control_d3_9_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_8_FFY_RST : STD_LOGIC; 
  signal d4_13_FFX_RST : STD_LOGIC; 
  signal d4_23_FFX_RST : STD_LOGIC; 
  signal d4_15_FFY_RST : STD_LOGIC; 
  signal d4_15_FFX_RST : STD_LOGIC; 
  signal d4_31_FFY_RST : STD_LOGIC; 
  signal d4_31_FFX_RST : STD_LOGIC; 
  signal d4_17_FFY_RST : STD_LOGIC; 
  signal d4_17_FFX_RST : STD_LOGIC; 
  signal d4_25_FFY_RST : STD_LOGIC; 
  signal d4_25_FFX_RST : STD_LOGIC; 
  signal d4_19_FFY_RST : STD_LOGIC; 
  signal d4_19_FFX_RST : STD_LOGIC; 
  signal d4_27_FFY_RST : STD_LOGIC; 
  signal d4_27_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_rd_en_FFY_RST : STD_LOGIC; 
  signal d4_29_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_5_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_9_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_control_d0_9_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_7_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_8_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_5_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_9_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_control_d1_9_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_27_FFY_RST : STD_LOGIC; 
  signal mac_control_lrxmcast_FFY_RST : STD_LOGIC; 
  signal rx_input_GMII_rx_dvll_FFY_RST : STD_LOGIC; 
  signal mac_control_lrxucast_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_cell_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_28_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_validmcast_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_rst_FFY_RST : STD_LOGIC; 
  signal addr4ext_11_FFY_RST : STD_LOGIC; 
  signal addr4ext_11_FFX_RST : STD_LOGIC; 
  signal addr4ext_13_FFY_RST : STD_LOGIC; 
  signal addr4ext_13_FFX_RST : STD_LOGIC; 
  signal addr4ext_15_FFY_RST : STD_LOGIC; 
  signal addr4ext_15_FFX_RST : STD_LOGIC; 
  signal d4_11_FFY_RST : STD_LOGIC; 
  signal d4_11_FFX_RST : STD_LOGIC; 
  signal rxallf_FFY_RST : STD_LOGIC; 
  signal d4_21_FFY_RST : STD_LOGIC; 
  signal d4_21_FFX_RST : STD_LOGIC; 
  signal d4_23_FFY_RST : STD_LOGIC; 
  signal d4_13_FFY_RST : STD_LOGIC; 
  signal d4_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxbcastl_FFY_RST : STD_LOGIC; 
  signal clkslen_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_10_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_11_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_12_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_11_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_13_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_5_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_7_FFX_RST : STD_LOGIC; 
  signal clkio_bufg_CE : STD_LOGIC; 
  signal clk_bufg_CE : STD_LOGIC; 
  signal clkrx_bufg_CE : STD_LOGIC; 
  signal PWR_VCC_0_FROM : STD_LOGIC; 
  signal PWR_VCC_0_GROM : STD_LOGIC; 
  signal PWR_VCC_1_FROM : STD_LOGIC; 
  signal PWR_VCC_1_GROM : STD_LOGIC; 
  signal PWR_VCC_2_FROM : STD_LOGIC; 
  signal PWR_VCC_2_GROM : STD_LOGIC; 
  signal PWR_VCC_3_FROM : STD_LOGIC; 
  signal PWR_VCC_3_GROM : STD_LOGIC; 
  signal PWR_VCC_4_FROM : STD_LOGIC; 
  signal PWR_VCC_4_GROM : STD_LOGIC; 
  signal PWR_VCC_5_FROM : STD_LOGIC; 
  signal PWR_VCC_6_FROM : STD_LOGIC; 
  signal PWR_VCC_7_FROM : STD_LOGIC; 
  signal PWR_VCC_8_FROM : STD_LOGIC; 
  signal PWR_VCC_8_GROM : STD_LOGIC; 
  signal PWR_VCC_9_FROM : STD_LOGIC; 
  signal PWR_VCC_9_GROM : STD_LOGIC; 
  signal PWR_VCC_10_FROM : STD_LOGIC; 
  signal PWR_VCC_10_GROM : STD_LOGIC; 
  signal PWR_VCC_11_FROM : STD_LOGIC; 
  signal PWR_VCC_11_GROM : STD_LOGIC; 
  signal PWR_VCC_12_FROM : STD_LOGIC; 
  signal PWR_VCC_12_GROM : STD_LOGIC; 
  signal PWR_VCC_13_FROM : STD_LOGIC; 
  signal PWR_VCC_13_GROM : STD_LOGIC; 
  signal PWR_VCC_14_FROM : STD_LOGIC; 
  signal PWR_VCC_14_GROM : STD_LOGIC; 
  signal PWR_VCC_15_FROM : STD_LOGIC; 
  signal PWR_VCC_15_GROM : STD_LOGIC; 
  signal PWR_VCC_16_FROM : STD_LOGIC; 
  signal PWR_VCC_16_GROM : STD_LOGIC; 
  signal PWR_VCC_17_FROM : STD_LOGIC; 
  signal PWR_VCC_17_GROM : STD_LOGIC; 
  signal PWR_VCC_18_FROM : STD_LOGIC; 
  signal PWR_VCC_18_GROM : STD_LOGIC; 
  signal PWR_VCC_19_FROM : STD_LOGIC; 
  signal PWR_VCC_19_GROM : STD_LOGIC; 
  signal PWR_VCC_20_FROM : STD_LOGIC; 
  signal PWR_VCC_21_FROM : STD_LOGIC; 
  signal PWR_VCC_22_FROM : STD_LOGIC; 
  signal PWR_VCC_22_GROM : STD_LOGIC; 
  signal PWR_VCC_23_FROM : STD_LOGIC; 
  signal PWR_VCC_24_FROM : STD_LOGIC; 
  signal PWR_VCC_24_GROM : STD_LOGIC; 
  signal PWR_VCC_25_FROM : STD_LOGIC; 
  signal PWR_VCC_26_FROM : STD_LOGIC; 
  signal PWR_VCC_26_GROM : STD_LOGIC; 
  signal PWR_VCC_27_FROM : STD_LOGIC; 
  signal PWR_VCC_27_GROM : STD_LOGIC; 
  signal PWR_VCC_28_FROM : STD_LOGIC; 
  signal PWR_VCC_29_FROM : STD_LOGIC; 
  signal PWR_VCC_29_GROM : STD_LOGIC; 
  signal PWR_VCC_30_FROM : STD_LOGIC; 
  signal PWR_VCC_30_GROM : STD_LOGIC; 
  signal PWR_VCC_31_FROM : STD_LOGIC; 
  signal PWR_VCC_31_GROM : STD_LOGIC; 
  signal PWR_VCC_32_FROM : STD_LOGIC; 
  signal PWR_VCC_32_GROM : STD_LOGIC; 
  signal PWR_VCC_33_FROM : STD_LOGIC; 
  signal PWR_VCC_34_FROM : STD_LOGIC; 
  signal PWR_VCC_34_GROM : STD_LOGIC; 
  signal PWR_VCC_35_FROM : STD_LOGIC; 
  signal PWR_VCC_35_GROM : STD_LOGIC; 
  signal PWR_VCC_36_FROM : STD_LOGIC; 
  signal PWR_VCC_36_GROM : STD_LOGIC; 
  signal PWR_VCC_37_FROM : STD_LOGIC; 
  signal PWR_VCC_37_GROM : STD_LOGIC; 
  signal PWR_VCC_38_FROM : STD_LOGIC; 
  signal PWR_VCC_38_GROM : STD_LOGIC; 
  signal PWR_GND_0_GROM : STD_LOGIC; 
  signal PWR_GND_1_GROM : STD_LOGIC; 
  signal PWR_GND_2_GROM : STD_LOGIC; 
  signal PWR_GND_3_GROM : STD_LOGIC; 
  signal PWR_GND_4_GROM : STD_LOGIC; 
  signal PWR_GND_5_GROM : STD_LOGIC; 
  signal PWR_GND_6_GROM : STD_LOGIC; 
  signal PWR_GND_7_GROM : STD_LOGIC; 
  signal PWR_GND_8_GROM : STD_LOGIC; 
  signal PWR_GND_9_GROM : STD_LOGIC; 
  signal PWR_GND_10_GROM : STD_LOGIC; 
  signal PWR_GND_11_GROM : STD_LOGIC; 
  signal PWR_GND_12_GROM : STD_LOGIC; 
  signal PWR_GND_13_GROM : STD_LOGIC; 
  signal PWR_GND_14_GROM : STD_LOGIC; 
  signal PWR_GND_15_GROM : STD_LOGIC; 
  signal PWR_GND_16_GROM : STD_LOGIC; 
  signal PWR_GND_17_GROM : STD_LOGIC; 
  signal PWR_GND_18_GROM : STD_LOGIC; 
  signal PWR_GND_19_GROM : STD_LOGIC; 
  signal PWR_GND_20_GROM : STD_LOGIC; 
  signal PWR_GND_21_GROM : STD_LOGIC; 
  signal PWR_GND_22_GROM : STD_LOGIC; 
  signal PWR_GND_23_GROM : STD_LOGIC; 
  signal PWR_GND_24_GROM : STD_LOGIC; 
  signal PWR_GND_25_GROM : STD_LOGIC; 
  signal PWR_GND_26_GROM : STD_LOGIC; 
  signal PWR_GND_27_GROM : STD_LOGIC; 
  signal PWR_GND_28_GROM : STD_LOGIC; 
  signal VCC : STD_LOGIC; 
  signal GND : STD_LOGIC; 
  signal rx_input_fifo_dout : STD_LOGIC_VECTOR ( 9 downto 9 ); 
  signal slowclock_clkcnt : STD_LOGIC_VECTOR ( 2 downto 0 ); 
  signal rx_input_fifo_fifodout : STD_LOGIC_VECTOR ( 8 downto 0 ); 
  signal rx_input_fifo_control_dinl : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal tx_input_dinint : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_input_dh : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_input_dl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal txbp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_din : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_lmacaddr : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal rxbp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal memcontroller_qn : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal q2 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal q3 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_output_bp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rxfbbp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_output_bpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_output_crcl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal tx_output_data : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal tx_output_outsell : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rx_input_data : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal rx_input_memio_endbyte : STD_LOGIC_VECTOR ( 2 downto 0 ); 
  signal mac_control_addr : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal tx_input_CNT : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_crcl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_datal : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal rx_input_memio_crccomb_n0118 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal rx_input_memio_crccomb_Mxor_n0007_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal mac_control_PHY_status_MII_Interface_statecnt : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal mac_control_PHY_status_miiaddr : STD_LOGIC_VECTOR ( 4 downto 0 ); 
  signal tx_output_crc_loigc_n0118 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal tx_output_crc_loigc_n0124 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal tx_output_crc_loigc_n0122 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal mac_control_PHY_status_MII_Interface_dreg : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_PHY_status_dout : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_PHY_status_din : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_bp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_bpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_phyaddr : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_dout : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal addr2ext : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal txfbbp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_fifo_control_d1 : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal rx_input_fifo_control_d0 : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal rx_input_fifo_control_d3 : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal rx_input_fifo_control_d2 : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_n0007_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_18_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_crc_loigc_n0115 : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_input_memio_crccomb_Mxor_CO_7_Xo : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal mac_control_PHY_status_MII_Interface_n0078 : STD_LOGIC_VECTOR ( 5 downto 1 ); 
  signal macaddr : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal rx_input_memio_crccomb_n0104 : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_input_memio_crccomb_n0115 : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_7_Xo : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal mac_control_phydi : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_rxfifowerr_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_crcll : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_dout : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_crccomb_Mxor_CO_26_Xo : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal rx_input_memio_crccomb_n0122 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal tx_output_crc_loigc_n0104 : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_9_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_output_fifo_wrcount : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal addr4ext : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal d4 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal tx_fifocheck_fbbpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_crccomb_n0124 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal rx_input_memio_addrchk_macaddrl : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal rx_output_len : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_output_n0070 : STD_LOGIC_VECTOR ( 15 downto 2 ); 
  signal rx_output_n0060 : STD_LOGIC_VECTOR ( 15 downto 2 ); 
  signal rx_output_lenr : STD_LOGIC_VECTOR ( 15 downto 2 ); 
  signal rx_input_memio_crccomb_Mxor_CO_9_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal memcontroller_clknum : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal rx_input_memio_addrchk_datal : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal rx_input_memio_addrchk_mcast : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_crcsell : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal tx_output_ncrcbytel : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal rx_input_memio_crccomb_n0056 : STD_LOGIC_VECTOR ( 2 downto 2 ); 
  signal rx_input_memio_addrchk_bcast : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal rx_input_memio_addrchk_maceq : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal rx_fifocheck_diff : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_output_crc_loigc_n0056 : STD_LOGIC_VECTOR ( 2 downto 2 ); 
  signal mac_control_phydo : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_phystat : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_txfifowerr_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_rxphyerr_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_rxoferr_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_rxcrcerr_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_txf_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_rxf_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal tx_output_addrl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_output_bcntl : STD_LOGIC_VECTOR ( 15 downto 1 ); 
  signal rx_output_bpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_output_mdl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal tx_output_datal : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_23_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_outselll : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal tx_output_ltxd : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_12_Xo : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal rx_output_fifodout : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_GMII_rxdl : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal tx_input_dinl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal memcontroller_addrn : STD_LOGIC_VECTOR ( 16 downto 0 ); 
  signal memcontroller_dnl2 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_fifoin : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal rx_output_fifodin : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal addr3ext : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal addr1ext : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal d1 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_dnl1 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_addrchk_lmaceq : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal rx_fifocheck_fbbpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_fifocheck_bpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_fifocheck_bpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_fifocheck_diff : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_input_n0074 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_bcntl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_doutl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_26_Xo : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal tx_output_crc_loigc_Mxor_CO_13_Xo : STD_LOGIC_VECTOR ( 2 downto 2 ); 
  signal rx_input_memio_crccomb_Mxor_CO_18_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_input_memio_crccomb_Mxor_CO_23_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_input_memio_crccomb_Mxor_CO_12_Xo : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal rx_input_memio_crccomb_Mxor_CO_13_Xo : STD_LOGIC_VECTOR ( 2 downto 2 ); 
  signal mac_control_PHY_status_addrl : STD_LOGIC_VECTOR ( 4 downto 0 ); 
  signal tx_output_n0034 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_n0048 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_fifo_control_ldata : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal mac_control_PHY_status_MII_Interface_n0014 : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal rx_output_n0046 : STD_LOGIC_VECTOR ( 15 downto 2 ); 
  signal rx_input_memio_addrchk_lmcast : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_ncrcbyte : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal memcontroller_ADDREXT : STD_LOGIC_VECTOR ( 16 downto 0 ); 
  signal rx_input_memio_addrchk_lbcast : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal tx_output_ldata : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal memcontroller_ts : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_dnout : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_q : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_dn : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal tx_output_addr_n0000 : STD_LOGIC_VECTOR ( 15 downto 1 ); 
  signal mac_control_rxcrcerr_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal rx_input_memio_n0043 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_rxoferr_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal mac_control_rxphyerr_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal mac_control_rxfifowerr_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal mac_control_txfifowerr_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal rx_output_lbp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_fifocheck_n0001 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_fifocheck_n0001 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_txf_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal rx_input_memio_n0042 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_rxf_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal tx_output_crcsel : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_input_memio_lma : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_lmd : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_output_lma : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal slowclock_clkcnt_n0000 : STD_LOGIC_VECTOR ( 2 downto 1 ); 
  signal tx_input_n0032 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_input_ldinint : STD_LOGIC_VECTOR ( 15 downto 0 ); 
begin
  rx_input_fifo_fifo_BU534 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2442,
      ADR1 => rx_input_fifo_fifo_N2443,
      ADR2 => rx_input_fifo_fifo_N2441,
      ADR3 => rx_input_fifo_fifo_N2444,
      O => rx_input_fifo_fifo_N5329_GROM
    );
  rx_input_fifo_fifo_N5329_YUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N5329_GROM,
      O => rx_input_fifo_fifo_N5329
    );
  rx_input_fifo_fifo_BU229 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_full,
      ADR2 => rx_input_ince,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2364_FROM
    );
  rx_input_fifo_fifo_BU235 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_full,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_ince,
      O => rx_input_fifo_fifo_N2364_GROM
    );
  rx_input_fifo_fifo_N2364_XUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2364_FROM,
      O => rx_input_fifo_fifo_N2364
    );
  rx_input_fifo_fifo_N2364_YUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2364_GROM,
      O => rx_input_fifo_fifo_N23
    );
  rx_input_fifo_fifo_full_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_full_FFX_SET
    );
  rx_input_fifo_fifo_BU435 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N4913,
      CE => rx_input_fifo_fifo_N4912,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_full_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_full
    );
  rx_input_fifo_fifo_BU434 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_full_CYINIT,
      I1 => rx_input_fifo_fifo_full_FROM,
      O => rx_input_fifo_fifo_N4913
    );
  rx_input_fifo_fifo_full_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_full_FROM
    );
  rx_input_fifo_fifo_full_CYINIT_4 : X_BUF
    port map (
      I => rx_input_fifo_fifo_BU431_O,
      O => rx_input_fifo_fifo_full_CYINIT
    );
  rx_input_fifo_fifo_N2427_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2427_FFY_SET
    );
  rx_input_fifo_fifo_BU429 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2417,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N2427_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2427
    );
  rx_input_fifo_fifo_N2427_LOGIC_ZERO_5 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N2427_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU428 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2427_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2427_CYINIT,
      SEL => rx_input_fifo_fifo_N4892,
      O => rx_input_fifo_fifo_N4902
    );
  rx_input_fifo_fifo_BU427 : X_LUT4
    generic map(
      INIT => X"99C3"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2418,
      ADR1 => rx_input_fifo_fifo_N2478,
      ADR2 => rx_input_fifo_fifo_N2428,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N4892
    );
  rx_input_fifo_fifo_BU430 : X_LUT4
    generic map(
      INIT => X"99C3"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2417,
      ADR1 => rx_input_fifo_fifo_N2477,
      ADR2 => rx_input_fifo_fifo_N2427,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N4891
    );
  rx_input_fifo_fifo_N2427_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2427_CYMUXG,
      O => rx_input_fifo_fifo_BU431_O
    );
  rx_input_fifo_fifo_BU431 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2427_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N4902,
      SEL => rx_input_fifo_fifo_N4891,
      O => rx_input_fifo_fifo_N2427_CYMUXG
    );
  rx_input_fifo_fifo_N2427_CYINIT_6 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4903,
      O => rx_input_fifo_fifo_N2427_CYINIT
    );
  rx_input_fifo_fifo_N2478_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2478_FFY_SET
    );
  rx_input_fifo_fifo_BU371 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N4730,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2478_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2477
    );
  rx_input_fifo_fifo_N2478_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2478_FFX_RST
    );
  rx_input_fifo_fifo_BU364 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N4690,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2478_FFX_RST,
      O => rx_input_fifo_fifo_N2478
    );
  rx_input_fifo_fifo_BU363 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N3,
      ADR1 => rx_input_fifo_fifo_N2,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4690
    );
  rx_input_fifo_fifo_BU370 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4730
    );
  rx_input_fifo_fifo_N3_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N3_FFX_RST
    );
  rx_input_fifo_fifo_BU294 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3943,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N3_FFX_RST,
      O => rx_input_fifo_fifo_N3
    );
  rx_input_fifo_fifo_N3_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N3_FFY_RST
    );
  rx_input_fifo_fifo_BU299 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3944,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N3_FFY_RST,
      O => rx_input_fifo_fifo_N2
    );
  rx_input_fifo_fifo_BU291 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N3,
      IB => rx_input_fifo_fifo_N3_CYINIT,
      SEL => rx_input_fifo_fifo_N3985,
      O => rx_input_fifo_fifo_N3987
    );
  rx_input_fifo_fifo_BU292 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N3_CYINIT,
      I1 => rx_input_fifo_fifo_N3985,
      O => rx_input_fifo_fifo_N3943
    );
  rx_input_fifo_fifo_BU290 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3985
    );
  rx_input_fifo_fifo_BU296 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3990
    );
  rx_input_fifo_fifo_BU297 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N3987,
      I1 => rx_input_fifo_fifo_N3990,
      O => rx_input_fifo_fifo_N3944
    );
  rx_input_fifo_fifo_N3_CYINIT_7 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3982,
      O => rx_input_fifo_fifo_N3_CYINIT
    );
  rx_input_fifo_fifo_N2417_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2417_FFX_SET
    );
  rx_input_fifo_fifo_BU394 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2397,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N2417_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2417
    );
  rx_input_fifo_fifo_N2417_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2417_FFY_RST
    );
  rx_input_fifo_fifo_BU392 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2398,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2417_FFY_RST,
      O => rx_input_fifo_fifo_N2418
    );
  rx_input_fifo_fifo_N2428_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2428_FFY_RST
    );
  rx_input_fifo_fifo_BU423 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2419,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2428_FFY_RST,
      O => rx_input_fifo_fifo_N2429
    );
  rx_input_fifo_fifo_N2428_LOGIC_ZERO_8 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N2428_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU422 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2428_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2428_CYINIT,
      SEL => rx_input_fifo_fifo_N4894,
      O => rx_input_fifo_fifo_N4904
    );
  rx_input_fifo_fifo_BU421 : X_LUT4
    generic map(
      INIT => X"A5C3"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2420,
      ADR1 => rx_input_fifo_fifo_N2430,
      ADR2 => rx_input_fifo_fifo_N2480,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N4894
    );
  rx_input_fifo_fifo_BU424 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2429,
      ADR1 => rx_input_fifo_fifo_N2479,
      ADR2 => rx_input_fifo_fifo_N2419,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N4893
    );
  rx_input_fifo_fifo_N2428_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2428_CYMUXG,
      O => rx_input_fifo_fifo_N4903
    );
  rx_input_fifo_fifo_BU425 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2428_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N4904,
      SEL => rx_input_fifo_fifo_N4893,
      O => rx_input_fifo_fifo_N2428_CYMUXG
    );
  rx_input_fifo_fifo_N2428_CYINIT_9 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4905,
      O => rx_input_fifo_fifo_N2428_CYINIT
    );
  rx_input_fifo_fifo_N2438_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2438_FFY_SET
    );
  rx_input_fifo_fifo_BU480 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2397,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2438_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2437
    );
  rx_input_fifo_fifo_N2467_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2467_FFY_SET
    );
  rx_input_fifo_fifo_BU456 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2467_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2468
    );
  rx_input_rx_nearf_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_rx_nearf_FFY_RST
    );
  rx_input_fifo_fifo_BU614 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N6323,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_rx_nearf_FFY_RST,
      O => rx_input_rx_nearf
    );
  rx_input_fifo_fifo_BU605 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2468,
      IB => rx_input_rx_nearf_CYINIT,
      SEL => rx_input_fifo_fifo_N6356,
      O => rx_input_fifo_fifo_N6359
    );
  rx_input_fifo_fifo_BU604 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2468,
      ADR1 => rx_input_fifo_fifo_N2448,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N6356
    );
  rx_input_fifo_fifo_BU610 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2467,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N2447,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N6362
    );
  rx_input_fifo_fifo_BU612 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N6359,
      I1 => rx_input_fifo_fifo_N6362,
      O => rx_input_fifo_fifo_N6323
    );
  rx_input_rx_nearf_CYINIT_10 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N6355,
      O => rx_input_rx_nearf_CYINIT
    );
  rx_input_fifo_fifo_BU498 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N2438,
      ADR2 => rx_input_fifo_fifo_N2437,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N5349
    );
  rx_input_fifo_fifo_BU349 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N5,
      ADR1 => rx_input_fifo_fifo_N4,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4610
    );
  rx_input_fifo_fifo_BU356 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N4,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N3,
      O => rx_input_fifo_fifo_N4650
    );
  rx_input_fifo_fifo_BU279 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N5,
      IB => rx_input_fifo_fifo_N5_CYINIT,
      SEL => rx_input_fifo_fifo_N3975,
      O => rx_input_fifo_fifo_N3977
    );
  rx_input_fifo_fifo_BU280 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N5_CYINIT,
      I1 => rx_input_fifo_fifo_N3975,
      O => rx_input_fifo_fifo_N3941
    );
  rx_input_fifo_fifo_BU278 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N5,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3975
    );
  rx_input_fifo_fifo_BU284 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N4,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3980
    );
  rx_input_fifo_fifo_N5_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N5_CYMUXG,
      O => rx_input_fifo_fifo_N3982
    );
  rx_input_fifo_fifo_BU285 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N4,
      IB => rx_input_fifo_fifo_N3977,
      SEL => rx_input_fifo_fifo_N3980,
      O => rx_input_fifo_fifo_N5_CYMUXG
    );
  rx_input_fifo_fifo_BU286 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N3977,
      I1 => rx_input_fifo_fifo_N3980,
      O => rx_input_fifo_fifo_N3942
    );
  rx_input_fifo_fifo_N5_CYINIT_11 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3972,
      O => rx_input_fifo_fifo_N5_CYINIT
    );
  rx_input_fifo_fifo_N2431_LOGIC_ZERO_12 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N2431_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU416 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2431_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2431_CYINIT,
      SEL => rx_input_fifo_fifo_N4896,
      O => rx_input_fifo_fifo_N4906
    );
  rx_input_fifo_fifo_BU415 : X_LUT4
    generic map(
      INIT => X"E12D"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2432,
      ADR1 => rx_input_fifo_fifo_full,
      ADR2 => rx_input_fifo_fifo_N2482,
      ADR3 => rx_input_fifo_fifo_N2422,
      O => rx_input_fifo_fifo_N4896
    );
  rx_input_fifo_fifo_BU418 : X_LUT4
    generic map(
      INIT => X"E12D"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2431,
      ADR1 => rx_input_fifo_fifo_full,
      ADR2 => rx_input_fifo_fifo_N2481,
      ADR3 => rx_input_fifo_fifo_N2421,
      O => rx_input_fifo_fifo_N4895
    );
  rx_input_fifo_fifo_N2431_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2431_CYMUXG,
      O => rx_input_fifo_fifo_N4905
    );
  rx_input_fifo_fifo_BU419 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2431_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N4906,
      SEL => rx_input_fifo_fifo_N4895,
      O => rx_input_fifo_fifo_N2431_CYMUXG
    );
  rx_input_fifo_fifo_N2431_CYINIT_13 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4907,
      O => rx_input_fifo_fifo_N2431_CYINIT
    );
  rx_input_fifo_fifo_N2469_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2469_FFY_SET
    );
  rx_input_fifo_fifo_BU452 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N5,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2469_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2470
    );
  rx_input_fifo_fifo_BU599 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2470,
      IB => rx_input_fifo_fifo_N6355_CYINIT,
      SEL => rx_input_fifo_fifo_N6348,
      O => rx_input_fifo_fifo_N6351
    );
  rx_input_fifo_fifo_BU598 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2470,
      ADR1 => rx_input_fifo_fifo_N2450,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N6348
    );
  rx_input_fifo_fifo_BU601 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2469,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N2449,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N6352
    );
  rx_input_fifo_fifo_N6355_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N6355_CYMUXG,
      O => rx_input_fifo_fifo_N6355
    );
  rx_input_fifo_fifo_BU602 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2469,
      IB => rx_input_fifo_fifo_N6351,
      SEL => rx_input_fifo_fifo_N6352,
      O => rx_input_fifo_fifo_N6355_CYMUXG
    );
  rx_input_fifo_fifo_N6355_CYINIT_14 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N6347,
      O => rx_input_fifo_fifo_N6355_CYINIT
    );
  rx_input_fifo_fifo_BU504 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2438,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N2439,
      ADR3 => rx_input_fifo_fifo_N2437,
      O => rx_input_fifo_fifo_N5348
    );
  rx_input_fifo_fifo_BU510 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2440,
      ADR1 => rx_input_fifo_fifo_N2438,
      ADR2 => rx_input_fifo_fifo_N2439,
      ADR3 => rx_input_fifo_fifo_N2437,
      O => rx_input_fifo_fifo_N2449_GROM
    );
  rx_input_fifo_fifo_N2449_YUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2449_GROM,
      O => rx_input_fifo_fifo_N5330
    );
  rx_input_fifo_fifo_BU426 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2418,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2428_FFX_RST,
      O => rx_input_fifo_fifo_N2428
    );
  rx_input_fifo_fifo_N2428_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2428_FFX_RST
    );
  rx_input_fifo_fifo_BU335 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N6,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N7,
      O => rx_input_fifo_fifo_N4530
    );
  rx_input_fifo_fifo_BU342 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N6,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N5,
      O => rx_input_fifo_fifo_N4570
    );
  rx_input_fifo_fifo_BU267 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N7,
      IB => rx_input_fifo_fifo_N7_CYINIT,
      SEL => rx_input_fifo_fifo_N3965,
      O => rx_input_fifo_fifo_N3967
    );
  rx_input_fifo_fifo_BU268 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N7_CYINIT,
      I1 => rx_input_fifo_fifo_N3965,
      O => rx_input_fifo_fifo_N3939
    );
  rx_input_fifo_fifo_BU266 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N7,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3965
    );
  rx_input_fifo_fifo_BU272 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N6,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3970
    );
  rx_input_fifo_fifo_N7_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N7_CYMUXG,
      O => rx_input_fifo_fifo_N3972
    );
  rx_input_fifo_fifo_BU273 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N6,
      IB => rx_input_fifo_fifo_N3967,
      SEL => rx_input_fifo_fifo_N3970,
      O => rx_input_fifo_fifo_N7_CYMUXG
    );
  rx_input_fifo_fifo_BU274 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N3967,
      I1 => rx_input_fifo_fifo_N3970,
      O => rx_input_fifo_fifo_N3940
    );
  rx_input_fifo_fifo_N7_CYINIT_15 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3962,
      O => rx_input_fifo_fifo_N7_CYINIT
    );
  rx_input_fifo_fifo_N2432_LOGIC_ZERO_16 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N2432_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU410 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2432_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2432_CYINIT,
      SEL => rx_input_fifo_fifo_N4898,
      O => rx_input_fifo_fifo_N4908
    );
  rx_input_fifo_fifo_BU409 : X_LUT4
    generic map(
      INIT => X"C3A5"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2434,
      ADR1 => rx_input_fifo_fifo_N2424,
      ADR2 => rx_input_fifo_fifo_N2484,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N4898
    );
  rx_input_fifo_fifo_BU412 : X_LUT4
    generic map(
      INIT => X"99C3"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2423,
      ADR1 => rx_input_fifo_fifo_N2483,
      ADR2 => rx_input_fifo_fifo_N2433,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N4897
    );
  rx_input_fifo_fifo_N2432_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2432_CYMUXG,
      O => rx_input_fifo_fifo_N4907
    );
  rx_input_fifo_fifo_BU413 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2432_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N4908,
      SEL => rx_input_fifo_fifo_N4897,
      O => rx_input_fifo_fifo_N2432_CYMUXG
    );
  rx_input_fifo_fifo_N2432_CYINIT_17 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4909,
      O => rx_input_fifo_fifo_N2432_CYINIT
    );
  rx_input_fifo_fifo_BU593 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2472,
      IB => rx_input_fifo_fifo_N6347_CYINIT,
      SEL => rx_input_fifo_fifo_N6340,
      O => rx_input_fifo_fifo_N6343
    );
  rx_input_fifo_fifo_BU592 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2472,
      ADR1 => rx_input_fifo_fifo_N2452,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N6340
    );
  rx_input_fifo_fifo_BU595 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2471,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N2451,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N6344
    );
  rx_input_fifo_fifo_N6347_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N6347_CYMUXG,
      O => rx_input_fifo_fifo_N6347
    );
  rx_input_fifo_fifo_BU596 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2471,
      IB => rx_input_fifo_fifo_N6343,
      SEL => rx_input_fifo_fifo_N6344,
      O => rx_input_fifo_fifo_N6347_CYMUXG
    );
  rx_input_fifo_fifo_N6347_CYINIT_18 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N6339,
      O => rx_input_fifo_fifo_N6347_CYINIT
    );
  rx_input_fifo_fifo_BU516 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N2441,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N5330,
      O => rx_input_fifo_fifo_N5346
    );
  rx_input_fifo_fifo_BU522 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N5330,
      ADR1 => rx_input_fifo_fifo_N2441,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N2442,
      O => rx_input_fifo_fifo_N5345
    );
  rx_input_fifo_fifo_BU328 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N8,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N7,
      O => rx_input_fifo_fifo_N4490
    );
  rx_input_fifo_fifo_BU321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N8,
      ADR2 => rx_input_fifo_fifo_N9,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4450
    );
  rx_input_fifo_fifo_BU255 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N9,
      IB => rx_input_fifo_fifo_N9_CYINIT,
      SEL => rx_input_fifo_fifo_N3955,
      O => rx_input_fifo_fifo_N3957
    );
  rx_input_fifo_fifo_BU256 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N9_CYINIT,
      I1 => rx_input_fifo_fifo_N3955,
      O => rx_input_fifo_fifo_N3937
    );
  rx_input_fifo_fifo_BU254 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N9,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3955
    );
  rx_input_fifo_fifo_BU260 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N8,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3960
    );
  rx_input_fifo_fifo_N9_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N9_CYMUXG,
      O => rx_input_fifo_fifo_N3962
    );
  rx_input_fifo_fifo_BU261 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N8,
      IB => rx_input_fifo_fifo_N3957,
      SEL => rx_input_fifo_fifo_N3960,
      O => rx_input_fifo_fifo_N9_CYMUXG
    );
  rx_input_fifo_fifo_BU262 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N3957,
      I1 => rx_input_fifo_fifo_N3960,
      O => rx_input_fifo_fifo_N3938
    );
  rx_input_fifo_fifo_N9_CYINIT_19 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3952,
      O => rx_input_fifo_fifo_N9_CYINIT
    );
  rx_input_fifo_fifo_N2434_LOGIC_ONE_20 : X_ONE
    port map (
      O => rx_input_fifo_fifo_N2434_LOGIC_ONE
    );
  rx_input_fifo_fifo_N2434_LOGIC_ZERO_21 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N2434_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU404 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2434_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2434_LOGIC_ONE,
      SEL => rx_input_fifo_fifo_N4900,
      O => rx_input_fifo_fifo_N4910
    );
  rx_input_fifo_fifo_BU403 : X_LUT4
    generic map(
      INIT => X"99C3"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2426,
      ADR1 => rx_input_fifo_fifo_N2486,
      ADR2 => rx_input_fifo_fifo_N2436,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N4900
    );
  rx_input_fifo_fifo_BU406 : X_LUT4
    generic map(
      INIT => X"99C3"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2425,
      ADR1 => rx_input_fifo_fifo_N2485,
      ADR2 => rx_input_fifo_fifo_N2435,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N4899
    );
  rx_input_fifo_fifo_N2434_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2434_CYMUXG,
      O => rx_input_fifo_fifo_N4909
    );
  rx_input_fifo_fifo_BU407 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2434_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N4910,
      SEL => rx_input_fifo_fifo_N4899,
      O => rx_input_fifo_fifo_N2434_CYMUXG
    );
  rx_input_fifo_fifo_N2443_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2443_FFY_RST
    );
  rx_input_fifo_fifo_BU466 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2404,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2443_FFY_RST,
      O => rx_input_fifo_fifo_N2444
    );
  rx_input_fifo_fifo_BU587 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2474,
      IB => rx_input_fifo_fifo_N6339_CYINIT,
      SEL => rx_input_fifo_fifo_N6332,
      O => rx_input_fifo_fifo_N6335
    );
  rx_input_fifo_fifo_BU586 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2474,
      ADR1 => rx_input_fifo_fifo_N2454,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N6332
    );
  rx_input_fifo_fifo_BU589 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2473,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N2453,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N6336
    );
  rx_input_fifo_fifo_N6339_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N6339_CYMUXG,
      O => rx_input_fifo_fifo_N6339
    );
  rx_input_fifo_fifo_BU590 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2473,
      IB => rx_input_fifo_fifo_N6335,
      SEL => rx_input_fifo_fifo_N6336,
      O => rx_input_fifo_fifo_N6339_CYMUXG
    );
  rx_input_fifo_fifo_N6339_CYINIT_22 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N6331,
      O => rx_input_fifo_fifo_N6339_CYINIT
    );
  rx_input_fifo_fifo_BU478 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2398,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2438_FFX_RST,
      O => rx_input_fifo_fifo_N2438
    );
  rx_input_fifo_fifo_N2438_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2438_FFX_RST
    );
  rx_input_fifo_fifo_BU528 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2442,
      ADR1 => rx_input_fifo_fifo_N5330,
      ADR2 => rx_input_fifo_fifo_N2443,
      ADR3 => rx_input_fifo_fifo_N2441,
      O => rx_input_fifo_fifo_N5344
    );
  rx_input_fifo_fifo_BU540 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N5329,
      ADR2 => rx_input_fifo_fifo_N5330,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N5343
    );
  rx_input_fifo_fifo_BU307 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N10,
      ADR1 => rx_input_fifo_fifo_N11,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4370
    );
  rx_input_fifo_fifo_BU314 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N10,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N9,
      O => rx_input_fifo_fifo_N4410
    );
  rx_input_fifo_fifo_N11_LOGIC_ZERO_23 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N11_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU243 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N11,
      IB => rx_input_fifo_fifo_N11_CYINIT,
      SEL => rx_input_fifo_fifo_N3945,
      O => rx_input_fifo_fifo_N3947
    );
  rx_input_fifo_fifo_BU244 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N11_CYINIT,
      I1 => rx_input_fifo_fifo_N3945,
      O => rx_input_fifo_fifo_N3935
    );
  rx_input_fifo_fifo_BU242 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N11,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3945
    );
  rx_input_fifo_fifo_BU248 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N10,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3950
    );
  rx_input_fifo_fifo_N11_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N11_CYMUXG,
      O => rx_input_fifo_fifo_N3952
    );
  rx_input_fifo_fifo_BU249 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N10,
      IB => rx_input_fifo_fifo_N3947,
      SEL => rx_input_fifo_fifo_N3950,
      O => rx_input_fifo_fifo_N11_CYMUXG
    );
  rx_input_fifo_fifo_BU250 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N3947,
      I1 => rx_input_fifo_fifo_N3950,
      O => rx_input_fifo_fifo_N3936
    );
  rx_input_fifo_fifo_N11_CYINIT_24 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N11_LOGIC_ZERO,
      O => rx_input_fifo_fifo_N11_CYINIT
    );
  rx_input_fifo_fifo_BU397 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_ince,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N2436_GROM
    );
  rx_input_fifo_fifo_N2436_YUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2436_GROM,
      O => rx_input_fifo_fifo_N4912
    );
  rx_input_fifo_fifo_N2475_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2475_FFY_SET
    );
  rx_input_fifo_fifo_BU440 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N11,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2475_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2476
    );
  rx_input_fifo_fifo_N6331_LOGIC_ONE_25 : X_ONE
    port map (
      O => rx_input_fifo_fifo_N6331_LOGIC_ONE
    );
  rx_input_fifo_fifo_BU581 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2476,
      IB => rx_input_fifo_fifo_N6331_LOGIC_ONE,
      SEL => rx_input_fifo_fifo_N6324,
      O => rx_input_fifo_fifo_N6327
    );
  rx_input_fifo_fifo_BU580 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2476,
      ADR1 => rx_input_fifo_fifo_N2456,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N6324
    );
  rx_input_fifo_fifo_BU583 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2475,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N2455,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N6328
    );
  rx_input_fifo_fifo_N6331_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N6331_CYMUXG,
      O => rx_input_fifo_fifo_N6331
    );
  rx_input_fifo_fifo_BU584 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2475,
      IB => rx_input_fifo_fifo_N6327,
      SEL => rx_input_fifo_fifo_N6328,
      O => rx_input_fifo_fifo_N6331_CYMUXG
    );
  rx_input_fifo_fifo_BU546 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N5330,
      ADR1 => rx_input_fifo_fifo_N2445,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N5329,
      O => rx_input_fifo_fifo_N5342
    );
  rx_input_fifo_fifo_BU552 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2445,
      ADR1 => rx_input_fifo_fifo_N2446,
      ADR2 => rx_input_fifo_fifo_N5330,
      ADR3 => rx_input_fifo_fifo_N5329,
      O => rx_input_fifo_fifo_N5341
    );
  rx_input_fifo_fifo_BU458 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2467_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2467
    );
  rx_input_fifo_fifo_N2467_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2467_FFX_SET
    );
  rx_input_fifo_fifo_BU28 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_empty,
      ADR3 => rx_input_fifo_rd_en,
      O => rx_input_fifo_fifo_N2362_FROM
    );
  rx_input_fifo_fifo_BU34 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_empty,
      ADR3 => rx_input_fifo_rd_en,
      O => rx_input_fifo_fifo_N2362_GROM
    );
  rx_input_fifo_fifo_N2362_XUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2362_FROM,
      O => rx_input_fifo_fifo_N2362
    );
  rx_input_fifo_fifo_N2362_YUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2362_GROM,
      O => rx_input_fifo_fifo_N22
    );
  rx_input_fifo_fifo_BU572 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N5349,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2447_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2448
    );
  rx_input_fifo_fifo_N2447_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2447_FFY_SET
    );
  rx_input_fifo_fifo_BU41 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_empty,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_rd_en,
      O => rx_input_fifo_fifo_N2724
    );
  rx_input_fifo_fifo_BU219 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_empty_CYINIT,
      I1 => rx_input_fifo_fifo_empty_FROM,
      O => rx_input_fifo_fifo_N3647
    );
  rx_input_fifo_fifo_empty_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_empty_FROM
    );
  rx_input_fifo_fifo_empty_CYINIT_26 : X_BUF
    port map (
      I => rx_input_fifo_fifo_BU216_O,
      O => rx_input_fifo_fifo_empty_CYINIT
    );
  mac_control_lmacaddr_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_27_FFY_RST
    );
  mac_control_lmacaddr_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_27_FFY_RST,
      O => mac_control_lmacaddr(26)
    );
  mac_control_lmacaddr_37_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_37_FFY_RST
    );
  mac_control_lmacaddr_36 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_37_FFY_RST,
      O => mac_control_lmacaddr(36)
    );
  mac_control_lmacaddr_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_45_FFY_RST
    );
  mac_control_lmacaddr_44 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_45_FFY_RST,
      O => mac_control_lmacaddr(44)
    );
  mac_control_lmacaddr_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_29_FFY_RST
    );
  mac_control_lmacaddr_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_29_FFY_RST,
      O => mac_control_lmacaddr(28)
    );
  mac_control_lmacaddr_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_39_FFY_RST
    );
  mac_control_lmacaddr_38 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_39_FFY_RST,
      O => mac_control_lmacaddr(38)
    );
  mac_control_lmacaddr_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_47_FFY_RST
    );
  mac_control_lmacaddr_46 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_47_FFY_RST,
      O => mac_control_lmacaddr(46)
    );
  rxbp_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_11_FFY_RST
    );
  rx_input_memio_BPOUT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_10_59,
      CE => rxbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_11_FFY_RST,
      O => rxbp(10)
    );
  rxbp_11_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxbp_11_CEMUXNOT
    );
  rxbp_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_13_FFY_RST
    );
  rx_input_memio_BPOUT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_12_57,
      CE => rxbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_13_FFY_RST,
      O => rxbp(12)
    );
  rxbp_13_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxbp_13_CEMUXNOT
    );
  rxbp_15_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxbp_15_CEMUXNOT
    );
  rx_output_fifo_BU144 : X_LUT4
    generic map(
      INIT => X"EEEE"
    )
    port map (
      ADR0 => rx_output_fifo_empty,
      ADR1 => rx_output_denll,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N2579_FROM
    );
  rx_output_fifo_BU22 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_denll,
      ADR2 => rx_output_fifo_empty,
      ADR3 => VCC,
      O => rx_output_fifo_N2579_GROM
    );
  rx_output_fifo_N2579_XUSED : X_BUF
    port map (
      I => rx_output_fifo_N2579_FROM,
      O => rx_output_fifo_N2579
    );
  rx_output_fifo_N2579_YUSED : X_BUF
    port map (
      I => rx_output_fifo_N2579_GROM,
      O => rx_output_fifo_N18
    );
  rx_output_fifo_BU29 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_denll,
      ADR2 => rx_output_fifo_empty,
      ADR3 => VCC,
      O => rx_output_fifo_N1835
    );
  rx_output_fifo_BU16 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_denll,
      ADR2 => rx_output_fifo_empty,
      ADR3 => VCC,
      O => rx_output_invalid_GROM
    );
  rx_output_invalid_YUSED : X_BUF
    port map (
      I => rx_output_invalid_GROM,
      O => rx_output_fifo_N1515
    );
  q2_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_1_FFY_RST
    );
  memcontroller_Q2_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(0),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_1_FFY_RST,
      O => q2(0)
    );
  mac_control_Ker52136_2_27 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => mac_control_bitcnt_104,
      ADR1 => mac_control_bitcnt_106,
      ADR2 => VCC,
      ADR3 => mac_control_bitcnt_105,
      O => mac_control_Ker52136_2_GROM
    );
  mac_control_Ker52136_2_YUSED : X_BUF
    port map (
      I => mac_control_Ker52136_2_GROM,
      O => mac_control_Ker52136_2
    );
  q3_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_1_FFY_RST
    );
  memcontroller_Q3_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(0),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_1_FFY_RST,
      O => q3(0)
    );
  q2_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_7_FFY_RST
    );
  memcontroller_Q2_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(6),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_7_FFY_RST,
      O => q2(6)
    );
  q3_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_3_FFY_RST
    );
  memcontroller_Q3_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(2),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_3_FFY_RST,
      O => q3(2)
    );
  q2_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_9_FFY_RST
    );
  memcontroller_Q2_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(8),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_9_FFY_RST,
      O => q2(8)
    );
  q3_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_5_FFY_RST
    );
  memcontroller_Q3_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(4),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_5_FFY_RST,
      O => q3(4)
    );
  rxfbbp_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_11_FFY_RST
    );
  rx_output_FBBP_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(10),
      CE => rxfbbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_11_FFY_RST,
      O => rxfbbp(10)
    );
  rxfbbp_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_11_CEMUXNOT
    );
  q3_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_7_FFY_RST
    );
  memcontroller_Q3_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(6),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_7_FFY_RST,
      O => q3(6)
    );
  rxfbbp_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_13_FFY_RST
    );
  rx_output_FBBP_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(12),
      CE => rxfbbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_13_FFY_RST,
      O => rxfbbp(12)
    );
  rxfbbp_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_13_CEMUXNOT
    );
  q3_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_9_FFY_RST
    );
  memcontroller_Q3_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(8),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_9_FFY_RST,
      O => q3(8)
    );
  rxfbbp_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_15_FFY_RST
    );
  rx_output_FBBP_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(14),
      CE => rxfbbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_15_FFY_RST,
      O => rxfbbp(14)
    );
  rxfbbp_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_15_CEMUXNOT
    );
  rxfifowerrsr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfifowerrsr_FFY_RST
    );
  slowclock_RXFIFOWERRSR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_rxfifowerrl,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfifowerrsr_FFY_RST,
      O => rxfifowerrsr
    );
  tx_output_bpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_11_FFY_RST
    );
  tx_output_bpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(10),
      CE => tx_output_bpl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_11_FFY_RST,
      O => tx_output_bpl(10)
    );
  tx_output_bpl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bpl_11_CEMUXNOT
    );
  tx_output_bpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_13_FFY_RST
    );
  tx_output_bpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(12),
      CE => tx_output_bpl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_13_FFY_RST,
      O => tx_output_bpl(12)
    );
  tx_output_bpl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bpl_13_CEMUXNOT
    );
  tx_output_bpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_15_FFY_RST
    );
  tx_output_bpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(14),
      CE => tx_output_bpl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_15_FFY_RST,
      O => tx_output_bpl(14)
    );
  tx_output_bpl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bpl_15_CEMUXNOT
    );
  rx_input_fifo_fifo_BU282 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3941,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N5_FFX_RST,
      O => rx_input_fifo_fifo_N5
    );
  rx_input_fifo_fifo_N5_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N5_FFX_RST
    );
  tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2_28 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => tx_output_data(5),
      ADR1 => VCC,
      ADR2 => tx_output_crcl(26),
      ADR3 => tx_output_crcl(28),
      O => tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2_FROM
    );
  tx_output_crc_loigc_Mxor_CO_25_Xo_1_1_2_29 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => tx_output_data(5),
      ADR1 => VCC,
      ADR2 => tx_output_crcl(17),
      ADR3 => tx_output_crcl(26),
      O => tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2_GROM
    );
  tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2_FROM,
      O => tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2
    );
  tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2_GROM,
      O => tx_output_crc_loigc_Mxor_CO_25_Xo_1_1_2
    );
  tx_output_outsell_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outsell_2_FFY_RST
    );
  tx_output_outsell_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_outsel_3_Q,
      CE => tx_output_outsell_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outsell_2_FFY_RST,
      O => tx_output_outsell(3)
    );
  tx_output_cs_Out1132 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_cs_FFd11,
      ADR1 => tx_output_cs_FFd14,
      ADR2 => tx_output_cs_FFd10,
      ADR3 => tx_output_cs_FFd13,
      O => tx_output_outsell_2_FROM
    );
  tx_output_cs_Out1160 : X_LUT4
    generic map(
      INIT => X"0040"
    )
    port map (
      ADR0 => tx_output_cs_Out1160_2,
      ADR1 => tx_output_CHOICE1634,
      ADR2 => tx_output_CHOICE1641,
      ADR3 => tx_output_cs_Out1160_SW0_1,
      O => tx_output_outsel_3_Q
    );
  tx_output_outsell_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_outsell_2_CEMUXNOT
    );
  tx_output_outsell_2_XUSED : X_BUF
    port map (
      I => tx_output_outsell_2_FROM,
      O => tx_output_CHOICE1634
    );
  rx_input_fifo_fifo_BU390 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2399,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2420_FFY_RST,
      O => rx_input_fifo_fifo_N2419
    );
  rx_input_fifo_fifo_N2420_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2420_FFY_RST
    );
  slowclock_txfifowerrl_LOGIC_ZERO_30 : X_ZERO
    port map (
      O => slowclock_txfifowerrl_LOGIC_ZERO
    );
  slowclock_txfifowerrl_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => slowclock_txfifowerrl_GROM
    );
  rx_input_memio_fifofulll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_fifofulll_FFY_RST
    );
  rx_input_memio_fifofulll_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfifofull,
      CE => rx_input_memio_fifofulll_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_fifofulll_FFY_RST,
      O => rx_input_memio_fifofulll
    );
  rx_input_memio_fifofulll_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_fifofulll_CEMUXNOT
    );
  rx_input_memio_endbyte_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_endbyte_1_FFY_RST
    );
  rx_input_memio_endbyte_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_endbyte_1_FFY_RST,
      O => rx_input_memio_endbyte(0)
    );
  rx_input_memio_endbyte_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_endbyte_2_FFY_RST
    );
  rx_input_memio_endbyte_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_endbyte_2_FFY_RST,
      O => rx_input_memio_endbyte(2)
    );
  rx_output_nfl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_nfl_FFY_RST
    );
  rx_output_nfl_32 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_nf,
      CE => rx_output_nfl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_nfl_FFY_RST,
      O => rx_output_nfl
    );
  rx_output_nfl_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_nfl_CEMUXNOT
    );
  mac_control_addr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_1_FFY_RST
    );
  mac_control_addr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_Mshreg_sinlll_102,
      CE => mac_control_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_addr_1_FFY_RST,
      O => mac_control_addr(0)
    );
  mac_control_addr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_3_FFY_RST
    );
  mac_control_addr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(1),
      CE => mac_control_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_addr_3_FFY_RST,
      O => mac_control_addr(2)
    );
  mac_control_addr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_5_FFY_RST
    );
  mac_control_addr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(3),
      CE => mac_control_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_addr_5_FFY_RST,
      O => mac_control_addr(4)
    );
  mac_control_addr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_7_FFY_RST
    );
  mac_control_addr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(5),
      CE => mac_control_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_addr_7_FFY_RST,
      O => mac_control_addr(6)
    );
  rx_input_fifo_fifo_BU420 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2420,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2431_FFY_RST,
      O => rx_input_fifo_fifo_N2430
    );
  rx_input_fifo_fifo_N2431_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2431_FFY_RST
    );
  tx_input_Ker3448049 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_input_CNT(11),
      ADR1 => tx_input_CNT(10),
      ADR2 => tx_input_CNT(9),
      ADR3 => tx_input_CNT(8),
      O => tx_input_CHOICE1710_FROM
    );
  tx_input_Ker34480111 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => tx_input_CNT(11),
      ADR1 => tx_input_CNT(8),
      ADR2 => tx_input_CNT(10),
      ADR3 => tx_input_CNT(9),
      O => tx_input_CHOICE1710_GROM
    );
  tx_input_CHOICE1710_XUSED : X_BUF
    port map (
      I => tx_input_CHOICE1710_FROM,
      O => tx_input_CHOICE1710
    );
  tx_input_CHOICE1710_YUSED : X_BUF
    port map (
      I => tx_input_CHOICE1710_GROM,
      O => tx_input_CHOICE1729
    );
  tx_input_Ker3448062 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_input_CNT(12),
      ADR1 => tx_input_CNT(13),
      ADR2 => tx_input_CNT(14),
      ADR3 => tx_input_CNT(15),
      O => tx_input_CHOICE1717_FROM
    );
  tx_input_Ker34480116 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => tx_input_CNT(12),
      ADR1 => tx_input_CNT(13),
      ADR2 => tx_input_CNT(15),
      ADR3 => tx_input_CNT(14),
      O => tx_input_CHOICE1717_GROM
    );
  tx_input_CHOICE1717_XUSED : X_BUF
    port map (
      I => tx_input_CHOICE1717_FROM,
      O => tx_input_CHOICE1717
    );
  tx_input_CHOICE1717_YUSED : X_BUF
    port map (
      I => tx_input_CHOICE1717_GROM,
      O => tx_input_CHOICE1732
    );
  tx_input_Ker34480137 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_input_N81681,
      ADR3 => tx_input_Ker34480137_2,
      O => tx_input_cs_FFd10_FROM
    );
  tx_input_cs_FFd10_In_33 : X_LUT4
    generic map(
      INIT => X"FAFE"
    )
    port map (
      ADR0 => tx_input_cs_FFd11,
      ADR1 => tx_input_cs_FFd6,
      ADR2 => tx_input_N69350,
      ADR3 => tx_input_N73800,
      O => tx_input_cs_FFd10_In
    );
  tx_input_cs_FFd10_XUSED : X_BUF
    port map (
      I => tx_input_cs_FFd10_FROM,
      O => tx_input_N73800
    );
  mac_control_din_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_11_FFY_RST
    );
  mac_control_din_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_11_FFY_RST,
      O => mac_control_din(10)
    );
  rx_input_fifo_fifo_N2497_LOGIC_ZERO_34 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N2497_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU213 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2497_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2497_CYINIT,
      SEL => rx_input_fifo_fifo_N3626,
      O => rx_input_fifo_fifo_N3636
    );
  rx_input_fifo_fifo_BU212 : X_LUT4
    generic map(
      INIT => X"A599"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2398,
      ADR1 => rx_input_fifo_fifo_N2498,
      ADR2 => rx_input_fifo_fifo_N2478,
      ADR3 => rx_input_fifo_fifo_empty,
      O => rx_input_fifo_fifo_N3626
    );
  rx_input_fifo_fifo_BU215 : X_LUT4
    generic map(
      INIT => X"9C93"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2477,
      ADR1 => rx_input_fifo_fifo_N2397,
      ADR2 => rx_input_fifo_fifo_empty,
      ADR3 => rx_input_fifo_fifo_N2497,
      O => rx_input_fifo_fifo_N3625
    );
  rx_input_fifo_fifo_N2497_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2497_CYMUXG,
      O => rx_input_fifo_fifo_BU216_O
    );
  rx_input_fifo_fifo_BU216 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2497_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N3636,
      SEL => rx_input_fifo_fifo_N3625,
      O => rx_input_fifo_fifo_N2497_CYMUXG
    );
  rx_input_fifo_fifo_N2497_CYINIT_35 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3637,
      O => rx_input_fifo_fifo_N2497_CYINIT
    );
  rx_input_fifo_fifo_BU177 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N12,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3600
    );
  rx_input_fifo_fifo_BU170 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N13,
      ADR2 => rx_input_fifo_fifo_N12,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3560
    );
  rx_input_fifo_fifo_BU98 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N13,
      IB => rx_input_fifo_fifo_N13_CYINIT,
      SEL => rx_input_fifo_fifo_N2855,
      O => rx_input_fifo_fifo_N2857
    );
  rx_input_fifo_fifo_BU99 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N13_CYINIT,
      I1 => rx_input_fifo_fifo_N2855,
      O => rx_input_fifo_fifo_N2813
    );
  rx_input_fifo_fifo_BU97 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N13,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2855
    );
  rx_input_fifo_fifo_BU103 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N12,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2860
    );
  rx_input_fifo_fifo_BU104 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N2857,
      I1 => rx_input_fifo_fifo_N2860,
      O => rx_input_fifo_fifo_N2814
    );
  rx_input_fifo_fifo_N13_CYINIT_36 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2852,
      O => rx_input_fifo_fifo_N13_CYINIT
    );
  rx_input_fifo_fifo_N2499_LOGIC_ZERO_37 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N2499_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU207 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2499_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2499_CYINIT,
      SEL => rx_input_fifo_fifo_N3628,
      O => rx_input_fifo_fifo_N3638
    );
  rx_input_fifo_fifo_BU206 : X_LUT4
    generic map(
      INIT => X"CA35"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2500,
      ADR1 => rx_input_fifo_fifo_N2480,
      ADR2 => rx_input_fifo_fifo_empty,
      ADR3 => rx_input_fifo_fifo_N2400,
      O => rx_input_fifo_fifo_N3628
    );
  rx_input_fifo_fifo_BU209 : X_LUT4
    generic map(
      INIT => X"A5C3"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2479,
      ADR1 => rx_input_fifo_fifo_N2499,
      ADR2 => rx_input_fifo_fifo_N2399,
      ADR3 => rx_input_fifo_fifo_empty,
      O => rx_input_fifo_fifo_N3627
    );
  rx_input_fifo_fifo_N2499_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2499_CYMUXG,
      O => rx_input_fifo_fifo_N3637
    );
  rx_input_fifo_fifo_BU210 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2499_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N3638,
      SEL => rx_input_fifo_fifo_N3627,
      O => rx_input_fifo_fifo_N2499_CYMUXG
    );
  rx_input_fifo_fifo_N2499_CYINIT_38 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3639,
      O => rx_input_fifo_fifo_N2499_CYINIT
    );
  rx_input_fifo_fifo_BU156 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N14,
      ADR1 => rx_input_fifo_fifo_N15,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3480
    );
  rx_input_fifo_fifo_BU163 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N14,
      ADR1 => rx_input_fifo_fifo_N13,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3520
    );
  rx_input_fifo_fifo_BU86 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N15,
      IB => rx_input_fifo_fifo_N15_CYINIT,
      SEL => rx_input_fifo_fifo_N2845,
      O => rx_input_fifo_fifo_N2847
    );
  rx_input_fifo_fifo_BU87 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N15_CYINIT,
      I1 => rx_input_fifo_fifo_N2845,
      O => rx_input_fifo_fifo_N2811
    );
  rx_input_fifo_fifo_BU85 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N15,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2845
    );
  rx_input_fifo_fifo_BU91 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N14,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2850
    );
  rx_input_fifo_fifo_N15_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N15_CYMUXG,
      O => rx_input_fifo_fifo_N2852
    );
  rx_input_fifo_fifo_BU92 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N14,
      IB => rx_input_fifo_fifo_N2847,
      SEL => rx_input_fifo_fifo_N2850,
      O => rx_input_fifo_fifo_N15_CYMUXG
    );
  rx_input_fifo_fifo_BU93 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N2847,
      I1 => rx_input_fifo_fifo_N2850,
      O => rx_input_fifo_fifo_N2812
    );
  rx_input_fifo_fifo_N15_CYINIT_39 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2842,
      O => rx_input_fifo_fifo_N15_CYINIT
    );
  rx_input_fifo_fifo_N2500_LOGIC_ZERO_40 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N2500_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU201 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2500_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2500_CYINIT,
      SEL => rx_input_fifo_fifo_N3630,
      O => rx_input_fifo_fifo_N3640
    );
  rx_input_fifo_fifo_BU200 : X_LUT4
    generic map(
      INIT => X"D287"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_empty,
      ADR1 => rx_input_fifo_fifo_N2482,
      ADR2 => rx_input_fifo_fifo_N2402,
      ADR3 => rx_input_fifo_fifo_N2502,
      O => rx_input_fifo_fifo_N3630
    );
  rx_input_fifo_fifo_BU203 : X_LUT4
    generic map(
      INIT => X"AC53"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2481,
      ADR1 => rx_input_fifo_fifo_N2501,
      ADR2 => rx_input_fifo_fifo_empty,
      ADR3 => rx_input_fifo_fifo_N2401,
      O => rx_input_fifo_fifo_N3629
    );
  rx_input_fifo_fifo_N2500_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2500_CYMUXG,
      O => rx_input_fifo_fifo_N3639
    );
  rx_input_fifo_fifo_BU204 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2500_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N3640,
      SEL => rx_input_fifo_fifo_N3629,
      O => rx_input_fifo_fifo_N2500_CYMUXG
    );
  rx_input_fifo_fifo_N2500_CYINIT_41 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3641,
      O => rx_input_fifo_fifo_N2500_CYINIT
    );
  rx_input_fifo_fifo_BU149 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N15,
      ADR1 => rx_input_fifo_fifo_N16,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3440
    );
  rx_input_fifo_fifo_BU142 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N16,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N17,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3400
    );
  rx_input_fifo_fifo_BU74 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N17,
      IB => rx_input_fifo_fifo_N17_CYINIT,
      SEL => rx_input_fifo_fifo_N2835,
      O => rx_input_fifo_fifo_N2837
    );
  rx_input_fifo_fifo_BU75 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N17_CYINIT,
      I1 => rx_input_fifo_fifo_N2835,
      O => rx_input_fifo_fifo_N2809
    );
  rx_input_fifo_fifo_BU73 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N17,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2835
    );
  rx_input_fifo_fifo_BU79 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N16,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2840
    );
  rx_input_fifo_fifo_N17_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N17_CYMUXG,
      O => rx_input_fifo_fifo_N2842
    );
  rx_input_fifo_fifo_BU80 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N16,
      IB => rx_input_fifo_fifo_N2837,
      SEL => rx_input_fifo_fifo_N2840,
      O => rx_input_fifo_fifo_N17_CYMUXG
    );
  rx_input_fifo_fifo_BU81 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N2837,
      I1 => rx_input_fifo_fifo_N2840,
      O => rx_input_fifo_fifo_N2810
    );
  rx_input_fifo_fifo_N17_CYINIT_42 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2832,
      O => rx_input_fifo_fifo_N17_CYINIT
    );
  rx_input_fifo_fifo_N2502_LOGIC_ZERO_43 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N2502_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU195 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2502_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2502_CYINIT,
      SEL => rx_input_fifo_fifo_N3632,
      O => rx_input_fifo_fifo_N3642
    );
  rx_input_fifo_fifo_BU194 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2504,
      ADR1 => rx_input_fifo_fifo_N2404,
      ADR2 => rx_input_fifo_fifo_N2484,
      ADR3 => rx_input_fifo_fifo_empty,
      O => rx_input_fifo_fifo_N3632
    );
  rx_input_fifo_fifo_BU197 : X_LUT4
    generic map(
      INIT => X"9C93"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2483,
      ADR1 => rx_input_fifo_fifo_N2403,
      ADR2 => rx_input_fifo_fifo_empty,
      ADR3 => rx_input_fifo_fifo_N2503,
      O => rx_input_fifo_fifo_N3631
    );
  rx_input_fifo_fifo_N2502_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2502_CYMUXG,
      O => rx_input_fifo_fifo_N3641
    );
  rx_input_fifo_fifo_BU198 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2502_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N3642,
      SEL => rx_input_fifo_fifo_N3631,
      O => rx_input_fifo_fifo_N2502_CYMUXG
    );
  rx_input_fifo_fifo_N2502_CYINIT_44 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3643,
      O => rx_input_fifo_fifo_N2502_CYINIT
    );
  rx_input_fifo_fifo_BU128 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N18,
      ADR1 => rx_input_fifo_fifo_N19,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3320
    );
  rx_input_fifo_fifo_BU135 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N17,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N18,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3360
    );
  rx_input_fifo_fifo_BU62 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N19,
      IB => rx_input_fifo_fifo_N19_CYINIT,
      SEL => rx_input_fifo_fifo_N2825,
      O => rx_input_fifo_fifo_N2827
    );
  rx_input_fifo_fifo_BU63 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N19_CYINIT,
      I1 => rx_input_fifo_fifo_N2825,
      O => rx_input_fifo_fifo_N2807
    );
  rx_input_fifo_fifo_BU61 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N19,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2825
    );
  rx_input_fifo_fifo_BU67 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N18,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2830
    );
  rx_input_fifo_fifo_N19_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N19_CYMUXG,
      O => rx_input_fifo_fifo_N2832
    );
  rx_input_fifo_fifo_BU68 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N18,
      IB => rx_input_fifo_fifo_N2827,
      SEL => rx_input_fifo_fifo_N2830,
      O => rx_input_fifo_fifo_N19_CYMUXG
    );
  rx_input_fifo_fifo_BU69 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N2827,
      I1 => rx_input_fifo_fifo_N2830,
      O => rx_input_fifo_fifo_N2808
    );
  rx_input_fifo_fifo_N19_CYINIT_45 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2822,
      O => rx_input_fifo_fifo_N19_CYINIT
    );
  rx_input_fifo_fifo_N2504_LOGIC_ONE_46 : X_ONE
    port map (
      O => rx_input_fifo_fifo_N2504_LOGIC_ONE
    );
  rx_input_fifo_fifo_N2504_LOGIC_ZERO_47 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N2504_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU189 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2504_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2504_LOGIC_ONE,
      SEL => rx_input_fifo_fifo_N3634,
      O => rx_input_fifo_fifo_N3644
    );
  rx_input_fifo_fifo_BU188 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2506,
      ADR1 => rx_input_fifo_fifo_N2406,
      ADR2 => rx_input_fifo_fifo_N2486,
      ADR3 => rx_input_fifo_fifo_empty,
      O => rx_input_fifo_fifo_N3634
    );
  rx_input_fifo_fifo_BU191 : X_LUT4
    generic map(
      INIT => X"E41B"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_empty,
      ADR1 => rx_input_fifo_fifo_N2505,
      ADR2 => rx_input_fifo_fifo_N2485,
      ADR3 => rx_input_fifo_fifo_N2405,
      O => rx_input_fifo_fifo_N3633
    );
  rx_input_fifo_fifo_N2504_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2504_CYMUXG,
      O => rx_input_fifo_fifo_N3643
    );
  rx_input_fifo_fifo_BU192 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N2504_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N3644,
      SEL => rx_input_fifo_fifo_N3633,
      O => rx_input_fifo_fifo_N2504_CYMUXG
    );
  rx_input_fifo_fifo_BU114 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N21,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N20,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3240
    );
  rx_input_fifo_fifo_BU121 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N20,
      ADR3 => rx_input_fifo_fifo_N19,
      O => rx_input_fifo_fifo_N3280
    );
  rx_input_fifo_fifo_N21_LOGIC_ZERO_48 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N21_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU50 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N21,
      IB => rx_input_fifo_fifo_N21_CYINIT,
      SEL => rx_input_fifo_fifo_N2815,
      O => rx_input_fifo_fifo_N2817
    );
  rx_input_fifo_fifo_BU51 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N21_CYINIT,
      I1 => rx_input_fifo_fifo_N2815,
      O => rx_input_fifo_fifo_N2805
    );
  rx_input_fifo_fifo_BU49 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N21,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2815
    );
  rx_input_fifo_fifo_BU55 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N20,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2820
    );
  rx_input_fifo_fifo_N21_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N21_CYMUXG,
      O => rx_input_fifo_fifo_N2822
    );
  rx_input_fifo_fifo_BU56 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N20,
      IB => rx_input_fifo_fifo_N2817,
      SEL => rx_input_fifo_fifo_N2820,
      O => rx_input_fifo_fifo_N21_CYMUXG
    );
  rx_input_fifo_fifo_BU57 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N2817,
      I1 => rx_input_fifo_fifo_N2820,
      O => rx_input_fifo_fifo_N2806
    );
  rx_input_fifo_fifo_N21_CYINIT_49 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N21_LOGIC_ZERO,
      O => rx_input_fifo_fifo_N21_CYINIT
    );
  rx_input_fifo_fifo_BU182 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_empty,
      ADR3 => rx_input_fifo_rd_en,
      O => rx_input_fifo_fifo_N2505_GROM
    );
  rx_input_fifo_fifo_N2505_YUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2505_GROM,
      O => rx_input_fifo_fifo_N3646
    );
  slowclock_n00021 : X_LUT4
    generic map(
      INIT => X"8080"
    )
    port map (
      ADR0 => slowclock_clkcnt(1),
      ADR1 => slowclock_clkcnt(0),
      ADR2 => slowclock_clkcnt(2),
      ADR3 => VCC,
      O => slowclock_n0002_FROM
    );
  slowclock_n00051 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => slowclock_clkcnt(1),
      ADR1 => slowclock_clkcnt(0),
      ADR2 => VCC,
      ADR3 => slowclock_clkcnt(2),
      O => slowclock_n0002_GROM
    );
  slowclock_n0002_XUSED : X_BUF
    port map (
      I => slowclock_n0002_FROM,
      O => slowclock_n0002
    );
  slowclock_n0002_YUSED : X_BUF
    port map (
      I => slowclock_n0002_GROM,
      O => slowclock_n0005
    );
  rx_input_fifo_control_dinl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_dinl_9_CEMUXNOT
    );
  tx_input_dh_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_13_FFY_RST
    );
  tx_input_dh_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(12),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_13_FFY_RST,
      O => tx_input_dh(12)
    );
  tx_input_dh_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_15_FFY_RST
    );
  tx_input_dh_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(14),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_15_FFY_RST,
      O => tx_input_dh(14)
    );
  mac_control_n007050_SW0 : X_LUT4
    generic map(
      INIT => X"F5FF"
    )
    port map (
      ADR0 => mac_control_CHOICE1616,
      ADR1 => VCC,
      ADR2 => mac_control_ledtx_cnt_153,
      ADR3 => mac_control_CHOICE1609,
      O => mac_control_N81797_FROM
    );
  mac_control_n00391 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_151,
      ADR1 => mac_control_ledtx_cnt_152,
      ADR2 => mac_control_ledtx_cnt_150,
      ADR3 => mac_control_N81797,
      O => mac_control_N81797_GROM
    );
  mac_control_N81797_XUSED : X_BUF
    port map (
      I => mac_control_N81797_FROM,
      O => mac_control_N81797
    );
  mac_control_N81797_YUSED : X_BUF
    port map (
      I => mac_control_N81797_GROM,
      O => mac_control_n0039
    );
  rx_input_GMII_lince1 : X_LUT4
    generic map(
      INIT => X"F3F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_GMII_rx_dvll,
      ADR2 => rx_input_GMII_ro,
      ADR3 => rx_input_GMII_rx_dvl,
      O => rx_input_GMII_lince
    );
  rx_input_GMII_dvdelta1 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_GMII_rx_dvll,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_GMII_rx_dvl,
      O => rx_input_ince_GROM
    );
  rx_input_ince_YUSED : X_BUF
    port map (
      I => rx_input_ince_GROM,
      O => rx_input_GMII_dvdelta
    );
  txbp_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_11_FFY_RST
    );
  tx_input_bp_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_26,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_11_FFY_RST,
      O => txbp(10)
    );
  tx_input_dl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_13_FFY_RST
    );
  tx_input_dl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(12),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_13_FFY_RST,
      O => tx_input_dl(12)
    );
  txbp_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_13_FFY_RST
    );
  tx_input_bp_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_28,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_13_FFY_RST,
      O => txbp(12)
    );
  rx_input_fifo_fifo_BU574 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2437,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2447_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2447
    );
  rx_input_fifo_fifo_N2447_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2447_FFX_SET
    );
  txbp_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_15_FFY_RST
    );
  tx_input_bp_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_30,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_15_FFY_RST,
      O => txbp(14)
    );
  mac_control_n007150_SW0 : X_LUT4
    generic map(
      INIT => X"DDFF"
    )
    port map (
      ADR0 => mac_control_CHOICE1593,
      ADR1 => mac_control_ledrx_cnt_165,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE1586,
      O => mac_control_N81777_FROM
    );
  mac_control_n00411 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_162,
      ADR1 => mac_control_ledrx_cnt_164,
      ADR2 => mac_control_ledrx_cnt_163,
      ADR3 => mac_control_N81777,
      O => mac_control_N81777_GROM
    );
  mac_control_N81777_XUSED : X_BUF
    port map (
      I => mac_control_N81777_FROM,
      O => mac_control_N81777
    );
  mac_control_N81777_YUSED : X_BUF
    port map (
      I => mac_control_N81777_GROM,
      O => mac_control_n0041
    );
  rx_input_memio_Ker411851 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => rx_input_endf,
      ADR1 => rx_input_invalid,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_cs_FFd1_FROM
    );
  rx_input_memio_addrchk_cs_FFd1_In1 : X_LUT4
    generic map(
      INIT => X"00B8"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd2,
      ADR1 => rx_input_memio_brdy,
      ADR2 => rx_input_memio_addrchk_cs_FFd1,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_addrchk_cs_FFd1_In
    );
  rx_input_memio_addrchk_cs_FFd1_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_cs_FFd1_FROM,
      O => rx_input_memio_brdy
    );
  rx_input_memio_addrchk_rxucastl_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_rxucastl_CEMUXNOT
    );
  rx_input_fifo_fifo_BU357 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N4650,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2480_FFY_RST,
      O => rx_input_fifo_fifo_N2479
    );
  rx_input_fifo_fifo_N2480_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2480_FFY_RST
    );
  mac_control_lmacaddr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_11_FFY_RST
    );
  mac_control_lmacaddr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_11_FFY_RST,
      O => mac_control_lmacaddr(10)
    );
  mac_control_lmacaddr_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_21_FFY_RST
    );
  mac_control_lmacaddr_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_21_FFY_RST,
      O => mac_control_lmacaddr(20)
    );
  mac_control_lmacaddr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_13_FFY_RST
    );
  mac_control_lmacaddr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_13_FFY_RST,
      O => mac_control_lmacaddr(12)
    );
  rx_input_fifo_fifo_BU288 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3942,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N5_FFY_RST,
      O => rx_input_fifo_fifo_N4
    );
  rx_input_fifo_fifo_N5_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N5_FFY_RST
    );
  mac_control_lmacaddr_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_23_FFY_RST
    );
  mac_control_lmacaddr_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_23_FFY_RST,
      O => mac_control_lmacaddr(22)
    );
  mac_control_lmacaddr_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_31_FFY_RST
    );
  mac_control_lmacaddr_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_31_FFY_RST,
      O => mac_control_lmacaddr(30)
    );
  mac_control_lmacaddr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_15_FFY_RST
    );
  mac_control_lmacaddr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_15_FFY_RST,
      O => mac_control_lmacaddr(14)
    );
  mac_control_lmacaddr_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_33_FFY_RST
    );
  mac_control_lmacaddr_32 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_33_FFY_RST,
      O => mac_control_lmacaddr(32)
    );
  mac_control_lmacaddr_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_41_FFY_RST
    );
  mac_control_lmacaddr_40 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_41_FFY_RST,
      O => mac_control_lmacaddr(40)
    );
  mac_control_lmacaddr_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_17_FFY_RST
    );
  mac_control_lmacaddr_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_17_FFY_RST,
      O => mac_control_lmacaddr(16)
    );
  mac_control_lmacaddr_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_25_FFY_RST
    );
  mac_control_lmacaddr_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_25_FFY_RST,
      O => mac_control_lmacaddr(24)
    );
  mac_control_lmacaddr_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_35_FFY_RST
    );
  mac_control_lmacaddr_34 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_35_FFY_RST,
      O => mac_control_lmacaddr(34)
    );
  rx_input_fifo_fifo_BU350 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N4610,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2480_FFX_RST,
      O => rx_input_fifo_fifo_N2480
    );
  rx_input_fifo_fifo_N2480_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2480_FFX_RST
    );
  mac_control_lmacaddr_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_43_FFY_RST
    );
  mac_control_lmacaddr_42 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_43_FFY_RST,
      O => mac_control_lmacaddr(42)
    );
  mac_control_lmacaddr_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_19_FFY_RST
    );
  mac_control_lmacaddr_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_19_FFY_RST,
      O => mac_control_lmacaddr(18)
    );
  rx_fifocheck_n000263 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_fifocheck_CHOICE1789,
      ADR2 => rx_fifocheck_CHOICE1796,
      ADR3 => VCC,
      O => rx_fifocheck_CHOICE1797_FROM
    );
  rx_fifocheck_n000292 : X_LUT4
    generic map(
      INIT => X"F8F0"
    )
    port map (
      ADR0 => rx_fifocheck_CHOICE1774,
      ADR1 => rx_fifocheck_CHOICE1781,
      ADR2 => rx_fifocheck_n0003,
      ADR3 => rx_fifocheck_CHOICE1797,
      O => rx_fifocheck_CHOICE1797_GROM
    );
  rx_fifocheck_CHOICE1797_XUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1797_FROM,
      O => rx_fifocheck_CHOICE1797
    );
  rx_fifocheck_CHOICE1797_YUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1797_GROM,
      O => rx_fifocheck_N74128
    );
  rx_fifocheck_n000249 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(11),
      ADR1 => rx_fifocheck_diff(9),
      ADR2 => rx_fifocheck_diff(10),
      ADR3 => rx_fifocheck_diff(8),
      O => rx_fifocheck_CHOICE1789_GROM
    );
  rx_fifocheck_CHOICE1789_YUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1789_GROM,
      O => rx_fifocheck_CHOICE1789
    );
  tx_output_cs_Out1160_SW0_1_50 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16,
      ADR2 => tx_output_cs_FFd8,
      ADR3 => VCC,
      O => tx_output_cs_Out1160_SW0_1_FROM
    );
  tx_output_n00251 : X_LUT4
    generic map(
      INIT => X"5550"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => tx_output_crcenl,
      ADR3 => tx_output_cs_FFd16,
      O => tx_output_cs_Out1160_SW0_1_GROM
    );
  tx_output_cs_Out1160_SW0_1_XUSED : X_BUF
    port map (
      I => tx_output_cs_Out1160_SW0_1_FROM,
      O => tx_output_cs_Out1160_SW0_1
    );
  tx_output_cs_Out1160_SW0_1_YUSED : X_BUF
    port map (
      I => tx_output_cs_Out1160_SW0_1_GROM,
      O => tx_output_n0025
    );
  tx_output_cs_Out149 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd6,
      ADR1 => tx_output_cs_FFd10,
      ADR2 => tx_output_cs_FFd9,
      ADR3 => tx_output_cs_FFd8,
      O => tx_output_CHOICE1679_FROM
    );
  tx_output_cs_Out1145 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_cs_FFd9,
      ADR1 => tx_output_cs_FFd17,
      ADR2 => tx_output_cs_FFd12,
      ADR3 => tx_output_cs_FFd15,
      O => tx_output_CHOICE1679_GROM
    );
  tx_output_CHOICE1679_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1679_FROM,
      O => tx_output_CHOICE1679
    );
  tx_output_CHOICE1679_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1679_GROM,
      O => tx_output_CHOICE1641
    );
  tx_output_ldata_3_18_SW0 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd4,
      ADR2 => VCC,
      ADR3 => tx_output_cs_FFd5,
      O => tx_output_N81625_FROM
    );
  tx_output_cs_Out1421 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd5,
      ADR1 => tx_output_cs_FFd7,
      ADR2 => tx_output_cs_FFd3,
      ADR3 => tx_output_cs_FFd4,
      O => tx_output_N81625_GROM
    );
  tx_output_N81625_XUSED : X_BUF
    port map (
      I => tx_output_N81625_FROM,
      O => tx_output_N81625
    );
  tx_output_N81625_YUSED : X_BUF
    port map (
      I => tx_output_N81625_GROM,
      O => tx_output_CHOICE1683
    );
  tx_output_n0034_5_1 : X_LUT4
    generic map(
      INIT => X"DDEE"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0056(2),
      ADR1 => tx_output_cs_FFd16,
      ADR2 => VCC,
      ADR3 => tx_output_crc_loigc_Mxor_CO_5_Xo_1_1_2,
      O => tx_output_n0034(5)
    );
  tx_output_cs_Out1426 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd1,
      ADR1 => tx_output_cs_FFd15,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_cs_FFd2,
      O => tx_output_crcl_5_GROM
    );
  tx_output_crcl_5_YUSED : X_BUF
    port map (
      I => tx_output_crcl_5_GROM,
      O => tx_output_CHOICE1686
    );
  tx_output_crc_loigc_Mxor_n0005_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(3),
      ADR1 => tx_output_crcl(28),
      ADR2 => tx_output_crc_loigc_n0104(0),
      ADR3 => tx_output_crc_loigc_n0122(1),
      O => tx_output_crcl_4_FROM
    );
  tx_output_n0034_4_1 : X_LUT4
    generic map(
      INIT => X"AFFA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => VCC,
      ADR2 => tx_output_crc_loigc_Mxor_CO_4_Xo_1_1_2,
      ADR3 => tx_output_crc_loigc_n0056(2),
      O => tx_output_n0034(4)
    );
  tx_output_crcl_4_XUSED : X_BUF
    port map (
      I => tx_output_crcl_4_FROM,
      O => tx_output_crc_loigc_n0056(2)
    );
  tx_output_crc_loigc_Mxor_n0007_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(6),
      ADR1 => tx_output_data(2),
      ADR2 => tx_output_crcl(29),
      ADR3 => tx_output_crcl(25),
      O => tx_output_crc_loigc_Mxor_n0007_Xo_0_FROM
    );
  tx_output_crc_loigc_Mxor_n0021_Result1 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => tx_output_crcl(29),
      ADR1 => tx_output_data(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_output_crc_loigc_Mxor_n0007_Xo_0_GROM
    );
  tx_output_crc_loigc_Mxor_n0007_Xo_0_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_n0007_Xo_0_FROM,
      O => tx_output_crc_loigc_Mxor_n0007_Xo(0)
    );
  tx_output_crc_loigc_Mxor_n0007_Xo_0_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_n0007_Xo_0_GROM,
      O => tx_output_crc_loigc_n0118(0)
    );
  tx_output_cs_Out13_2_51 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd8,
      ADR2 => tx_output_cs_FFd17,
      ADR3 => tx_output_cs_FFd4,
      O => tx_output_outsell_0_FROM
    );
  tx_output_cs_Out13 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => tx_output_cs_FFd5,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd6,
      ADR3 => tx_output_cs_Out13_2,
      O => tx_output_outsel_0_Q
    );
  tx_output_outsell_0_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_outsell_0_CEMUXNOT
    );
  tx_output_outsell_0_XUSED : X_BUF
    port map (
      I => tx_output_outsell_0_FROM,
      O => tx_output_cs_Out13_2
    );
  mac_control_n0035194_SW0 : X_LUT4
    generic map(
      INIT => X"8080"
    )
    port map (
      ADR0 => mac_control_CHOICE2770,
      ADR1 => mac_control_CHOICE2777,
      ADR2 => mac_control_n0035194_SW0_2,
      ADR3 => VCC,
      O => mac_control_N81689_FROM
    );
  mac_control_n0035194 : X_LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_141,
      ADR1 => mac_control_CHOICE2732,
      ADR2 => mac_control_CHOICE2739,
      ADR3 => mac_control_N81689,
      O => mac_control_N81689_GROM
    );
  mac_control_N81689_XUSED : X_BUF
    port map (
      I => mac_control_N81689_FROM,
      O => mac_control_N81689
    );
  mac_control_N81689_YUSED : X_BUF
    port map (
      I => mac_control_N81689_GROM,
      O => mac_control_N79380
    );
  rx_input_memio_n001610 : X_LUT4
    generic map(
      INIT => X"0400"
    )
    port map (
      ADR0 => rx_input_data(1),
      ADR1 => rx_input_data(0),
      ADR2 => rx_input_data(3),
      ADR3 => rx_input_data(2),
      O => rx_input_memio_CHOICE1447_GROM
    );
  rx_input_memio_CHOICE1447_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1447_GROM,
      O => rx_input_memio_CHOICE1447
    );
  rx_input_memio_n001618 : X_LUT4
    generic map(
      INIT => X"0080"
    )
    port map (
      ADR0 => rx_input_data(6),
      ADR1 => rx_input_data(7),
      ADR2 => rx_input_data(4),
      ADR3 => rx_input_data(5),
      O => rx_input_memio_CHOICE1451_GROM
    );
  rx_input_memio_CHOICE1451_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1451_GROM,
      O => rx_input_memio_CHOICE1451
    );
  rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2_52 : X_LUT4
    generic map(
      INIT => X"9696"
    )
    port map (
      ADR0 => rx_input_memio_crcl(31),
      ADR1 => rx_input_memio_datal(0),
      ADR2 => rx_input_memio_crcl(10),
      ADR3 => VCC,
      O => rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2_FROM
    );
  rx_input_memio_crccomb_Mxor_CO_30_Xo_1_1_2_53 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => rx_input_memio_crcl(31),
      ADR1 => rx_input_memio_datal(0),
      ADR2 => VCC,
      ADR3 => rx_input_memio_crcl(22),
      O => rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2
    );
  rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2_GROM,
      O => rx_input_memio_crccomb_Mxor_CO_30_Xo_1_1_2
    );
  rx_input_memio_n005915 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => rx_input_memio_crcll(4),
      ADR1 => rx_input_memio_crcll(7),
      ADR2 => rx_input_memio_crcll(6),
      ADR3 => rx_input_memio_crcll(5),
      O => rx_input_memio_CHOICE2917_FROM
    );
  rx_input_memio_n0059143_2_54 : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_CHOICE2922,
      ADR2 => rx_input_memio_CHOICE2913,
      ADR3 => rx_input_memio_CHOICE2917,
      O => rx_input_memio_CHOICE2917_GROM
    );
  rx_input_memio_CHOICE2917_XUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE2917_FROM,
      O => rx_input_memio_CHOICE2917
    );
  rx_input_memio_CHOICE2917_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE2917_GROM,
      O => rx_input_memio_n0059143_2
    );
  rx_input_memio_n005932 : X_LUT4
    generic map(
      INIT => X"0080"
    )
    port map (
      ADR0 => rx_input_memio_crcll(8),
      ADR1 => rx_input_memio_crcll(10),
      ADR2 => rx_input_memio_crcll(11),
      ADR3 => rx_input_memio_crcll(9),
      O => rx_input_memio_CHOICE2922_GROM
    );
  rx_input_memio_CHOICE2922_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE2922_GROM,
      O => rx_input_memio_CHOICE2922
    );
  rx_input_memio_n005940 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => rx_input_memio_crcll(13),
      ADR1 => rx_input_memio_crcll(14),
      ADR2 => rx_input_memio_crcll(12),
      ADR3 => rx_input_memio_crcll(15),
      O => rx_input_memio_CHOICE2926_GROM
    );
  rx_input_memio_CHOICE2926_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE2926_GROM,
      O => rx_input_memio_CHOICE2926
    );
  slowclock_lclken_LOGIC_ONE_55 : X_ONE
    port map (
      O => slowclock_lclken_LOGIC_ONE
    );
  rx_input_memio_n005975 : X_LUT4
    generic map(
      INIT => X"0100"
    )
    port map (
      ADR0 => rx_input_memio_crcll(19),
      ADR1 => rx_input_memio_crcll(17),
      ADR2 => rx_input_memio_crcll(16),
      ADR3 => rx_input_memio_crcll(18),
      O => rx_input_memio_CHOICE2934_FROM
    );
  rx_input_memio_n0059143_SW0_2_56 : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_CHOICE2926,
      ADR2 => rx_input_memio_CHOICE2941,
      ADR3 => rx_input_memio_CHOICE2934,
      O => rx_input_memio_CHOICE2934_GROM
    );
  rx_input_memio_CHOICE2934_XUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE2934_FROM,
      O => rx_input_memio_CHOICE2934
    );
  rx_input_memio_CHOICE2934_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE2934_GROM,
      O => rx_input_memio_n0059143_SW0_2
    );
  rx_input_fifo_fifo_BU258 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3937,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N9_FFX_RST,
      O => rx_input_fifo_fifo_N9
    );
  rx_input_fifo_fifo_N9_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N9_FFX_RST
    );
  rx_input_memio_n005988 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_input_memio_crcll(22),
      ADR1 => rx_input_memio_crcll(20),
      ADR2 => rx_input_memio_crcll(21),
      ADR3 => rx_input_memio_crcll(23),
      O => rx_input_memio_CHOICE2941_GROM
    );
  rx_input_memio_CHOICE2941_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE2941_GROM,
      O => rx_input_memio_CHOICE2941
    );
  mac_control_n001220_1_57 : X_LUT4
    generic map(
      INIT => X"CFCF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => clkslen,
      ADR3 => VCC,
      O => mac_control_n001220_1_GROM
    );
  mac_control_n001220_1_YUSED : X_BUF
    port map (
      I => mac_control_n001220_1_GROM,
      O => mac_control_n001220_1
    );
  rx_input_memio_crccomb_Mxor_CO_0_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(30),
      ADR1 => rx_input_memio_crcl(24),
      ADR2 => rx_input_memio_datal(7),
      ADR3 => rx_input_memio_datal(1),
      O => rx_input_memio_crcl_0_FROM
    );
  rx_input_memio_n0048_0_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_0_Q,
      O => rx_input_memio_n0048(0)
    );
  rx_input_memio_crcl_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_0_FROM,
      O => rx_input_memio_crc_0_Q
    );
  tx_fifocheck_fbbpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_3_FFY_RST
    );
  tx_fifocheck_fbbpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_3_FFY_RST,
      O => tx_fifocheck_fbbpl(2)
    );
  tx_fifocheck_fbbpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_5_FFY_RST
    );
  tx_fifocheck_fbbpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_5_FFY_RST,
      O => tx_fifocheck_fbbpl(4)
    );
  tx_fifocheck_fbbpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_7_FFY_RST
    );
  tx_fifocheck_fbbpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_7_FFY_RST,
      O => tx_fifocheck_fbbpl(6)
    );
  tx_fifocheck_fbbpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_9_FFY_RST
    );
  tx_fifocheck_fbbpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_9_FFY_RST,
      O => tx_fifocheck_fbbpl(8)
    );
  mac_control_phydo_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_11_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(10),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_11_FFY_RST,
      O => mac_control_phydo(10)
    );
  mac_control_phydo_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_13_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(12),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_13_FFY_RST,
      O => mac_control_phydo(12)
    );
  mac_control_phydo_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_15_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(14),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_15_FFY_RST,
      O => mac_control_phydo(14)
    );
  mac_control_Mmux_n0017_Result_29_42_SW0_1_58 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => mac_control_phyaddr(29),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_n0103,
      O => mac_control_Mmux_n0017_Result_29_42_SW0_1_FROM
    );
  mac_control_Mmux_n0017_Result_26_42_SW0_1_59 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyaddr(26),
      ADR2 => VCC,
      ADR3 => mac_control_n0103,
      O => mac_control_Mmux_n0017_Result_29_42_SW0_1_GROM
    );
  mac_control_Mmux_n0017_Result_29_42_SW0_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_29_42_SW0_1_FROM,
      O => mac_control_Mmux_n0017_Result_29_42_SW0_1
    );
  mac_control_Mmux_n0017_Result_29_42_SW0_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_29_42_SW0_1_GROM,
      O => mac_control_Mmux_n0017_Result_26_42_SW0_1
    );
  rx_input_fifo_fifo_BU408 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2424,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2434_FFY_RST,
      O => rx_input_fifo_fifo_N2434
    );
  rx_input_fifo_fifo_N2434_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2434_FFY_RST
    );
  tx_output_cs_Out1435_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_CHOICE1683,
      ADR1 => tx_output_cs_FFd11,
      ADR2 => tx_output_CHOICE1686,
      ADR3 => tx_output_CHOICE1679,
      O => tx_output_ltxen3_FROM
    );
  tx_output_cs_Out1435 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd14,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_cs_FFd13,
      ADR3 => tx_output_N81669,
      O => tx_output_ltxen
    );
  tx_output_ltxen3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_ltxen3_CEMUXNOT
    );
  tx_output_ltxen3_XUSED : X_BUF
    port map (
      I => tx_output_ltxen3_FROM,
      O => tx_output_N81669
    );
  mac_control_n00301 : X_LUT4
    generic map(
      INIT => X"2200"
    )
    port map (
      ADR0 => mac_control_N52143,
      ADR1 => mac_control_addr(0),
      ADR2 => VCC,
      ADR3 => mac_control_N52100,
      O => mac_control_n0030_FROM
    );
  mac_control_n00131 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_N52100,
      ADR3 => mac_control_N52132,
      O => mac_control_n0030_GROM
    );
  mac_control_n0030_XUSED : X_BUF
    port map (
      I => mac_control_n0030_FROM,
      O => mac_control_n0030
    );
  mac_control_n0030_YUSED : X_BUF
    port map (
      I => mac_control_n0030_GROM,
      O => mac_control_n0013
    );
  mac_control_n01031 : X_LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      ADR0 => mac_control_addr(4),
      ADR1 => mac_control_addr(2),
      ADR2 => mac_control_addr(3),
      ADR3 => mac_control_N52236,
      O => mac_control_n0103_FROM
    );
  mac_control_Mmux_n0017_Result_24_47_SW0 : X_LUT4
    generic map(
      INIT => X"FEEE"
    )
    port map (
      ADR0 => mac_control_CHOICE2186,
      ADR1 => mac_control_CHOICE2183,
      ADR2 => mac_control_phyaddr(24),
      ADR3 => mac_control_n0103,
      O => mac_control_n0103_GROM
    );
  mac_control_n0103_XUSED : X_BUF
    port map (
      I => mac_control_n0103_FROM,
      O => mac_control_n0103
    );
  mac_control_n0103_YUSED : X_BUF
    port map (
      I => mac_control_n0103_GROM,
      O => mac_control_N81789
    );
  mac_control_bitcnt_inst_sum_256_60 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_109_CYINIT,
      I1 => mac_control_bitcnt_inst_lut3_191,
      O => mac_control_bitcnt_inst_sum_256
    );
  mac_control_bitcnt_inst_lut3_1911 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_Mshreg_scslll_103,
      ADR2 => mac_control_bitcnt_109,
      ADR3 => VCC,
      O => mac_control_bitcnt_inst_lut3_191
    );
  mac_control_n00161 : X_LUT4
    generic map(
      INIT => X"5400"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => mac_control_sclkdelta,
      ADR2 => mac_control_Mshreg_scslll_103,
      ADR3 => clkslen,
      O => mac_control_bitcnt_109_GROM
    );
  mac_control_bitcnt_109_YUSED : X_BUF
    port map (
      I => mac_control_bitcnt_109_GROM,
      O => mac_control_n0016
    );
  mac_control_bitcnt_109_CYINIT_61 : X_BUF
    port map (
      I => mac_control_bitcnt_inst_cy_292,
      O => mac_control_bitcnt_109_CYINIT
    );
  mac_control_n00501 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => clkslen,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_rst,
      ADR3 => VCC,
      O => mac_control_n0050_GROM
    );
  mac_control_n0050_YUSED : X_BUF
    port map (
      I => mac_control_n0050_GROM,
      O => mac_control_n0050
    );
  mac_control_n00421 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => clkslen,
      ADR1 => mac_control_txf_rst,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_n0042_GROM
    );
  mac_control_n0042_YUSED : X_BUF
    port map (
      I => mac_control_n0042_GROM,
      O => mac_control_n0042
    );
  mac_control_n00511 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => clkslen,
      ADR3 => rxphyerrsr,
      O => mac_control_n0051_GROM
    );
  mac_control_n0051_YUSED : X_BUF
    port map (
      I => mac_control_n0051_GROM,
      O => mac_control_n0051
    );
  mac_control_n00431 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => clkslen,
      ADR3 => txfsr,
      O => mac_control_n0043_GROM
    );
  mac_control_n0043_YUSED : X_BUF
    port map (
      I => mac_control_n0043_GROM,
      O => mac_control_n0043
    );
  rx_input_fifo_fifo_BU382 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2403,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2423_FFX_RST,
      O => rx_input_fifo_fifo_N2423
    );
  rx_input_fifo_fifo_N2423_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2423_FFX_RST
    );
  mac_control_n00337 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_123,
      ADR1 => mac_control_phyrstcnt_121,
      ADR2 => mac_control_phyrstcnt_122,
      ADR3 => mac_control_phyrstcnt_124,
      O => mac_control_CHOICE2959_FROM
    );
  mac_control_n003310 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_119,
      ADR1 => mac_control_phyrstcnt_120,
      ADR2 => mac_control_phyrstcnt_110,
      ADR3 => mac_control_CHOICE2959,
      O => mac_control_CHOICE2959_GROM
    );
  mac_control_CHOICE2959_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2959_FROM,
      O => mac_control_CHOICE2959
    );
  mac_control_CHOICE2959_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2959_GROM,
      O => mac_control_CHOICE2960
    );
  mac_control_n00521 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => mac_control_rxoferr_rst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => clkslen,
      O => mac_control_n0052_GROM
    );
  mac_control_n0052_YUSED : X_BUF
    port map (
      I => mac_control_n0052_GROM,
      O => mac_control_n0052
    );
  mac_control_n00601 : X_LUT4
    generic map(
      INIT => X"5000"
    )
    port map (
      ADR0 => mac_control_bitcnt_109,
      ADR1 => VCC,
      ADR2 => mac_control_sclkdeltall,
      ADR3 => mac_control_N52138,
      O => mac_control_n0060_FROM
    );
  mac_control_Mmux_n0017_Result_26_77_1_62 : X_LUT4
    generic map(
      INIT => X"FF0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_dout(25),
      ADR3 => mac_control_n0060,
      O => mac_control_n0060_GROM
    );
  mac_control_n0060_XUSED : X_BUF
    port map (
      I => mac_control_n0060_FROM,
      O => mac_control_n0060
    );
  mac_control_n0060_YUSED : X_BUF
    port map (
      I => mac_control_n0060_GROM,
      O => mac_control_Mmux_n0017_Result_26_77_1
    );
  mac_control_din_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_15_FFY_RST
    );
  mac_control_din_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_15_FFY_RST,
      O => mac_control_din(14)
    );
  rx_input_fifo_fifo_BU388 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2400,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2420_FFX_RST,
      O => rx_input_fifo_fifo_N2420
    );
  rx_input_fifo_fifo_N2420_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2420_FFX_RST
    );
  mac_control_din_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_31_FFY_RST
    );
  mac_control_din_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(29),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_31_FFY_RST,
      O => mac_control_din(30)
    );
  mac_control_din_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_17_FFY_RST
    );
  mac_control_din_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_17_FFY_RST,
      O => mac_control_din(16)
    );
  mac_control_din_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_19_FFY_RST
    );
  mac_control_din_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(17),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_19_FFY_RST,
      O => mac_control_din(18)
    );
  mac_control_din_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_29_FFY_RST
    );
  mac_control_din_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(27),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_29_FFY_RST,
      O => mac_control_din(28)
    );
  rx_input_memio_crccomb_Mxor_n0021_Result1 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_datal(2),
      ADR2 => rx_input_memio_crcl(29),
      ADR3 => VCC,
      O => rx_input_memio_crccomb_n0118_0_FROM
    );
  rx_input_memio_crccomb_Mxor_n0007_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(29),
      ADR1 => rx_input_memio_crcl(25),
      ADR2 => rx_input_memio_datal(2),
      ADR3 => rx_input_memio_datal(6),
      O => rx_input_memio_crccomb_n0118_0_GROM
    );
  rx_input_memio_crccomb_n0118_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_n0118_0_FROM,
      O => rx_input_memio_crccomb_n0118(0)
    );
  rx_input_memio_crccomb_n0118_0_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_n0118_0_GROM,
      O => rx_input_memio_crccomb_Mxor_n0007_Xo(0)
    );
  mac_control_PHY_status_MII_Interface_n001124_2_63 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_mdccnt_33,
      ADR1 => mac_control_PHY_status_MII_Interface_mdccnt_32,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_mdccnt_34,
      O => mac_control_PHY_status_MII_Interface_n001124_2_GROM
    );
  mac_control_PHY_status_MII_Interface_n001124_2_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n001124_2_GROM,
      O => mac_control_PHY_status_MII_Interface_n001124_2
    );
  rx_input_fifo_fifo_BU476 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2399,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2439_FFX_RST,
      O => rx_input_fifo_fifo_N2439
    );
  rx_input_fifo_fifo_N2439_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2439_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_sout142_SW0 : X_LUT4
    generic map(
      INIT => X"F533"
    )
    port map (
      ADR0 => mac_control_PHY_status_miiaddr(0),
      ADR1 => mac_control_PHY_status_miiaddr(1),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(1),
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(0),
      O => mac_control_PHY_status_MII_Interface_N81705_FROM
    );
  mac_control_PHY_status_MII_Interface_sout142 : X_LUT4
    generic map(
      INIT => X"0020"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR3 => mac_control_PHY_status_MII_Interface_N81705,
      O => mac_control_PHY_status_MII_Interface_N81705_GROM
    );
  mac_control_PHY_status_MII_Interface_N81705_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81705_FROM,
      O => mac_control_PHY_status_MII_Interface_N81705
    );
  mac_control_PHY_status_MII_Interface_N81705_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81705_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2526
    );
  rx_input_memio_cs_FFd15_In_SW1 : X_LUT4
    generic map(
      INIT => X"1333"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => rx_input_memio_cs_FFd10,
      ADR2 => rx_input_memio_CHOICE1447,
      ADR3 => rx_input_memio_CHOICE1451,
      O => rx_input_memio_cs_FFd15_FROM
    );
  rx_input_memio_cs_FFd15_In_64 : X_LUT4
    generic map(
      INIT => X"A0B1"
    )
    port map (
      ADR0 => rx_input_invalid,
      ADR1 => rx_input_endf,
      ADR2 => rx_input_memio_cs_FFd15,
      ADR3 => rx_input_memio_N81863,
      O => rx_input_memio_cs_FFd15_In
    );
  rx_input_memio_cs_FFd15_XUSED : X_BUF
    port map (
      I => rx_input_memio_cs_FFd15_FROM,
      O => rx_input_memio_N81863
    );
  tx_output_crc_loigc_Mxor_CO_3_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0118(1),
      ADR1 => tx_output_crc_loigc_n0122(0),
      ADR2 => tx_output_crc_loigc_n0124(0),
      ADR3 => tx_output_crc_loigc_n0124(1),
      O => tx_output_crcl_3_FROM
    );
  tx_output_n0034_3_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_3_Q,
      O => tx_output_n0034(3)
    );
  tx_output_crcl_3_XUSED : X_BUF
    port map (
      I => tx_output_crcl_3_FROM,
      O => tx_output_crc_3_Q
    );
  rx_input_fifo_fifo_BU474 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2400,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2439_FFY_RST,
      O => rx_input_fifo_fifo_N2440
    );
  rx_input_fifo_fifo_N2439_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2439_FFY_RST
    );
  mac_control_PHY_status_n00151_1_65 : X_LUT4
    generic map(
      INIT => X"CCFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => clkslen,
      O => mac_control_PHY_status_n00151_1_GROM
    );
  mac_control_PHY_status_n00151_1_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_n00151_1_GROM,
      O => mac_control_PHY_status_n00151_1
    );
  mac_control_PHY_status_dout_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_3_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(2),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_3_FFY_RST,
      O => mac_control_PHY_status_dout(2)
    );
  mac_control_PHY_status_dout_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_5_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(4),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_5_FFY_RST,
      O => mac_control_PHY_status_dout(4)
    );
  mac_control_PHY_status_dout_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_7_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(6),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_7_FFY_RST,
      O => mac_control_PHY_status_dout(6)
    );
  mac_control_PHY_status_dout_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_9_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(8),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_9_FFY_RST,
      O => mac_control_PHY_status_dout(8)
    );
  mac_control_PHY_status_MII_Interface_sout273_SW1 : X_LUT4
    generic map(
      INIT => X"CECF"
    )
    port map (
      ADR0 => mac_control_PHY_status_din(14),
      ADR1 => mac_control_PHY_status_MII_Interface_CHOICE2546,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(4),
      O => mac_control_PHY_status_MII_Interface_N82067_FROM
    );
  mac_control_PHY_status_MII_Interface_sout273 : X_LUT4
    generic map(
      INIT => X"EFE0"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_CHOICE2532,
      ADR1 => mac_control_PHY_status_MII_Interface_N82069,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(1),
      ADR3 => mac_control_PHY_status_MII_Interface_N82067,
      O => mac_control_PHY_status_MII_Interface_N82067_GROM
    );
  mac_control_PHY_status_MII_Interface_N82067_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N82067_FROM,
      O => mac_control_PHY_status_MII_Interface_N82067
    );
  mac_control_PHY_status_MII_Interface_N82067_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N82067_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2555
    );
  rx_input_memio_bpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_13_FFY_RST
    );
  rx_input_memio_bpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(12),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_13_FFY_RST,
      O => rx_input_memio_bpl(12)
    );
  rx_input_memio_cs_FFd16_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_RESET_1,
      O => rx_input_memio_cs_FFd16_FFY_SET
    );
  rx_input_memio_cs_FFd16_66 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_memio_cs_FFd16_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_memio_cs_FFd16_FFY_SET,
      RST => GND,
      O => rx_input_memio_cs_FFd16
    );
  rx_input_memio_cs_FFd16_In_SW0 : X_LUT4
    generic map(
      INIT => X"FFDF"
    )
    port map (
      ADR0 => rx_input_memio_CHOICE1451,
      ADR1 => rx_input_endf,
      ADR2 => rx_input_memio_CHOICE1447,
      ADR3 => rx_input_invalid,
      O => rx_input_memio_cs_FFd16_FROM
    );
  rx_input_memio_cs_FFd16_In_67 : X_LUT4
    generic map(
      INIT => X"FEFA"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd3,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => rx_input_memio_cs_FFd1,
      ADR3 => rx_input_memio_N70785,
      O => rx_input_memio_cs_FFd16_In
    );
  rx_input_memio_cs_FFd16_XUSED : X_BUF
    port map (
      I => rx_input_memio_cs_FFd16_FROM,
      O => rx_input_memio_N70785
    );
  rx_input_fifo_fifo_BU417 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2421,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2431_FFX_RST,
      O => rx_input_fifo_fifo_N2431
    );
  rx_input_fifo_fifo_N2431_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2431_FFX_RST
    );
  mac_control_Mmux_n0017_Result_18_42_SW0_1_68 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => mac_control_phyaddr(18),
      ADR1 => VCC,
      ADR2 => mac_control_n0103,
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_18_42_SW0_1_FROM
    );
  mac_control_Mmux_n0017_Result_20_42_SW0_1_69 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => mac_control_n0103,
      ADR1 => mac_control_phyaddr(20),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_18_42_SW0_1_GROM
    );
  mac_control_Mmux_n0017_Result_18_42_SW0_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_18_42_SW0_1_FROM,
      O => mac_control_Mmux_n0017_Result_18_42_SW0_1
    );
  mac_control_Mmux_n0017_Result_18_42_SW0_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_18_42_SW0_1_GROM,
      O => mac_control_Mmux_n0017_Result_20_42_SW0_1
    );
  rx_input_fifo_RESET_1_70 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => RESET_IBUF_2,
      O => rx_input_fifo_RESET_1_GROM
    );
  rx_input_fifo_RESET_1_YUSED : X_BUF
    port map (
      I => rx_input_fifo_RESET_1_GROM,
      O => rx_input_fifo_RESET_1
    );
  rxf_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxf_CEMUXNOT
    );
  mac_control_phyaddr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_3_FFY_RST
    );
  mac_control_phyaddr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_3_FFY_RST,
      O => mac_control_phyaddr(2)
    );
  mac_control_phyaddr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_5_FFY_RST
    );
  mac_control_phyaddr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_5_FFY_RST,
      O => mac_control_phyaddr(4)
    );
  mac_control_phyaddr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_7_FFY_RST
    );
  mac_control_phyaddr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_7_FFY_RST,
      O => mac_control_phyaddr(6)
    );
  mac_control_phyaddr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_9_FFY_RST
    );
  mac_control_phyaddr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_9_FFY_RST,
      O => mac_control_phyaddr(8)
    );
  slowclock_rxoferrl_71 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_rxoferrl_GROM,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => rxoferr,
      SRST => slowclock_rxoferrl_LOGIC_ZERO,
      O => slowclock_rxoferrl
    );
  slowclock_rxoferrl_LOGIC_ZERO_72 : X_ZERO
    port map (
      O => slowclock_rxoferrl_LOGIC_ZERO
    );
  slowclock_rxoferrl_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => slowclock_rxoferrl_GROM
    );
  rx_input_memio_crcrst_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcrst_CEMUXNOT
    );
  rx_input_memio_dout_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_1_FFY_RST
    );
  rx_input_memio_dout_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_1_FFY_RST,
      O => rx_input_memio_dout(0)
    );
  txfbbp_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_11_FFY_RST
    );
  tx_output_FBBP_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(10),
      CE => txfbbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_11_FFY_RST,
      O => txfbbp(10)
    );
  txfbbp_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => txfbbp_11_CEMUXNOT
    );
  rx_input_memio_dout_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_3_FFY_RST
    );
  rx_input_memio_dout_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_3_FFY_RST,
      O => rx_input_memio_dout(2)
    );
  txfbbp_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_13_FFY_RST
    );
  tx_output_FBBP_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(12),
      CE => txfbbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_13_FFY_RST,
      O => txfbbp(12)
    );
  txfbbp_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => txfbbp_13_CEMUXNOT
    );
  txfbbp_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_15_FFY_RST
    );
  tx_output_FBBP_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(14),
      CE => txfbbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_15_FFY_RST,
      O => txfbbp(14)
    );
  txfbbp_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => txfbbp_15_CEMUXNOT
    );
  rx_input_memio_dout_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_7_FFY_RST
    );
  rx_input_memio_dout_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_7_FFY_RST,
      O => rx_input_memio_dout(6)
    );
  rx_input_memio_dout_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_9_FFY_RST
    );
  rx_input_memio_dout_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_9_FFY_RST,
      O => rx_input_memio_dout(8)
    );
  mac_control_PHY_status_MII_Interface_Ker372431 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => clkslen,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_N37245_FROM
    );
  mac_control_PHY_status_MII_Interface_n00101 : X_LUT4
    generic map(
      INIT => X"AE00"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => MDC_OBUF,
      ADR2 => mac_control_PHY_status_MII_Interface_mdccnt_37,
      ADR3 => mac_control_PHY_status_MII_Interface_N37245,
      O => mac_control_PHY_status_MII_Interface_N37245_GROM
    );
  mac_control_PHY_status_MII_Interface_N37245_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N37245_FROM,
      O => mac_control_PHY_status_MII_Interface_N37245
    );
  mac_control_PHY_status_MII_Interface_N37245_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N37245_GROM,
      O => mac_control_PHY_status_MII_Interface_n0010
    );
  mac_control_PHY_status_MII_Interface_Ker372381 : X_LUT4
    generic map(
      INIT => X"8800"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(1),
      O => mac_control_PHY_status_MII_Interface_N37240_FROM
    );
  mac_control_PHY_status_MII_Interface_sout312 : X_LUT4
    generic map(
      INIT => X"B800"
    )
    port map (
      ADR0 => mac_control_PHY_status_din(0),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR2 => mac_control_PHY_status_din(8),
      ADR3 => mac_control_PHY_status_MII_Interface_N37240,
      O => mac_control_PHY_status_MII_Interface_N37240_GROM
    );
  mac_control_PHY_status_MII_Interface_N37240_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N37240_FROM,
      O => mac_control_PHY_status_MII_Interface_N37240
    );
  mac_control_PHY_status_MII_Interface_N37240_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N37240_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2562
    );
  tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2_73 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => tx_output_data(0),
      ADR1 => VCC,
      ADR2 => tx_output_crcl(22),
      ADR3 => tx_output_crcl(31),
      O => tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2_FROM
    );
  tx_output_crc_loigc_Mxor_CO_18_Xo_2_1_2_74 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => tx_output_data(0),
      ADR1 => tx_output_crcl(31),
      ADR2 => VCC,
      ADR3 => tx_output_crcl(10),
      O => tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2_GROM
    );
  tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2_FROM,
      O => tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2
    );
  tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2_GROM,
      O => tx_output_crc_loigc_Mxor_CO_18_Xo_2_1_2
    );
  tx_output_TXF1 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_ltxen3,
      ADR2 => tx_output_ltxen2,
      ADR3 => VCC,
      O => txf_GROM
    );
  txf_YUSED : X_BUF
    port map (
      I => txf_GROM,
      O => txf
    );
  rx_input_fifo_control_ldata_1_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d1(1),
      ADR1 => rx_input_fifo_control_cs_FFd1,
      ADR2 => rx_input_fifo_control_cs_FFd2,
      ADR3 => rx_input_fifo_control_d0(1),
      O => rx_input_fifo_control_CHOICE1462_FROM
    );
  rx_input_fifo_control_ldata_0_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_d0(0),
      ADR1 => rx_input_fifo_control_cs_FFd1,
      ADR2 => rx_input_fifo_control_d1(0),
      ADR3 => rx_input_fifo_control_cs_FFd2,
      O => rx_input_fifo_control_CHOICE1462_GROM
    );
  rx_input_fifo_control_CHOICE1462_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1462_FROM,
      O => rx_input_fifo_control_CHOICE1462
    );
  rx_input_fifo_control_CHOICE1462_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1462_GROM,
      O => rx_input_fifo_control_CHOICE1455
    );
  rx_input_fifo_fifo_BU454 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N4,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2469_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2469
    );
  rx_input_fifo_fifo_N2469_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2469_FFX_SET
    );
  rx_input_fifo_control_ldata_0_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_d2(0),
      ADR1 => rx_input_fifo_control_cs_FFd3,
      ADR2 => rx_input_fifo_control_cs_FFd4,
      ADR3 => rx_input_fifo_control_d3(0),
      O => rx_input_data_0_FROM
    );
  rx_input_fifo_control_ldata_0_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1455,
      ADR3 => rx_input_fifo_control_CHOICE1458,
      O => rx_input_fifo_control_ldata(0)
    );
  rx_input_data_0_XUSED : X_BUF
    port map (
      I => rx_input_data_0_FROM,
      O => rx_input_fifo_control_CHOICE1458
    );
  rx_output_Ker331051 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_cs_FFd11,
      ADR2 => rx_output_cs_FFd1,
      ADR3 => VCC,
      O => rx_output_cs_FFd9_FROM
    );
  rx_output_cs_FFd9_In1 : X_LUT4
    generic map(
      INIT => X"88A8"
    )
    port map (
      ADR0 => rx_output_nf,
      ADR1 => rx_output_N33107,
      ADR2 => rx_output_cs_FFd5,
      ADR3 => rx_output_n0018,
      O => rx_output_cs_FFd9_In
    );
  rx_output_cs_FFd9_XUSED : X_BUF
    port map (
      I => rx_output_cs_FFd9_FROM,
      O => rx_output_N33107
    );
  rx_input_fifo_control_ldata_7_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd1,
      ADR1 => rx_input_fifo_control_d1(7),
      ADR2 => rx_input_fifo_control_cs_FFd2,
      ADR3 => rx_input_fifo_control_d0(7),
      O => rx_input_fifo_control_CHOICE1483_FROM
    );
  rx_input_fifo_control_ldata_2_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd1,
      ADR1 => rx_input_fifo_control_d0(2),
      ADR2 => rx_input_fifo_control_cs_FFd2,
      ADR3 => rx_input_fifo_control_d1(2),
      O => rx_input_fifo_control_CHOICE1483_GROM
    );
  rx_input_fifo_control_CHOICE1483_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1483_FROM,
      O => rx_input_fifo_control_CHOICE1483
    );
  rx_input_fifo_control_CHOICE1483_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1483_GROM,
      O => rx_input_fifo_control_CHOICE1518
    );
  rx_input_fifo_control_ldata_1_9 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd3,
      ADR1 => rx_input_fifo_control_cs_FFd4,
      ADR2 => rx_input_fifo_control_d2(1),
      ADR3 => rx_input_fifo_control_d3(1),
      O => rx_input_data_1_FROM
    );
  rx_input_fifo_control_ldata_1_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1462,
      ADR3 => rx_input_fifo_control_CHOICE1465,
      O => rx_input_fifo_control_ldata(1)
    );
  rx_input_data_1_XUSED : X_BUF
    port map (
      I => rx_input_data_1_FROM,
      O => rx_input_fifo_control_CHOICE1465
    );
  tx_output_n000724 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcnt_45,
      ADR1 => tx_output_bcnt_43,
      ADR2 => tx_output_bcnt_44,
      ADR3 => tx_output_bcnt_42,
      O => tx_output_CHOICE1656_GROM
    );
  tx_output_CHOICE1656_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1656_GROM,
      O => tx_output_CHOICE1656
    );
  rx_input_fifo_control_ldata_6_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d0(6),
      ADR1 => rx_input_fifo_control_cs_FFd2,
      ADR2 => rx_input_fifo_control_d1(6),
      ADR3 => rx_input_fifo_control_cs_FFd1,
      O => rx_input_fifo_control_CHOICE1490_FROM
    );
  rx_input_fifo_control_ldata_3_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd2,
      ADR1 => rx_input_fifo_control_cs_FFd1,
      ADR2 => rx_input_fifo_control_d0(3),
      ADR3 => rx_input_fifo_control_d1(3),
      O => rx_input_fifo_control_CHOICE1490_GROM
    );
  rx_input_fifo_control_CHOICE1490_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1490_FROM,
      O => rx_input_fifo_control_CHOICE1490
    );
  rx_input_fifo_control_CHOICE1490_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1490_GROM,
      O => rx_input_fifo_control_CHOICE1511
    );
  rx_input_fifo_control_ldata_2_9 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d2(2),
      ADR1 => rx_input_fifo_control_d3(2),
      ADR2 => rx_input_fifo_control_cs_FFd4,
      ADR3 => rx_input_fifo_control_cs_FFd3,
      O => rx_input_data_2_FROM
    );
  rx_input_fifo_control_ldata_2_10 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_control_CHOICE1518,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_control_CHOICE1521,
      O => rx_input_fifo_control_ldata(2)
    );
  rx_input_data_2_XUSED : X_BUF
    port map (
      I => rx_input_data_2_FROM,
      O => rx_input_fifo_control_CHOICE1521
    );
  tx_output_n000761 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcnt_51,
      ADR1 => tx_output_bcnt_53,
      ADR2 => tx_output_bcnt_52,
      ADR3 => tx_output_bcnt_50,
      O => tx_output_CHOICE1671_FROM
    );
  tx_output_n000774_SW0 : X_LUT4
    generic map(
      INIT => X"BFFF"
    )
    port map (
      ADR0 => tx_output_bcnt_41,
      ADR1 => tx_output_CHOICE1656,
      ADR2 => tx_output_CHOICE1664,
      ADR3 => tx_output_CHOICE1671,
      O => tx_output_CHOICE1671_GROM
    );
  tx_output_CHOICE1671_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1671_FROM,
      O => tx_output_CHOICE1671
    );
  tx_output_CHOICE1671_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1671_GROM,
      O => tx_output_N81677
    );
  rx_input_fifo_control_cs_FFd4_In_2_75 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd1,
      ADR1 => rx_input_fifo_control_cs_FFd4,
      ADR2 => rx_input_fifo_control_cs_FFd2,
      ADR3 => rx_input_fifo_control_cs_FFd3,
      O => rx_input_fifo_control_cs_FFd4_In_2_FROM
    );
  rx_input_fifo_control_ldata_4_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd2,
      ADR1 => rx_input_fifo_control_d0(4),
      ADR2 => rx_input_fifo_control_d1(4),
      ADR3 => rx_input_fifo_control_cs_FFd1,
      O => rx_input_fifo_control_cs_FFd4_In_2_GROM
    );
  rx_input_fifo_control_cs_FFd4_In_2_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_cs_FFd4_In_2_FROM,
      O => rx_input_fifo_control_cs_FFd4_In_2
    );
  rx_input_fifo_control_cs_FFd4_In_2_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_cs_FFd4_In_2_GROM,
      O => rx_input_fifo_control_CHOICE1497
    );
  rx_input_fifo_control_ldata_3_9 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d3(3),
      ADR1 => rx_input_fifo_control_cs_FFd3,
      ADR2 => rx_input_fifo_control_d2(3),
      ADR3 => rx_input_fifo_control_cs_FFd4,
      O => rx_input_data_3_FROM
    );
  rx_input_fifo_control_ldata_3_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1511,
      ADR3 => rx_input_fifo_control_CHOICE1514,
      O => rx_input_fifo_control_ldata(3)
    );
  rx_input_data_3_XUSED : X_BUF
    port map (
      I => rx_input_data_3_FROM,
      O => rx_input_fifo_control_CHOICE1514
    );
  tx_output_n000748 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcnt_46,
      ADR1 => tx_output_bcnt_47,
      ADR2 => tx_output_bcnt_48,
      ADR3 => tx_output_bcnt_49,
      O => tx_output_CHOICE1664_GROM
    );
  tx_output_CHOICE1664_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1664_GROM,
      O => tx_output_CHOICE1664
    );
  rx_input_fifo_control_ldata_8_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_d1(8),
      ADR1 => rx_input_fifo_control_cs_FFd2,
      ADR2 => rx_input_fifo_control_d0(8),
      ADR3 => rx_input_fifo_control_cs_FFd1,
      O => rx_input_fifo_control_CHOICE1476_FROM
    );
  rx_input_fifo_control_ldata_5_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd2,
      ADR1 => rx_input_fifo_control_cs_FFd1,
      ADR2 => rx_input_fifo_control_d1(5),
      ADR3 => rx_input_fifo_control_d0(5),
      O => rx_input_fifo_control_CHOICE1476_GROM
    );
  rx_input_fifo_control_CHOICE1476_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1476_FROM,
      O => rx_input_fifo_control_CHOICE1476
    );
  rx_input_fifo_control_CHOICE1476_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1476_GROM,
      O => rx_input_fifo_control_CHOICE1504
    );
  rx_input_fifo_control_ldata_4_9 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d2(4),
      ADR1 => rx_input_fifo_control_d3(4),
      ADR2 => rx_input_fifo_control_cs_FFd4,
      ADR3 => rx_input_fifo_control_cs_FFd3,
      O => rx_input_data_4_FROM
    );
  rx_input_fifo_control_ldata_4_10 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_control_CHOICE1497,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_control_CHOICE1500,
      O => rx_input_fifo_control_ldata(4)
    );
  rx_input_data_4_XUSED : X_BUF
    port map (
      I => rx_input_data_4_FROM,
      O => rx_input_fifo_control_CHOICE1500
    );
  rx_input_fifo_fifo_BU568 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2449_GROM,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2449_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2450
    );
  rx_input_fifo_fifo_N2449_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2449_FFY_SET
    );
  rx_input_fifo_control_ldata_5_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_d3(5),
      ADR1 => rx_input_fifo_control_cs_FFd4,
      ADR2 => rx_input_fifo_control_cs_FFd3,
      ADR3 => rx_input_fifo_control_d2(5),
      O => rx_input_data_5_FROM
    );
  rx_input_fifo_control_ldata_5_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1504,
      ADR3 => rx_input_fifo_control_CHOICE1507,
      O => rx_input_fifo_control_ldata(5)
    );
  rx_input_data_5_XUSED : X_BUF
    port map (
      I => rx_input_data_5_FROM,
      O => rx_input_fifo_control_CHOICE1507
    );
  rx_input_fifo_control_ldata_6_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_d2(6),
      ADR1 => rx_input_fifo_control_cs_FFd3,
      ADR2 => rx_input_fifo_control_cs_FFd4,
      ADR3 => rx_input_fifo_control_d3(6),
      O => rx_input_data_6_FROM
    );
  rx_input_fifo_control_ldata_6_10 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_control_CHOICE1490,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_control_CHOICE1493,
      O => rx_input_fifo_control_ldata(6)
    );
  rx_input_data_6_XUSED : X_BUF
    port map (
      I => rx_input_data_6_FROM,
      O => rx_input_fifo_control_CHOICE1493
    );
  rx_input_fifo_control_ldata_7_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_d3(7),
      ADR1 => rx_input_fifo_control_cs_FFd4,
      ADR2 => rx_input_fifo_control_cs_FFd3,
      ADR3 => rx_input_fifo_control_d2(7),
      O => rx_input_data_7_FROM
    );
  rx_input_fifo_control_ldata_7_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1483,
      ADR3 => rx_input_fifo_control_CHOICE1486,
      O => rx_input_fifo_control_ldata(7)
    );
  rx_input_data_7_XUSED : X_BUF
    port map (
      I => rx_input_data_7_FROM,
      O => rx_input_fifo_control_CHOICE1486
    );
  rx_input_fifo_control_ldata_9_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd2,
      ADR1 => rx_input_fifo_control_d1(9),
      ADR2 => rx_input_fifo_control_d0(9),
      ADR3 => rx_input_fifo_control_cs_FFd1,
      O => rx_input_fifo_control_CHOICE1469_GROM
    );
  rx_input_fifo_control_CHOICE1469_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1469_GROM,
      O => rx_input_fifo_control_CHOICE1469
    );
  rx_input_fifo_control_ldata_8_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_d2(8),
      ADR1 => rx_input_fifo_control_cs_FFd3,
      ADR2 => rx_input_fifo_control_d3(8),
      ADR3 => rx_input_fifo_control_cs_FFd4,
      O => rx_input_endf_FROM
    );
  rx_input_fifo_control_ldata_8_10 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_fifo_control_CHOICE1476,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_control_CHOICE1479,
      O => rx_input_fifo_control_ldata(8)
    );
  rx_input_endf_XUSED : X_BUF
    port map (
      I => rx_input_endf_FROM,
      O => rx_input_fifo_control_CHOICE1479
    );
  rx_input_fifo_control_ldata_9_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd3,
      ADR1 => rx_input_fifo_control_d2(9),
      ADR2 => rx_input_fifo_control_d3(9),
      ADR3 => rx_input_fifo_control_cs_FFd4,
      O => rx_input_invalid_FROM
    );
  rx_input_fifo_control_ldata_9_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1469,
      ADR3 => rx_input_fifo_control_CHOICE1472,
      O => rx_input_fifo_control_ldata(9)
    );
  rx_input_invalid_XUSED : X_BUF
    port map (
      I => rx_input_invalid_FROM,
      O => rx_input_fifo_control_CHOICE1472
    );
  mac_control_PHY_status_MII_Interface_sts28_SW0 : X_LUT4
    generic map(
      INIT => X"77FF"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(1),
      O => mac_control_PHY_status_MII_Interface_N81600_FROM
    );
  mac_control_PHY_status_MII_Interface_n0079_SW0 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(5),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(1),
      O => mac_control_PHY_status_MII_Interface_N81600_GROM
    );
  mac_control_PHY_status_MII_Interface_N81600_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81600_FROM,
      O => mac_control_PHY_status_MII_Interface_N81600
    );
  mac_control_PHY_status_MII_Interface_N81600_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81600_GROM,
      O => mac_control_PHY_status_MII_Interface_N69488
    );
  rx_input_memio_addrchk_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"4450"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => rx_input_memio_addrchk_cs_FFd3,
      ADR2 => rx_input_memio_addrchk_cs_FFd2,
      ADR3 => rx_input_memio_brdy,
      O => rx_input_memio_addrchk_cs_FFd2_In
    );
  rx_input_memio_addrchk_cs_FFd6_In10 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd4,
      ADR1 => rx_input_memio_addrchk_cs_FFd2,
      ADR2 => rx_input_memio_addrchk_cs_FFd1,
      ADR3 => rx_input_memio_addrchk_cs_FFd3,
      O => rx_input_memio_addrchk_cs_FFd2_GROM
    );
  rx_input_memio_addrchk_cs_FFd2_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_cs_FFd2_GROM,
      O => rx_input_memio_addrchk_CHOICE1550
    );
  tx_output_crc_loigc_Mxor_CO_6_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0115(0),
      ADR1 => tx_output_crc_loigc_n0124(0),
      ADR2 => tx_output_crc_loigc_Mxor_n0007_Xo(0),
      ADR3 => tx_output_crc_loigc_Mxor_CO_18_Xo(0),
      O => tx_output_crcl_6_FROM
    );
  tx_output_n0034_6_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16,
      ADR2 => VCC,
      ADR3 => tx_output_crc_6_Q,
      O => tx_output_n0034(6)
    );
  tx_output_crcl_6_XUSED : X_BUF
    port map (
      I => tx_output_crcl_6_FROM,
      O => tx_output_crc_6_Q
    );
  rx_input_memio_addrchk_cs_FFd6_In13 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd7,
      ADR1 => rx_input_memio_addrchk_CHOICE1550,
      ADR2 => rx_input_memio_addrchk_cs_FFd5,
      ADR3 => rx_input_memio_addrchk_cs_FFd6,
      O => rx_input_memio_addrchk_cs_FFd6_FROM
    );
  rx_input_memio_addrchk_cs_FFd6_In27 : X_LUT4
    generic map(
      INIT => X"F444"
    )
    port map (
      ADR0 => rx_input_memio_brdy,
      ADR1 => rx_input_memio_addrchk_cs_FFd6,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => rx_input_memio_addrchk_CHOICE1551,
      O => rx_input_memio_addrchk_cs_FFd6_In
    );
  rx_input_memio_addrchk_cs_FFd6_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_cs_FFd6_FROM,
      O => rx_input_memio_addrchk_CHOICE1551
    );
  rx_input_memio_crccomb_Mxor_CO_7_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(24),
      ADR1 => rx_input_memio_crcl(27),
      ADR2 => rx_input_memio_datal(4),
      ADR3 => rx_input_memio_datal(7),
      O => rx_input_memio_crccomb_Mxor_CO_7_Xo_1_FROM
    );
  rx_input_memio_crccomb_Mxor_CO_4_Xo_1_1_2_76 : X_LUT4
    generic map(
      INIT => X"9696"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0118(1),
      ADR1 => rx_input_memio_datal(4),
      ADR2 => rx_input_memio_crcl(27),
      ADR3 => VCC,
      O => rx_input_memio_crccomb_Mxor_CO_7_Xo_1_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_7_Xo_1_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_7_Xo_1_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_7_Xo(1)
    );
  rx_input_memio_crccomb_Mxor_CO_7_Xo_1_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_7_Xo_1_GROM,
      O => rx_input_memio_crccomb_Mxor_CO_4_Xo_1_1_2
    );
  mac_control_Ker52151 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_N52220,
      ADR1 => mac_control_addr(7),
      ADR2 => mac_control_N69420,
      ADR3 => mac_control_newcmd,
      O => mac_control_N52153_FROM
    );
  mac_control_n00341 : X_LUT4
    generic map(
      INIT => X"000C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => clkslen,
      ADR2 => RESET_IBUF,
      ADR3 => mac_control_N52153,
      O => mac_control_N52153_GROM
    );
  mac_control_N52153_XUSED : X_BUF
    port map (
      I => mac_control_N52153_FROM,
      O => mac_control_N52153
    );
  mac_control_N52153_YUSED : X_BUF
    port map (
      I => mac_control_N52153_GROM,
      O => mac_control_n0034
    );
  mac_control_Ker52136 : X_LUT4
    generic map(
      INIT => X"0044"
    )
    port map (
      ADR0 => mac_control_Ker52136_2,
      ADR1 => mac_control_bitcnt_107,
      ADR2 => VCC,
      ADR3 => mac_control_bitcnt_108,
      O => mac_control_N52138_FROM
    );
  mac_control_n001220 : X_LUT4
    generic map(
      INIT => X"2322"
    )
    port map (
      ADR0 => mac_control_CHOICE1171,
      ADR1 => mac_control_n001220_1,
      ADR2 => mac_control_n001220_SW0_1,
      ADR3 => mac_control_N52138,
      O => mac_control_N52138_GROM
    );
  mac_control_N52138_XUSED : X_BUF
    port map (
      I => mac_control_N52138_FROM,
      O => mac_control_N52138
    );
  mac_control_N52138_YUSED : X_BUF
    port map (
      I => mac_control_N52138_GROM,
      O => mac_control_N70898
    );
  mac_control_PHY_status_MII_Interface_n0004_77 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR2 => mac_control_PHY_status_MII_Interface_n0004_2,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(1),
      O => mac_control_PHY_status_MII_Interface_cs_FFd2_FROM
    );
  mac_control_PHY_status_MII_Interface_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd3,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_n0004,
      O => mac_control_PHY_status_MII_Interface_cs_FFd2_In
    );
  mac_control_PHY_status_MII_Interface_cs_FFd2_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd2_FROM,
      O => mac_control_PHY_status_MII_Interface_n0004
    );
  rx_input_fifo_fifo_BU276 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3940,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N7_FFY_RST,
      O => rx_input_fifo_fifo_N6
    );
  rx_input_fifo_fifo_N7_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N7_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_n0079_78 : X_LUT4
    generic map(
      INIT => X"1555"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR3 => mac_control_PHY_status_MII_Interface_N69488,
      O => mac_control_PHY_status_MII_Interface_statecnt_1_FROM
    );
  mac_control_PHY_status_MII_Interface_n0014_1_1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_n0078(1),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_n0079,
      O => mac_control_PHY_status_MII_Interface_n0014(1)
    );
  mac_control_PHY_status_MII_Interface_statecnt_1_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_statecnt_1_FROM,
      O => mac_control_PHY_status_MII_Interface_n0079
    );
  rx_input_fifo_fifo_BU343 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N4570,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2482_FFY_RST,
      O => rx_input_fifo_fifo_N2481
    );
  rx_input_fifo_fifo_N2482_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2482_FFY_RST
    );
  rx_input_fifo_fifo_BU570 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N5348,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2449_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2449
    );
  rx_input_fifo_fifo_N2449_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2449_FFX_SET
    );
  macaddr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_3_FFY_RST
    );
  mac_control_MACADDR_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(2),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_3_FFY_RST,
      O => macaddr(2)
    );
  macaddr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_5_FFY_RST
    );
  mac_control_MACADDR_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(4),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_5_FFY_RST,
      O => macaddr(4)
    );
  macaddr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_7_FFY_RST
    );
  mac_control_MACADDR_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(6),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_7_FFY_RST,
      O => macaddr(6)
    );
  macaddr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_9_FFY_RST
    );
  mac_control_MACADDR_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(8),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_9_FFY_RST,
      O => macaddr(8)
    );
  rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_2_79 : X_LUT4
    generic map(
      INIT => X"9696"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0115(0),
      ADR1 => rx_input_memio_crccomb_n0104(0),
      ADR2 => rx_input_memio_crcl(4),
      ADR3 => VCC,
      O => rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_2_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_2_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_2_GROM,
      O => rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_2
    );
  tx_input_Ker344911 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF_1,
      ADR2 => tx_input_den,
      ADR3 => VCC,
      O => tx_input_N34493_FROM
    );
  tx_input_n00201 : X_LUT4
    generic map(
      INIT => X"CCC8"
    )
    port map (
      ADR0 => tx_input_cs_FFd10,
      ADR1 => tx_input_N34493,
      ADR2 => tx_input_cs_FFd11,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_N34493_GROM
    );
  tx_input_N34493_XUSED : X_BUF
    port map (
      I => tx_input_N34493_FROM,
      O => tx_input_N34493
    );
  tx_input_N34493_YUSED : X_BUF
    port map (
      I => tx_input_N34493_GROM,
      O => tx_input_n0020
    );
  rx_output_n0043_SW0 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => rx_output_cs_FFd1,
      ADR1 => rx_output_cs_FFd11,
      ADR2 => VCC,
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_N69253_FROM
    );
  rx_output_n0043_80 : X_LUT4
    generic map(
      INIT => X"5554"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => rx_output_cs_FFd5,
      ADR2 => rx_output_cs_FFd17,
      ADR3 => rx_output_N69253,
      O => rx_output_N69253_GROM
    );
  rx_output_N69253_XUSED : X_BUF
    port map (
      I => rx_output_N69253_FROM,
      O => rx_output_N69253
    );
  rx_output_N69253_YUSED : X_BUF
    port map (
      I => rx_output_N69253_GROM,
      O => rx_output_n0043
    );
  tx_output_crc_loigc_Mxor_n0001_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_data(7),
      ADR3 => tx_output_crcl(24),
      O => tx_output_crc_loigc_n0122_1_FROM
    );
  tx_output_crc_loigc_Mxor_CO_7_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(24),
      ADR1 => tx_output_data(4),
      ADR2 => tx_output_crcl(27),
      ADR3 => tx_output_data(7),
      O => tx_output_crc_loigc_n0122_1_GROM
    );
  tx_output_crc_loigc_n0122_1_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0122_1_FROM,
      O => tx_output_crc_loigc_n0122(1)
    );
  tx_output_crc_loigc_n0122_1_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0122_1_GROM,
      O => tx_output_crc_loigc_Mxor_CO_7_Xo(1)
    );
  tx_output_crc_loigc_Mxor_CO_7_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_Mxor_CO_7_Xo(1),
      ADR1 => tx_output_crc_loigc_n0118(1),
      ADR2 => tx_output_crc_loigc_n0124(0),
      ADR3 => tx_output_crc_loigc_n0118(0),
      O => tx_output_crcl_7_FROM
    );
  tx_output_n0034_7_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_7_Q,
      O => tx_output_n0034(7)
    );
  tx_output_crcl_7_XUSED : X_BUF
    port map (
      I => tx_output_crcl_7_FROM,
      O => tx_output_crc_7_Q
    );
  mac_control_PHY_status_din_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_3_FFY_RST
    );
  mac_control_PHY_status_din_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(2),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_3_FFY_RST,
      O => mac_control_PHY_status_din(2)
    );
  mac_control_PHY_status_din_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_5_FFY_RST
    );
  mac_control_PHY_status_din_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(4),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_5_FFY_RST,
      O => mac_control_PHY_status_din(4)
    );
  mac_control_PHY_status_din_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_7_FFY_RST
    );
  mac_control_PHY_status_din_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(6),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_7_FFY_RST,
      O => mac_control_PHY_status_din(6)
    );
  rx_input_fifo_fifo_BU411 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2423,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2432_FFY_RST,
      O => rx_input_fifo_fifo_N2433
    );
  rx_input_fifo_fifo_N2432_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2432_FFY_RST
    );
  mac_control_PHY_status_din_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_9_FFY_RST
    );
  mac_control_PHY_status_din_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(8),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_9_FFY_RST,
      O => mac_control_PHY_status_din(8)
    );
  mac_control_Mmux_n0017_Result_5_107_SW0 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phyaddr(5),
      ADR1 => mac_control_rxfifowerr_cnt(5),
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_N52132,
      O => mac_control_N82133_FROM
    );
  mac_control_Mmux_n0017_Result_10_107_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(10),
      ADR1 => mac_control_phyaddr(10),
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_N52132,
      O => mac_control_N82133_GROM
    );
  mac_control_N82133_XUSED : X_BUF
    port map (
      I => mac_control_N82133_FROM,
      O => mac_control_N82133
    );
  mac_control_N82133_YUSED : X_BUF
    port map (
      I => mac_control_N82133_GROM,
      O => mac_control_N82121
    );
  rx_input_fifo_fifo_BU336 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N4530,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2482_FFX_RST,
      O => rx_input_fifo_fifo_N2482
    );
  rx_input_fifo_fifo_N2482_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2482_FFX_RST
    );
  rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2_81 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => rx_input_memio_datal(1),
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcl(30),
      ADR3 => rx_input_memio_crcl(15),
      O => rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2_FROM
    );
  rx_input_memio_crccomb_Mxor_n0000_Result1 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_memio_datal(1),
      ADR1 => rx_input_memio_crcl(30),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2
    );
  rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2_GROM,
      O => rx_input_memio_crccomb_n0104(0)
    );
  mac_control_Mmux_n0017_Result_25_42_SW0_1_82 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => mac_control_phyaddr(25),
      ADR1 => mac_control_n0103,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_25_42_SW0_1_FROM
    );
  mac_control_Mmux_n0017_Result_30_42_SW0_1_83 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0103,
      ADR2 => VCC,
      ADR3 => mac_control_phyaddr(30),
      O => mac_control_Mmux_n0017_Result_25_42_SW0_1_GROM
    );
  mac_control_Mmux_n0017_Result_25_42_SW0_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_25_42_SW0_1_FROM,
      O => mac_control_Mmux_n0017_Result_25_42_SW0_1
    );
  mac_control_Mmux_n0017_Result_25_42_SW0_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_25_42_SW0_1_GROM,
      O => mac_control_Mmux_n0017_Result_30_42_SW0_1
    );
  mac_control_Mmux_n0017_Result_28_42_SW0_1_84 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyaddr(28),
      ADR2 => VCC,
      ADR3 => mac_control_n0103,
      O => mac_control_Mmux_n0017_Result_28_42_SW0_1_FROM
    );
  mac_control_Mmux_n0017_Result_22_42_SW0_1_85 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyaddr(22),
      ADR2 => VCC,
      ADR3 => mac_control_n0103,
      O => mac_control_Mmux_n0017_Result_28_42_SW0_1_GROM
    );
  mac_control_Mmux_n0017_Result_28_42_SW0_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_28_42_SW0_1_FROM,
      O => mac_control_Mmux_n0017_Result_28_42_SW0_1
    );
  mac_control_Mmux_n0017_Result_28_42_SW0_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_28_42_SW0_1_GROM,
      O => mac_control_Mmux_n0017_Result_22_42_SW0_1
    );
  tx_input_fifofulll_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_fifofulll_CEMUXNOT
    );
  tx_output_crcl_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_8_FFY_RST
    );
  tx_output_crcl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(8),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_8_FFY_RST,
      O => tx_output_crcl(8)
    );
  tx_output_crc_loigc_Mxor_CO_8_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(0),
      ADR1 => tx_output_crc_loigc_n0115(0),
      ADR2 => tx_output_crc_loigc_n0122(0),
      ADR3 => tx_output_crc_loigc_Mxor_CO_7_Xo(1),
      O => tx_output_crcl_8_FROM
    );
  tx_output_n0034_8_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crc_8_Q,
      O => tx_output_n0034(8)
    );
  tx_output_crcl_8_XUSED : X_BUF
    port map (
      I => tx_output_crcl_8_FROM,
      O => tx_output_crc_8_Q
    );
  rx_input_fifo_fifo_BU384 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2402,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2421_FFY_RST,
      O => rx_input_fifo_fifo_N2422
    );
  rx_input_fifo_fifo_N2421_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2421_FFY_RST
    );
  rx_input_memio_n0059107 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => rx_input_memio_crcll(26),
      ADR1 => rx_input_memio_crcll(24),
      ADR2 => rx_input_memio_crcll(27),
      ADR3 => rx_input_memio_crcll(25),
      O => rx_input_memio_CHOICE2946_GROM
    );
  rx_input_memio_CHOICE2946_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE2946_GROM,
      O => rx_input_memio_CHOICE2946
    );
  rx_input_memio_n0059116 : X_LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      ADR0 => rx_input_memio_crcll(29),
      ADR1 => rx_input_memio_crcll(28),
      ADR2 => rx_input_memio_crcll(31),
      ADR3 => rx_input_memio_crcll(30),
      O => rx_input_memio_crcequal_FROM
    );
  rx_input_memio_n0059143 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_CHOICE2946,
      ADR1 => rx_input_memio_n0059143_2,
      ADR2 => rx_input_memio_n0059143_SW0_2,
      ADR3 => rx_input_memio_CHOICE2951,
      O => rx_input_memio_N80267
    );
  rx_input_memio_crcequal_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcequal_CEMUXNOT
    );
  rx_input_memio_crcequal_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcequal_FROM,
      O => rx_input_memio_CHOICE2951
    );
  mac_control_Mmux_n0017_Result_10_149_SW0 : X_LUT4
    generic map(
      INIT => X"0105"
    )
    port map (
      ADR0 => mac_control_CHOICE2449,
      ADR1 => mac_control_n0085,
      ADR2 => mac_control_CHOICE2432,
      ADR3 => mac_control_lmacaddr(10),
      O => mac_control_dout_10_FROM
    );
  mac_control_Mmux_n0017_Result_10_149 : X_LUT4
    generic map(
      INIT => X"0A3A"
    )
    port map (
      ADR0 => mac_control_dout(9),
      ADR1 => mac_control_addr(5),
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_N81665,
      O => mac_control_N77583
    );
  mac_control_dout_10_XUSED : X_BUF
    port map (
      I => mac_control_dout_10_FROM,
      O => mac_control_N81665
    );
  mac_control_PHY_status_phyaddrws_BYMUX : X_INV
    port map (
      I => mac_control_PHY_status_cs_FFd1,
      O => mac_control_PHY_status_phyaddrws_BYMUXNOT
    );
  mac_control_Mmux_n0017_Result_7_108_SW0 : X_LUT4
    generic map(
      INIT => X"F700"
    )
    port map (
      ADR0 => mac_control_sclkdeltall,
      ADR1 => mac_control_N52138,
      ADR2 => mac_control_bitcnt_109,
      ADR3 => mac_control_dout(6),
      O => mac_control_N82019_FROM
    );
  mac_control_Mmux_n0017_Result_11_108_SW0 : X_LUT4
    generic map(
      INIT => X"B0F0"
    )
    port map (
      ADR0 => mac_control_bitcnt_109,
      ADR1 => mac_control_sclkdeltall,
      ADR2 => mac_control_dout(10),
      ADR3 => mac_control_N52138,
      O => mac_control_N82019_GROM
    );
  mac_control_N82019_XUSED : X_BUF
    port map (
      I => mac_control_N82019_FROM,
      O => mac_control_N82019
    );
  mac_control_N82019_YUSED : X_BUF
    port map (
      I => mac_control_N82019_GROM,
      O => mac_control_N82013
    );
  rx_input_memio_crccomb_Mxor_CO_26_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(24),
      ADR1 => rx_input_memio_datal(7),
      ADR2 => rx_input_memio_crcl(28),
      ADR3 => rx_input_memio_datal(3),
      O => rx_input_memio_crccomb_Mxor_CO_26_Xo_1_FROM
    );
  rx_input_memio_crccomb_Mxor_n0001_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_datal(7),
      ADR3 => rx_input_memio_crcl(24),
      O => rx_input_memio_crccomb_Mxor_CO_26_Xo_1_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_26_Xo_1_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_26_Xo_1_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_26_Xo(1)
    );
  rx_input_memio_crccomb_Mxor_CO_26_Xo_1_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_26_Xo_1_GROM,
      O => rx_input_memio_crccomb_n0122(1)
    );
  tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2_86 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => tx_output_crcl(15),
      ADR1 => VCC,
      ADR2 => tx_output_data(1),
      ADR3 => tx_output_crcl(30),
      O => tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2_FROM
    );
  tx_output_crc_loigc_Mxor_n0000_Result1 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_crcl(30),
      ADR2 => VCC,
      ADR3 => tx_output_data(1),
      O => tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2_GROM
    );
  tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2_FROM,
      O => tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2
    );
  tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2_GROM,
      O => tx_output_crc_loigc_n0104(0)
    );
  tx_output_crc_loigc_Mxor_n0012_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_crcl(25),
      ADR3 => tx_output_data(6),
      O => tx_output_crc_loigc_n0122_0_FROM
    );
  tx_output_crc_loigc_Mxor_CO_9_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(28),
      ADR1 => tx_output_crcl(25),
      ADR2 => tx_output_data(3),
      ADR3 => tx_output_data(6),
      O => tx_output_crc_loigc_n0122_0_GROM
    );
  tx_output_crc_loigc_n0122_0_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0122_0_FROM,
      O => tx_output_crc_loigc_n0122(0)
    );
  tx_output_crc_loigc_n0122_0_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0122_0_GROM,
      O => tx_output_crc_loigc_Mxor_CO_9_Xo(0)
    );
  rx_output_fifo_nearfull_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifo_nearfull_CEMUXNOT
    );
  tx_output_crcl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_9_FFY_RST
    );
  tx_output_crcl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(9),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_9_FFY_RST,
      O => tx_output_crcl(9)
    );
  tx_output_crc_loigc_Mxor_CO_9_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0118(1),
      ADR1 => tx_output_crc_loigc_n0118(0),
      ADR2 => tx_output_crc_loigc_Mxor_CO_9_Xo(0),
      ADR3 => tx_output_crcl(1),
      O => tx_output_crcl_9_FROM
    );
  tx_output_n0034_9_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16,
      ADR2 => VCC,
      ADR3 => tx_output_crc_9_Q,
      O => tx_output_n0034(9)
    );
  tx_output_crcl_9_XUSED : X_BUF
    port map (
      I => tx_output_crcl_9_FROM,
      O => tx_output_crc_9_Q
    );
  addr4ext_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_3_FFY_RST
    );
  tx_input_MA_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_18,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_3_FFY_RST,
      O => addr4ext(2)
    );
  addr4ext_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_5_FFY_RST
    );
  tx_input_MA_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_20,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_5_FFY_RST,
      O => addr4ext(4)
    );
  addr4ext_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_7_FFY_RST
    );
  tx_input_MA_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_22,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_7_FFY_RST,
      O => addr4ext(6)
    );
  addr4ext_9_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_9_FFY_RST
    );
  tx_input_MA_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_24,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_9_FFY_RST,
      O => addr4ext(8)
    );
  d4_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_3_FFY_RST
    );
  tx_input_MD_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(2),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_3_FFY_RST,
      O => d4(2)
    );
  d4_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_5_FFY_RST
    );
  tx_input_MD_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(4),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_5_FFY_RST,
      O => d4(4)
    );
  d4_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_7_FFY_RST
    );
  tx_input_MD_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(6),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_7_FFY_RST,
      O => d4(6)
    );
  d4_9_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_9_FFY_RST
    );
  tx_input_MD_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(8),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_9_FFY_RST,
      O => d4(8)
    );
  tx_fifocheck_fbbpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_11_FFY_RST
    );
  tx_fifocheck_fbbpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_11_FFY_RST,
      O => tx_fifocheck_fbbpl(10)
    );
  tx_fifocheck_fbbpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_13_FFY_RST
    );
  tx_fifocheck_fbbpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_13_FFY_RST,
      O => tx_fifocheck_fbbpl(12)
    );
  tx_fifocheck_fbbpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_15_FFY_RST
    );
  tx_fifocheck_fbbpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_15_FFY_RST,
      O => tx_fifocheck_fbbpl(14)
    );
  rx_output_cs_FFd12_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd12_FFY_RST
    );
  rx_output_cs_FFd11_87 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd12,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd12_FFY_RST,
      O => rx_output_cs_FFd11
    );
  rx_output_cs_FFd14_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd14_FFY_RST
    );
  rx_output_cs_FFd13_88 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd14,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd14_FFY_RST,
      O => rx_output_cs_FFd13
    );
  rx_output_cs_FFd16_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd16_FFY_RST
    );
  rx_output_cs_FFd15_89 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd16,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd16_FFY_RST,
      O => rx_output_cs_FFd15
    );
  rx_input_fifo_fifo_BU270 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3939,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N7_FFX_RST,
      O => rx_input_fifo_fifo_N7
    );
  rx_input_fifo_fifo_N7_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N7_FFX_RST
    );
  rx_output_cs_Out41 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => rx_output_cs_FFd7,
      ADR1 => rx_output_cs_FFd8,
      ADR2 => VCC,
      ADR3 => rx_output_cs_FFd12,
      O => rx_output_cein
    );
  rx_output_n00331 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => rx_output_cs_FFd12,
      O => rx_output_ceinl_GROM
    );
  rx_output_ceinl_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_ceinl_CEMUXNOT
    );
  rx_output_ceinl_YUSED : X_BUF
    port map (
      I => rx_output_ceinl_GROM,
      O => rx_output_n0033
    );
  rx_output_cs_Out51 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_cs_FFd10,
      O => rx_output_fifo_reset_FROM
    );
  rx_output_n00341 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_cs_FFd10,
      ADR2 => RESET_IBUF,
      ADR3 => VCC,
      O => rx_output_fifo_reset_GROM
    );
  rx_output_fifo_reset_XUSED : X_BUF
    port map (
      I => rx_output_fifo_reset_FROM,
      O => rx_output_fifo_reset
    );
  rx_output_fifo_reset_YUSED : X_BUF
    port map (
      I => rx_output_fifo_reset_GROM,
      O => rx_output_n0034
    );
  rx_input_fifo_fifo_BU470 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2402,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2441_FFY_RST,
      O => rx_input_fifo_fifo_N2442
    );
  rx_input_fifo_fifo_N2441_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2441_FFY_RST
    );
  tx_input_cs_FFd6_In1 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_input_den,
      ADR3 => tx_input_cs_FFd7,
      O => tx_input_cs_FFd6_In
    );
  tx_input_n00211 : X_LUT4
    generic map(
      INIT => X"5040"
    )
    port map (
      ADR0 => RESET_IBUF_1,
      ADR1 => tx_input_cs_FFd6,
      ADR2 => tx_input_den,
      ADR3 => tx_input_cs_FFd7,
      O => tx_input_cs_FFd6_GROM
    );
  tx_input_cs_FFd6_YUSED : X_BUF
    port map (
      I => tx_input_cs_FFd6_GROM,
      O => tx_input_n0021
    );
  tx_input_n00231 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => tx_input_cs_FFd2,
      ADR1 => RESET_IBUF_1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_n0023_GROM
    );
  tx_input_n0023_YUSED : X_BUF
    port map (
      I => tx_input_n0023_GROM,
      O => tx_input_n0023
    );
  mac_control_n00101 : X_LUT4
    generic map(
      INIT => X"0080"
    )
    port map (
      ADR0 => mac_control_sclkdelta,
      ADR1 => mac_control_N52251,
      ADR2 => clkslen,
      ADR3 => RESET_IBUF,
      O => mac_control_n0010_FROM
    );
  mac_control_n001212 : X_LUT4
    generic map(
      INIT => X"0202"
    )
    port map (
      ADR0 => mac_control_sclkdelta,
      ADR1 => mac_control_N52251,
      ADR2 => mac_control_addr(7),
      ADR3 => VCC,
      O => mac_control_n0010_GROM
    );
  mac_control_n0010_XUSED : X_BUF
    port map (
      I => mac_control_n0010_FROM,
      O => mac_control_n0010
    );
  mac_control_n0010_YUSED : X_BUF
    port map (
      I => mac_control_n0010_GROM,
      O => mac_control_CHOICE1171
    );
  mac_control_n003557 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_129,
      ADR1 => mac_control_phyrstcnt_130,
      ADR2 => mac_control_phyrstcnt_131,
      ADR3 => mac_control_phyrstcnt_111,
      O => mac_control_CHOICE2746_FROM
    );
  mac_control_n003323 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_111,
      ADR1 => mac_control_phyrstcnt_129,
      ADR2 => mac_control_phyrstcnt_131,
      ADR3 => mac_control_phyrstcnt_130,
      O => mac_control_CHOICE2746_GROM
    );
  mac_control_CHOICE2746_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2746_FROM,
      O => mac_control_CHOICE2746
    );
  mac_control_CHOICE2746_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2746_GROM,
      O => mac_control_CHOICE2966
    );
  mac_control_n003544 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_126,
      ADR1 => mac_control_phyrstcnt_127,
      ADR2 => mac_control_phyrstcnt_125,
      ADR3 => mac_control_phyrstcnt_128,
      O => mac_control_CHOICE2739_FROM
    );
  mac_control_n003318 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_126,
      ADR1 => mac_control_phyrstcnt_128,
      ADR2 => mac_control_phyrstcnt_125,
      ADR3 => mac_control_phyrstcnt_127,
      O => mac_control_CHOICE2739_GROM
    );
  mac_control_CHOICE2739_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2739_FROM,
      O => mac_control_CHOICE2739
    );
  mac_control_CHOICE2739_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2739_GROM,
      O => mac_control_CHOICE2963
    );
  mac_control_n0035111 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_138,
      ADR1 => mac_control_phyrstcnt_137,
      ADR2 => mac_control_phyrstcnt_139,
      ADR3 => mac_control_phyrstcnt_136,
      O => mac_control_CHOICE2762_FROM
    );
  mac_control_n003351 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_136,
      ADR1 => mac_control_phyrstcnt_139,
      ADR2 => mac_control_phyrstcnt_137,
      ADR3 => mac_control_phyrstcnt_138,
      O => mac_control_CHOICE2762_GROM
    );
  mac_control_CHOICE2762_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2762_FROM,
      O => mac_control_CHOICE2762
    );
  mac_control_CHOICE2762_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2762_GROM,
      O => mac_control_CHOICE2974
    );
  mac_control_n003521 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_122,
      ADR1 => mac_control_phyrstcnt_124,
      ADR2 => mac_control_phyrstcnt_123,
      ADR3 => mac_control_phyrstcnt_121,
      O => mac_control_CHOICE2731_FROM
    );
  mac_control_n003526 : X_LUT4
    generic map(
      INIT => X"0100"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_120,
      ADR1 => mac_control_phyrstcnt_110,
      ADR2 => mac_control_phyrstcnt_119,
      ADR3 => mac_control_CHOICE2731,
      O => mac_control_CHOICE2731_GROM
    );
  mac_control_CHOICE2731_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2731_FROM,
      O => mac_control_CHOICE2731
    );
  mac_control_CHOICE2731_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2731_GROM,
      O => mac_control_CHOICE2732
    );
  mac_control_n003346 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_135,
      ADR1 => mac_control_phyrstcnt_134,
      ADR2 => mac_control_phyrstcnt_132,
      ADR3 => mac_control_phyrstcnt_133,
      O => mac_control_CHOICE2971_GROM
    );
  mac_control_CHOICE2971_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2971_GROM,
      O => mac_control_CHOICE2971
    );
  mac_control_n0035135 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_114,
      ADR1 => mac_control_phyrstcnt_140,
      ADR2 => mac_control_phyrstcnt_113,
      ADR3 => mac_control_phyrstcnt_112,
      O => mac_control_CHOICE2770_FROM
    );
  mac_control_n003363 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_140,
      ADR1 => mac_control_phyrstcnt_112,
      ADR2 => mac_control_phyrstcnt_113,
      ADR3 => mac_control_phyrstcnt_114,
      O => mac_control_CHOICE2770_GROM
    );
  mac_control_CHOICE2770_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2770_FROM,
      O => mac_control_CHOICE2770
    );
  mac_control_CHOICE2770_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2770_GROM,
      O => mac_control_CHOICE2978
    );
  mac_control_n0035148 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_116,
      ADR1 => mac_control_phyrstcnt_117,
      ADR2 => mac_control_phyrstcnt_118,
      ADR3 => mac_control_phyrstcnt_115,
      O => mac_control_CHOICE2777_FROM
    );
  mac_control_n003368 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_116,
      ADR1 => mac_control_phyrstcnt_115,
      ADR2 => mac_control_phyrstcnt_118,
      ADR3 => mac_control_phyrstcnt_117,
      O => mac_control_CHOICE2777_GROM
    );
  mac_control_CHOICE2777_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2777_FROM,
      O => mac_control_CHOICE2777
    );
  mac_control_CHOICE2777_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2777_GROM,
      O => mac_control_CHOICE2981
    );
  mac_control_n007025 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_145,
      ADR1 => mac_control_ledtx_cnt_142,
      ADR2 => mac_control_ledtx_cnt_143,
      ADR3 => mac_control_ledtx_cnt_144,
      O => mac_control_CHOICE1609_GROM
    );
  mac_control_CHOICE1609_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1609_GROM,
      O => mac_control_CHOICE1609
    );
  mac_control_n007050 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_151,
      ADR1 => mac_control_N81797,
      ADR2 => mac_control_ledtx_cnt_152,
      ADR3 => mac_control_ledtx_cnt_150,
      O => mac_control_N73201_FROM
    );
  mac_control_n00381 : X_LUT4
    generic map(
      INIT => X"2030"
    )
    port map (
      ADR0 => mac_control_ledtx_rst,
      ADR1 => RESET_IBUF,
      ADR2 => clkslen,
      ADR3 => mac_control_N73201,
      O => mac_control_N73201_GROM
    );
  mac_control_N73201_XUSED : X_BUF
    port map (
      I => mac_control_N73201_FROM,
      O => mac_control_N73201
    );
  mac_control_N73201_YUSED : X_BUF
    port map (
      I => mac_control_N73201_GROM,
      O => mac_control_n0038
    );
  rx_input_fifo_fifo_BU386 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2401,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2421_FFX_RST,
      O => rx_input_fifo_fifo_N2421
    );
  rx_input_fifo_fifo_N2421_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2421_FFX_RST
    );
  tx_output_crc_loigc_Mxor_CO_0_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(1),
      ADR1 => tx_output_crcl(30),
      ADR2 => tx_output_crcl(24),
      ADR3 => tx_output_data(7),
      O => tx_output_crcl_0_FROM
    );
  tx_output_n0034_0_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16,
      ADR2 => VCC,
      ADR3 => tx_output_crc_0_Q,
      O => tx_output_n0034(0)
    );
  tx_output_crcl_0_XUSED : X_BUF
    port map (
      I => tx_output_crcl_0_FROM,
      O => tx_output_crc_0_Q
    );
  mac_control_n007125 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_157,
      ADR1 => mac_control_ledrx_cnt_154,
      ADR2 => mac_control_ledrx_cnt_156,
      ADR3 => mac_control_ledrx_cnt_155,
      O => mac_control_CHOICE1586_GROM
    );
  mac_control_CHOICE1586_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1586_GROM,
      O => mac_control_CHOICE1586
    );
  mac_control_n007038 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_146,
      ADR1 => mac_control_ledtx_cnt_148,
      ADR2 => mac_control_ledtx_cnt_147,
      ADR3 => mac_control_ledtx_cnt_149,
      O => mac_control_CHOICE1616_GROM
    );
  mac_control_CHOICE1616_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1616_GROM,
      O => mac_control_CHOICE1616
    );
  mac_control_n003598 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_135,
      ADR1 => mac_control_phyrstcnt_133,
      ADR2 => mac_control_phyrstcnt_132,
      ADR3 => mac_control_phyrstcnt_134,
      O => mac_control_CHOICE2755_FROM
    );
  mac_control_n0035194_SW0_2_90 : X_LUT4
    generic map(
      INIT => X"A000"
    )
    port map (
      ADR0 => mac_control_CHOICE2746,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE2762,
      ADR3 => mac_control_CHOICE2755,
      O => mac_control_CHOICE2755_GROM
    );
  mac_control_CHOICE2755_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2755_FROM,
      O => mac_control_CHOICE2755
    );
  mac_control_CHOICE2755_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2755_GROM,
      O => mac_control_n0035194_SW0_2
    );
  mac_control_n007150 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_162,
      ADR1 => mac_control_ledrx_cnt_163,
      ADR2 => mac_control_N81777,
      ADR3 => mac_control_ledrx_cnt_164,
      O => mac_control_N73084_FROM
    );
  mac_control_n00401 : X_LUT4
    generic map(
      INIT => X"00D0"
    )
    port map (
      ADR0 => mac_control_N73084,
      ADR1 => mac_control_ledrx_rst,
      ADR2 => clkslen,
      ADR3 => RESET_IBUF,
      O => mac_control_N73084_GROM
    );
  mac_control_N73084_XUSED : X_BUF
    port map (
      I => mac_control_N73084_FROM,
      O => mac_control_N73084
    );
  mac_control_N73084_YUSED : X_BUF
    port map (
      I => mac_control_N73084_GROM,
      O => mac_control_n0040
    );
  mac_control_n007138 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_159,
      ADR1 => mac_control_ledrx_cnt_160,
      ADR2 => mac_control_ledrx_cnt_161,
      ADR3 => mac_control_ledrx_cnt_158,
      O => mac_control_CHOICE1593_GROM
    );
  mac_control_CHOICE1593_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1593_GROM,
      O => mac_control_CHOICE1593
    );
  slowclock_rxfl_LOGIC_ZERO_91 : X_ZERO
    port map (
      O => slowclock_rxfl_LOGIC_ZERO
    );
  slowclock_rxfl_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => slowclock_rxfl_GROM
    );
  slowclock_txfl_LOGIC_ZERO_92 : X_ZERO
    port map (
      O => slowclock_txfl_LOGIC_ZERO
    );
  slowclock_txfl_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => slowclock_txfl_GROM
    );
  tx_input_dh_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_3_FFY_RST
    );
  tx_input_dh_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(2),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_3_FFY_RST,
      O => tx_input_dh(2)
    );
  tx_input_dh_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_5_FFY_RST
    );
  tx_input_dh_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(4),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_5_FFY_RST,
      O => tx_input_dh(4)
    );
  rx_input_memio_crccomb_Mxor_n0003_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_datal(5),
      ADR3 => rx_input_memio_crcl(26),
      O => rx_input_memio_crccomb_n0118_1_FROM
    );
  rx_input_memio_crccomb_Mxor_CO_14_Xo_3_1_2_93 : X_LUT4
    generic map(
      INIT => X"C33C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcl(28),
      ADR2 => rx_input_memio_datal(3),
      ADR3 => rx_input_memio_crccomb_n0118(1),
      O => rx_input_memio_crccomb_n0118_1_GROM
    );
  rx_input_memio_crccomb_n0118_1_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_n0118_1_FROM,
      O => rx_input_memio_crccomb_n0118(1)
    );
  rx_input_memio_crccomb_n0118_1_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_n0118_1_GROM,
      O => rx_input_memio_crccomb_Mxor_CO_14_Xo_3_1_2
    );
  rx_input_fifo_fifo_BU450 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N6,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2472_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2471
    );
  rx_input_fifo_fifo_N2472_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2472_FFY_SET
    );
  rx_input_memio_crccomb_Mxor_n0011_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_datal(0),
      ADR3 => rx_input_memio_crcl(31),
      O => rx_input_memio_crccomb_n0124_0_FROM
    );
  rx_input_memio_crccomb_Mxor_CO_5_Xo_1_1_2_94 : X_LUT4
    generic map(
      INIT => X"C33C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crccomb_Mxor_n0007_Xo(0),
      ADR2 => rx_input_memio_crccomb_n0124(1),
      ADR3 => rx_input_memio_crccomb_n0124(0),
      O => rx_input_memio_crccomb_n0124_0_GROM
    );
  rx_input_memio_crccomb_n0124_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_n0124_0_FROM,
      O => rx_input_memio_crccomb_n0124(0)
    );
  rx_input_memio_crccomb_n0124_0_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_n0124_0_GROM,
      O => rx_input_memio_crccomb_Mxor_CO_5_Xo_1_1_2
    );
  tx_input_dh_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_9_FFY_RST
    );
  tx_input_dh_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(8),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_9_FFY_RST,
      O => tx_input_dh(8)
    );
  tx_input_dl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_1_FFY_RST
    );
  tx_input_dl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(0),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_1_FFY_RST,
      O => tx_input_dl(0)
    );
  tx_input_dl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_3_FFY_RST
    );
  tx_input_dl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(2),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_3_FFY_RST,
      O => tx_input_dl(2)
    );
  tx_input_dl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_5_FFY_RST
    );
  tx_input_dl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(4),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_5_FFY_RST,
      O => tx_input_dl(4)
    );
  tx_input_dl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_7_FFY_RST
    );
  tx_input_dl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(6),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_7_FFY_RST,
      O => tx_input_dl(6)
    );
  rx_input_fifo_fifo_BU414 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2422,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2432_FFX_RST,
      O => rx_input_fifo_fifo_N2432
    );
  rx_input_fifo_fifo_N2432_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2432_FFX_RST
    );
  tx_input_dl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_9_FFY_RST
    );
  tx_input_dl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(8),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_9_FFY_RST,
      O => tx_input_dl(8)
    );
  txbp_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_9_FFX_RST
    );
  tx_input_bp_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_25,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_9_FFX_RST,
      O => txbp(9)
    );
  MDC_OBUF_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MDC_OBUF_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_mdcint : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_37,
      CE => mac_control_PHY_status_MII_Interface_N37245,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MDC_OBUF_FFY_RST,
      O => MDC_OBUF
    );
  mac_control_Mmux_n0017_Result_10_107 : X_LUT4
    generic map(
      INIT => X"9910"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_N82121,
      ADR3 => mac_control_N52125,
      O => mac_control_CHOICE2448_FROM
    );
  mac_control_Mmux_n0017_Result_10_113 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_CHOICE2442,
      ADR1 => mac_control_N52244,
      ADR2 => mac_control_CHOICE2436,
      ADR3 => mac_control_CHOICE2448,
      O => mac_control_CHOICE2448_GROM
    );
  mac_control_CHOICE2448_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2448_FROM,
      O => mac_control_CHOICE2448
    );
  mac_control_CHOICE2448_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2448_GROM,
      O => mac_control_CHOICE2449
    );
  mac_control_lmacaddr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_1_FFX_RST
    );
  mac_control_lmacaddr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_1_FFX_RST,
      O => mac_control_lmacaddr(1)
    );
  mac_control_lmacaddr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_1_FFY_RST
    );
  mac_control_lmacaddr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_1_FFY_RST,
      O => mac_control_lmacaddr(0)
    );
  mac_control_lmacaddr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_3_FFX_RST
    );
  mac_control_lmacaddr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_3_FFX_RST,
      O => mac_control_lmacaddr(3)
    );
  mac_control_lmacaddr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_3_FFY_RST
    );
  mac_control_lmacaddr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_3_FFY_RST,
      O => mac_control_lmacaddr(2)
    );
  rx_input_fifo_fifo_BU472 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2401,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2441_FFX_RST,
      O => rx_input_fifo_fifo_N2441
    );
  rx_input_fifo_fifo_N2441_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2441_FFX_RST
    );
  mac_control_lmacaddr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_5_FFX_RST
    );
  mac_control_lmacaddr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_5_FFX_RST,
      O => mac_control_lmacaddr(5)
    );
  mac_control_lmacaddr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_5_FFY_RST
    );
  mac_control_lmacaddr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_5_FFY_RST,
      O => mac_control_lmacaddr(4)
    );
  mac_control_lmacaddr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_7_FFX_RST
    );
  mac_control_lmacaddr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_7_FFX_RST,
      O => mac_control_lmacaddr(7)
    );
  mac_control_lmacaddr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_7_FFY_RST
    );
  mac_control_lmacaddr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_7_FFY_RST,
      O => mac_control_lmacaddr(6)
    );
  mac_control_lmacaddr_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_9_FFX_RST
    );
  mac_control_lmacaddr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_9_FFX_RST,
      O => mac_control_lmacaddr(9)
    );
  mac_control_lmacaddr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_9_FFY_RST
    );
  mac_control_lmacaddr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_9_FFY_RST,
      O => mac_control_lmacaddr(8)
    );
  rxbp_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_1_FFX_RST
    );
  rx_input_memio_BPOUT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_1_68,
      CE => rxbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_1_FFX_RST,
      O => rxbp(1)
    );
  rxbp_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_1_FFY_RST
    );
  rx_input_memio_BPOUT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_0_69,
      CE => rxbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_1_FFY_RST,
      O => rxbp(0)
    );
  rxbp_1_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxbp_1_CEMUXNOT
    );
  rxbp_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_3_FFY_RST
    );
  rx_input_memio_BPOUT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_2_67,
      CE => rxbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_3_FFY_RST,
      O => rxbp(2)
    );
  rxbp_3_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxbp_3_CEMUXNOT
    );
  rxbp_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_5_FFY_RST
    );
  rx_input_memio_BPOUT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_4_65,
      CE => rxbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_5_FFY_RST,
      O => rxbp(4)
    );
  rxbp_5_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxbp_5_CEMUXNOT
    );
  rxbp_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_7_FFY_RST
    );
  rx_input_memio_BPOUT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_6_63,
      CE => rxbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_7_FFY_RST,
      O => rxbp(6)
    );
  rxbp_7_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxbp_7_CEMUXNOT
    );
  rxbp_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_9_FFY_RST
    );
  rx_input_memio_BPOUT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_8_61,
      CE => rxbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_9_FFY_RST,
      O => rxbp(8)
    );
  rxbp_9_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxbp_9_CEMUXNOT
    );
  rxfbbp_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_1_FFY_RST
    );
  rx_output_FBBP_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(0),
      CE => rxfbbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_1_FFY_RST,
      O => rxfbbp(0)
    );
  rxfbbp_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_1_CEMUXNOT
    );
  rxfbbp_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_3_FFY_RST
    );
  rx_output_FBBP_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(2),
      CE => rxfbbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_3_FFY_RST,
      O => rxfbbp(2)
    );
  rxfbbp_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_3_CEMUXNOT
    );
  rxfbbp_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_5_FFY_RST
    );
  rx_output_FBBP_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(4),
      CE => rxfbbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_5_FFY_RST,
      O => rxfbbp(4)
    );
  rxfbbp_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_5_CEMUXNOT
    );
  rxfbbp_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_7_CEMUXNOT
    );
  rxfbbp_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_9_FFY_RST
    );
  rx_output_FBBP_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(8),
      CE => rxfbbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_9_FFY_RST,
      O => rxfbbp(8)
    );
  rxfbbp_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_9_CEMUXNOT
    );
  mac_control_Mmux_n0017_Result_14_107 : X_LUT4
    generic map(
      INIT => X"8584"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => mac_control_N52125,
      ADR2 => mac_control_addr(1),
      ADR3 => mac_control_N82117,
      O => mac_control_CHOICE2486_FROM
    );
  mac_control_Mmux_n0017_Result_14_113 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_CHOICE2474,
      ADR1 => mac_control_N52244,
      ADR2 => mac_control_CHOICE2480,
      ADR3 => mac_control_CHOICE2486,
      O => mac_control_CHOICE2486_GROM
    );
  mac_control_CHOICE2486_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2486_FROM,
      O => mac_control_CHOICE2486
    );
  mac_control_CHOICE2486_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2486_GROM,
      O => mac_control_CHOICE2487
    );
  rx_input_memio_addrchk_macaddrl_1_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_1_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_3_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(2),
      CE => rx_input_memio_addrchk_macaddrl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_3_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(2)
    );
  rx_input_memio_addrchk_macaddrl_3_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_3_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_5_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(4),
      CE => rx_input_memio_addrchk_macaddrl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_5_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(4)
    );
  rx_input_memio_addrchk_macaddrl_5_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_5_CEMUXNOT
    );
  rx_input_fifo_fifo_BU448 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N7,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2472_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2472
    );
  rx_input_fifo_fifo_N2472_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2472_FFX_SET
    );
  rx_input_memio_addrchk_macaddrl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_7_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(6),
      CE => rx_input_memio_addrchk_macaddrl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_7_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(6)
    );
  rx_input_memio_addrchk_macaddrl_7_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_7_CEMUXNOT
    );
  rx_input_fifo_fifo_BU564 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N5345,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2451_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2452
    );
  rx_input_fifo_fifo_N2451_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2451_FFY_SET
    );
  rx_input_memio_addrchk_macaddrl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_9_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(8),
      CE => rx_input_memio_addrchk_macaddrl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_9_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(8)
    );
  rx_input_memio_addrchk_macaddrl_9_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_9_CEMUXNOT
    );
  mac_control_Mmux_n0017_Result_8_107_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phyaddr(8),
      ADR1 => mac_control_N52132,
      ADR2 => mac_control_rxfifowerr_cnt(8),
      ADR3 => mac_control_N52111,
      O => mac_control_N82129_FROM
    );
  mac_control_Mmux_n0017_Result_14_107_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phyaddr(14),
      ADR1 => mac_control_N52132,
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_rxfifowerr_cnt(14),
      O => mac_control_N82129_GROM
    );
  mac_control_N82129_XUSED : X_BUF
    port map (
      I => mac_control_N82129_FROM,
      O => mac_control_N82129
    );
  mac_control_N82129_YUSED : X_BUF
    port map (
      I => mac_control_N82129_GROM,
      O => mac_control_N82117
    );
  rx_output_n0046_2_SW0 : X_LUT4
    generic map(
      INIT => X"5533"
    )
    port map (
      ADR0 => rx_output_n0070(2),
      ADR1 => rx_output_len(2),
      ADR2 => VCC,
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_2_FROM
    );
  rx_output_n0046_2_Q : X_LUT4
    generic map(
      INIT => X"A0AF"
    )
    port map (
      ADR0 => rx_output_n0060(2),
      ADR1 => VCC,
      ADR2 => rx_output_len(0),
      ADR3 => rx_output_N69852,
      O => rx_output_n0046(2)
    );
  rx_output_lenr_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_2_CEMUXNOT
    );
  rx_output_lenr_2_XUSED : X_BUF
    port map (
      I => rx_output_lenr_2_FROM,
      O => rx_output_N69852
    );
  rx_input_memio_crccomb_Mxor_n0004_Result1 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_input_memio_crcl(27),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_datal(4),
      O => rx_input_memio_crcl_25_FROM
    );
  rx_input_memio_n0048_25_1 : X_LUT4
    generic map(
      INIT => X"F3FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crccomb_Mxor_CO_25_Xo_1_1_2,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crccomb_n0124(1),
      O => rx_input_memio_n0048(25)
    );
  rx_input_memio_crcl_25_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_25_FROM,
      O => rx_input_memio_crccomb_n0124(1)
    );
  rx_input_memio_crccomb_Mxor_CO_9_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(28),
      ADR1 => rx_input_memio_crcl(25),
      ADR2 => rx_input_memio_datal(3),
      ADR3 => rx_input_memio_datal(6),
      O => rx_input_memio_crccomb_Mxor_CO_9_Xo_0_FROM
    );
  rx_input_memio_crccomb_Mxor_n0012_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_datal(6),
      ADR3 => rx_input_memio_crcl(25),
      O => rx_input_memio_crccomb_Mxor_CO_9_Xo_0_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_9_Xo_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_9_Xo_0_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_9_Xo(0)
    );
  rx_input_memio_crccomb_Mxor_CO_9_Xo_0_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_9_Xo_0_GROM,
      O => rx_input_memio_crccomb_n0122(0)
    );
  tx_output_crc_loigc_Mxor_n0003_Result1 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_crcl(26),
      ADR2 => VCC,
      ADR3 => tx_output_data(5),
      O => tx_output_crc_loigc_n0118_1_FROM
    );
  tx_output_crc_loigc_Mxor_CO_4_Xo_1_1_2_95 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => tx_output_crcl(27),
      ADR1 => VCC,
      ADR2 => tx_output_data(4),
      ADR3 => tx_output_crc_loigc_n0118(1),
      O => tx_output_crc_loigc_n0118_1_GROM
    );
  tx_output_crc_loigc_n0118_1_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0118_1_FROM,
      O => tx_output_crc_loigc_n0118(1)
    );
  tx_output_crc_loigc_n0118_1_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0118_1_GROM,
      O => tx_output_crc_loigc_Mxor_CO_4_Xo_1_1_2
    );
  tx_output_crc_loigc_Mxor_n0011_Result1 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_crcl(31),
      ADR2 => tx_output_data(0),
      ADR3 => VCC,
      O => tx_output_crc_loigc_n0124_0_FROM
    );
  tx_output_crc_loigc_Mxor_CO_5_Xo_1_1_2_96 : X_LUT4
    generic map(
      INIT => X"C33C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_crc_loigc_Mxor_n0007_Xo(0),
      ADR2 => tx_output_crc_loigc_n0124(0),
      ADR3 => tx_output_crc_loigc_n0124(1),
      O => tx_output_crc_loigc_n0124_0_GROM
    );
  tx_output_crc_loigc_n0124_0_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0124_0_FROM,
      O => tx_output_crc_loigc_n0124(0)
    );
  tx_output_crc_loigc_n0124_0_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0124_0_GROM,
      O => tx_output_crc_loigc_Mxor_CO_5_Xo_1_1_2
    );
  rx_output_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd6_FFY_RST
    );
  rx_output_cs_FFd6_97 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd6_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd6_FFY_RST,
      O => rx_output_cs_FFd6
    );
  rx_output_cs_FFd6_In_SW0 : X_LUT4
    generic map(
      INIT => X"CC8C"
    )
    port map (
      ADR0 => rx_output_fifo_nearfull,
      ADR1 => rx_output_cs_FFd6,
      ADR2 => memcontroller_clknum(1),
      ADR3 => memcontroller_clknum(0),
      O => rx_output_cs_FFd6_FROM
    );
  rx_output_cs_FFd6_In_98 : X_LUT4
    generic map(
      INIT => X"CC80"
    )
    port map (
      ADR0 => rx_output_cs_FFd7,
      ADR1 => rx_output_nf,
      ADR2 => rx_output_fifo_full,
      ADR3 => rx_output_N70424,
      O => rx_output_cs_FFd6_In
    );
  rx_output_cs_FFd6_XUSED : X_BUF
    port map (
      I => rx_output_cs_FFd6_FROM,
      O => rx_output_N70424
    );
  rx_output_n0046_3_SW0 : X_LUT4
    generic map(
      INIT => X"05F5"
    )
    port map (
      ADR0 => rx_output_len(3),
      ADR1 => VCC,
      ADR2 => rx_output_len(1),
      ADR3 => rx_output_n0070(3),
      O => rx_output_lenr_3_FROM
    );
  rx_output_n0046_3_Q : X_LUT4
    generic map(
      INIT => X"88BB"
    )
    port map (
      ADR0 => rx_output_n0060(3),
      ADR1 => rx_output_len(0),
      ADR2 => VCC,
      ADR3 => rx_output_N69800,
      O => rx_output_n0046(3)
    );
  rx_output_lenr_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_3_CEMUXNOT
    );
  rx_output_lenr_3_XUSED : X_BUF
    port map (
      I => rx_output_lenr_3_FROM,
      O => rx_output_N69800
    );
  rx_output_n0046_4_SW0 : X_LUT4
    generic map(
      INIT => X"330F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_n0070(4),
      ADR2 => rx_output_len(4),
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_4_FROM
    );
  rx_output_n0046_4_Q : X_LUT4
    generic map(
      INIT => X"A0F5"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => VCC,
      ADR2 => rx_output_n0060(4),
      ADR3 => rx_output_N69904,
      O => rx_output_n0046(4)
    );
  rx_output_lenr_4_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_4_CEMUXNOT
    );
  rx_output_lenr_4_XUSED : X_BUF
    port map (
      I => rx_output_lenr_4_FROM,
      O => rx_output_N69904
    );
  rx_output_cs_FFd10_In5 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_output_cs_FFd8,
      ADR1 => rx_output_cs_FFd4,
      ADR2 => rx_output_cs_FFd5,
      ADR3 => rx_output_cs_FFd6,
      O => rx_output_CHOICE1557_FROM
    );
  rx_output_cs_Out64 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_output_cs_FFd2,
      ADR1 => rx_output_cs_FFd1,
      ADR2 => rx_output_cs_FFd6,
      ADR3 => rx_output_cs_FFd3,
      O => rx_output_CHOICE1557_GROM
    );
  rx_output_CHOICE1557_XUSED : X_BUF
    port map (
      I => rx_output_CHOICE1557_FROM,
      O => rx_output_CHOICE1557
    );
  rx_output_CHOICE1557_YUSED : X_BUF
    port map (
      I => rx_output_CHOICE1557_GROM,
      O => rx_output_CHOICE1525
    );
  rx_output_denl_LOGIC_ZERO_99 : X_ZERO
    port map (
      O => rx_output_denl_LOGIC_ZERO
    );
  rx_output_cs_Out68 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => rx_output_cs_FFd5,
      ADR1 => rx_output_cs_FFd8,
      ADR2 => VCC,
      ADR3 => rx_output_cs_FFd7,
      O => rx_output_denl_FROM
    );
  rx_output_cs_Out610 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => rx_output_cs_FFd9,
      ADR1 => rx_output_cs_FFd4,
      ADR2 => VCC,
      ADR3 => rx_output_CHOICE1528,
      O => rx_output_CHOICE1529
    );
  rx_output_denl_XUSED : X_BUF
    port map (
      I => rx_output_denl_FROM,
      O => rx_output_CHOICE1528
    );
  rx_output_n0046_5_SW0 : X_LUT4
    generic map(
      INIT => X"4477"
    )
    port map (
      ADR0 => rx_output_n0070(5),
      ADR1 => rx_output_len(1),
      ADR2 => VCC,
      ADR3 => rx_output_len(5),
      O => rx_output_lenr_5_FROM
    );
  rx_output_n0046_5_Q : X_LUT4
    generic map(
      INIT => X"A0AF"
    )
    port map (
      ADR0 => rx_output_n0060(5),
      ADR1 => VCC,
      ADR2 => rx_output_len(0),
      ADR3 => rx_output_N69956,
      O => rx_output_n0046(5)
    );
  rx_output_lenr_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_5_CEMUXNOT
    );
  rx_output_lenr_5_XUSED : X_BUF
    port map (
      I => rx_output_lenr_5_FROM,
      O => rx_output_N69956
    );
  rx_output_lenr_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_6_FFY_RST
    );
  rx_output_lenr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(6),
      CE => rx_output_lenr_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_6_FFY_RST,
      O => rx_output_lenr(6)
    );
  rx_output_n0046_6_SW0 : X_LUT4
    generic map(
      INIT => X"03CF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(1),
      ADR2 => rx_output_len(6),
      ADR3 => rx_output_n0070(6),
      O => rx_output_lenr_6_FROM
    );
  rx_output_n0046_6_Q : X_LUT4
    generic map(
      INIT => X"A0F5"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => VCC,
      ADR2 => rx_output_n0060(6),
      ADR3 => rx_output_N70008,
      O => rx_output_n0046(6)
    );
  rx_output_lenr_6_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_6_CEMUXNOT
    );
  rx_output_lenr_6_XUSED : X_BUF
    port map (
      I => rx_output_lenr_6_FROM,
      O => rx_output_N70008
    );
  mac_control_Mmux_n0017_Result_14_149_SW0 : X_LUT4
    generic map(
      INIT => X"0105"
    )
    port map (
      ADR0 => mac_control_CHOICE2487,
      ADR1 => mac_control_lmacaddr(14),
      ADR2 => mac_control_CHOICE2470,
      ADR3 => mac_control_n0085,
      O => mac_control_dout_14_FROM
    );
  mac_control_Mmux_n0017_Result_14_149 : X_LUT4
    generic map(
      INIT => X"0C5C"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_dout(13),
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_N81637,
      O => mac_control_N77791
    );
  mac_control_dout_14_XUSED : X_BUF
    port map (
      I => mac_control_dout_14_FROM,
      O => mac_control_N81637
    );
  mac_control_PHY_status_MII_Interface_sout27 : X_LUT4
    generic map(
      INIT => X"0E04"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_din(15),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR3 => mac_control_PHY_status_din(7),
      O => mac_control_PHY_status_MII_Interface_CHOICE2503_FROM
    );
  mac_control_PHY_status_MII_Interface_sout12 : X_LUT4
    generic map(
      INIT => X"A280"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR2 => mac_control_PHY_status_din(3),
      ADR3 => mac_control_PHY_status_din(11),
      O => mac_control_PHY_status_MII_Interface_CHOICE2503_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE2503_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2503_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2503
    );
  mac_control_PHY_status_MII_Interface_CHOICE2503_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2503_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2497
    );
  tx_output_crc_loigc_Mxor_CO_1_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_0_Q,
      ADR1 => tx_output_crcl(31),
      ADR2 => tx_output_data(0),
      ADR3 => tx_output_crc_loigc_n0122(0),
      O => tx_output_crcl_1_FROM
    );
  tx_output_n0034_1_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_1_Q,
      O => tx_output_n0034(1)
    );
  tx_output_crcl_1_XUSED : X_BUF
    port map (
      I => tx_output_crcl_1_FROM,
      O => tx_output_crc_1_Q
    );
  mac_control_PHY_status_MII_Interface_sout63 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_CHOICE2511_FROM
    );
  mac_control_PHY_status_MII_Interface_sout68 : X_LUT4
    generic map(
      INIT => X"CA00"
    )
    port map (
      ADR0 => mac_control_PHY_status_din(10),
      ADR1 => mac_control_PHY_status_din(2),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE2511,
      O => mac_control_PHY_status_MII_Interface_CHOICE2511_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE2511_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2511_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2511
    );
  mac_control_PHY_status_MII_Interface_CHOICE2511_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2511_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2512
    );
  rx_output_n0046_7_SW0 : X_LUT4
    generic map(
      INIT => X"550F"
    )
    port map (
      ADR0 => rx_output_n0070(7),
      ADR1 => VCC,
      ADR2 => rx_output_len(7),
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_7_FROM
    );
  rx_output_n0046_7_Q : X_LUT4
    generic map(
      INIT => X"A0AF"
    )
    port map (
      ADR0 => rx_output_n0060(7),
      ADR1 => VCC,
      ADR2 => rx_output_len(0),
      ADR3 => rx_output_N70112,
      O => rx_output_n0046(7)
    );
  rx_output_lenr_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_7_CEMUXNOT
    );
  rx_output_lenr_7_XUSED : X_BUF
    port map (
      I => rx_output_lenr_7_FROM,
      O => rx_output_N70112
    );
  mac_control_PHY_status_MII_Interface_sout73 : X_LUT4
    generic map(
      INIT => X"CCFE"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_CHOICE2497,
      ADR1 => mac_control_PHY_status_MII_Interface_CHOICE2512,
      ADR2 => mac_control_PHY_status_MII_Interface_CHOICE2503,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(0),
      O => mac_control_PHY_status_MII_Interface_CHOICE2513_FROM
    );
  mac_control_PHY_status_MII_Interface_sout498_2_100 : X_LUT4
    generic map(
      INIT => X"AFFF"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(1),
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE2513,
      O => mac_control_PHY_status_MII_Interface_CHOICE2513_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE2513_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2513_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2513
    );
  mac_control_PHY_status_MII_Interface_CHOICE2513_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2513_GROM,
      O => mac_control_PHY_status_MII_Interface_sout498_2
    );
  mac_control_Mmux_n0017_Result_3_108_1_101 : X_LUT4
    generic map(
      INIT => X"F0FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_dout(2),
      O => mac_control_Mmux_n0017_Result_3_108_1_FROM
    );
  mac_control_Mmux_n0017_Result_3_96_1_102 : X_LUT4
    generic map(
      INIT => X"F5F5"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => VCC,
      ADR2 => mac_control_addr(5),
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_3_108_1_GROM
    );
  mac_control_Mmux_n0017_Result_3_108_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_3_108_1_FROM,
      O => mac_control_Mmux_n0017_Result_3_108_1
    );
  mac_control_Mmux_n0017_Result_3_108_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_3_108_1_GROM,
      O => mac_control_Mmux_n0017_Result_3_96_1
    );
  mac_control_Mmux_n0017_Result_31_103_SW1 : X_LUT4
    generic map(
      INIT => X"0007"
    )
    port map (
      ADR0 => mac_control_N52132,
      ADR1 => mac_control_CHOICE1817,
      ADR2 => mac_control_CHOICE1821,
      ADR3 => mac_control_CHOICE1814,
      O => mac_control_dout_31_FROM
    );
  mac_control_Mmux_n0017_Result_31_103 : X_LUT4
    generic map(
      INIT => X"0A3A"
    )
    port map (
      ADR0 => mac_control_dout(30),
      ADR1 => mac_control_addr(5),
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_N82074,
      O => mac_control_N74276
    );
  mac_control_dout_31_XUSED : X_BUF
    port map (
      I => mac_control_dout_31_FROM,
      O => mac_control_N82074
    );
  mac_control_Mmux_n0017_Result_23_103_SW1 : X_LUT4
    generic map(
      INIT => X"0015"
    )
    port map (
      ADR0 => mac_control_CHOICE1870,
      ADR1 => mac_control_CHOICE1873,
      ADR2 => mac_control_N52132,
      ADR3 => mac_control_CHOICE1877,
      O => mac_control_dout_23_FROM
    );
  mac_control_Mmux_n0017_Result_23_103 : X_LUT4
    generic map(
      INIT => X"3074"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_n0060,
      ADR2 => mac_control_dout(22),
      ADR3 => mac_control_N82082,
      O => mac_control_N74572
    );
  mac_control_dout_23_XUSED : X_BUF
    port map (
      I => mac_control_dout_23_FROM,
      O => mac_control_N82082
    );
  rx_input_fifo_fifo_BU566 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N5346,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2451_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2451
    );
  rx_input_fifo_fifo_N2451_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2451_FFX_SET
    );
  rx_output_n0046_8_SW0 : X_LUT4
    generic map(
      INIT => X"05F5"
    )
    port map (
      ADR0 => rx_output_len(8),
      ADR1 => VCC,
      ADR2 => rx_output_len(1),
      ADR3 => rx_output_n0070(8),
      O => rx_output_lenr_8_FROM
    );
  rx_output_n0046_8_Q : X_LUT4
    generic map(
      INIT => X"A0F5"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => VCC,
      ADR2 => rx_output_n0060(8),
      ADR3 => rx_output_N70060,
      O => rx_output_n0046(8)
    );
  rx_output_lenr_8_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_8_CEMUXNOT
    );
  rx_output_lenr_8_XUSED : X_BUF
    port map (
      I => rx_output_lenr_8_FROM,
      O => rx_output_N70060
    );
  tx_input_cs_Out51 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => tx_input_cs_FFd4,
      ADR1 => VCC,
      ADR2 => tx_input_cs_FFd6,
      ADR3 => tx_input_cs_FFd11,
      O => tx_input_mrw_GROM
    );
  tx_input_mrw_YUSED : X_BUF
    port map (
      I => tx_input_mrw_GROM,
      O => tx_input_mrw
    );
  rx_output_n0046_9_SW0 : X_LUT4
    generic map(
      INIT => X"0F55"
    )
    port map (
      ADR0 => rx_output_len(9),
      ADR1 => VCC,
      ADR2 => rx_output_n0070(9),
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_9_FROM
    );
  rx_output_n0046_9_Q : X_LUT4
    generic map(
      INIT => X"A0F5"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => VCC,
      ADR2 => rx_output_n0060(9),
      ADR3 => rx_output_N70164,
      O => rx_output_n0046(9)
    );
  rx_output_lenr_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_9_CEMUXNOT
    );
  rx_output_lenr_9_XUSED : X_BUF
    port map (
      I => rx_output_lenr_9_FROM,
      O => rx_output_N70164
    );
  rx_input_memio_addrchk_n00504 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(41),
      ADR1 => rx_input_memio_addrchk_datal(43),
      ADR2 => rx_input_memio_addrchk_datal(40),
      ADR3 => rx_input_memio_addrchk_datal(42),
      O => rx_input_memio_addrchk_CHOICE1403_FROM
    );
  rx_input_memio_addrchk_n004911 : X_LUT4
    generic map(
      INIT => X"0010"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(42),
      ADR1 => rx_input_memio_addrchk_datal(43),
      ADR2 => rx_input_memio_addrchk_datal(40),
      ADR3 => rx_input_memio_addrchk_datal(41),
      O => rx_input_memio_addrchk_CHOICE1403_GROM
    );
  rx_input_memio_addrchk_CHOICE1403_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1403_FROM,
      O => rx_input_memio_addrchk_CHOICE1403
    );
  rx_input_memio_addrchk_CHOICE1403_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1403_GROM,
      O => rx_input_memio_addrchk_CHOICE1392
    );
  rx_input_memio_addrchk_n004924 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(46),
      ADR1 => rx_input_memio_addrchk_datal(47),
      ADR2 => rx_input_memio_addrchk_datal(44),
      ADR3 => rx_input_memio_addrchk_datal(45),
      O => rx_input_memio_addrchk_mcast_0_FROM
    );
  rx_input_memio_addrchk_n004925 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_CHOICE1392,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1399,
      O => rx_input_memio_addrchk_lmcast(0)
    );
  rx_input_memio_addrchk_mcast_0_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_mcast_0_CEMUXNOT
    );
  rx_input_memio_addrchk_mcast_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_mcast_0_FROM,
      O => rx_input_memio_addrchk_CHOICE1399
    );
  rx_input_fifo_fifo_BU322 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N4450,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2483_FFY_RST,
      O => rx_input_fifo_fifo_N2484
    );
  rx_input_fifo_fifo_N2483_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2483_FFY_RST
    );
  tx_output_ncrcbyte_7_10 : X_LUT4
    generic map(
      INIT => X"3B0A"
    )
    port map (
      ADR0 => tx_output_crcsell(3),
      ADR1 => tx_output_crcl(23),
      ADR2 => tx_output_crcl(31),
      ADR3 => tx_output_crcsell(2),
      O => tx_output_CHOICE1303_FROM
    );
  tx_output_ncrcbyte_0_10 : X_LUT4
    generic map(
      INIT => X"22F2"
    )
    port map (
      ADR0 => tx_output_crcsell(3),
      ADR1 => tx_output_crcl(24),
      ADR2 => tx_output_crcsell(2),
      ADR3 => tx_output_crcl(16),
      O => tx_output_CHOICE1303_GROM
    );
  tx_output_CHOICE1303_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1303_FROM,
      O => tx_output_CHOICE1303
    );
  tx_output_CHOICE1303_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1303_GROM,
      O => tx_output_CHOICE1380
    );
  tx_output_ncrcbyte_0_21 : X_LUT4
    generic map(
      INIT => X"30BA"
    )
    port map (
      ADR0 => tx_output_crcsell(1),
      ADR1 => tx_output_crcl(0),
      ADR2 => tx_output_crcsell(0),
      ADR3 => tx_output_crcl(8),
      O => tx_output_ncrcbytel_0_FROM
    );
  tx_output_ncrcbyte_0_22 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_CHOICE1380,
      ADR3 => tx_output_CHOICE1385,
      O => tx_output_ncrcbyte(0)
    );
  tx_output_ncrcbytel_0_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_ncrcbytel_0_CEMUXNOT
    );
  tx_output_ncrcbytel_0_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_0_FROM,
      O => tx_output_CHOICE1385
    );
  mac_control_PHY_status_dout_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_15_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(14),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_15_FFY_RST,
      O => mac_control_PHY_status_dout(14)
    );
  tx_output_ncrcbyte_3_10 : X_LUT4
    generic map(
      INIT => X"0CAE"
    )
    port map (
      ADR0 => tx_output_crcsell(3),
      ADR1 => tx_output_crcsell(2),
      ADR2 => tx_output_crcl(19),
      ADR3 => tx_output_crcl(27),
      O => tx_output_CHOICE1336_FROM
    );
  tx_output_ncrcbyte_1_10 : X_LUT4
    generic map(
      INIT => X"0ACE"
    )
    port map (
      ADR0 => tx_output_crcsell(3),
      ADR1 => tx_output_crcsell(2),
      ADR2 => tx_output_crcl(25),
      ADR3 => tx_output_crcl(17),
      O => tx_output_CHOICE1336_GROM
    );
  tx_output_CHOICE1336_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1336_FROM,
      O => tx_output_CHOICE1336
    );
  tx_output_CHOICE1336_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1336_GROM,
      O => tx_output_CHOICE1369
    );
  tx_output_ncrcbyte_1_21 : X_LUT4
    generic map(
      INIT => X"44F4"
    )
    port map (
      ADR0 => tx_output_crcl(9),
      ADR1 => tx_output_crcsell(1),
      ADR2 => tx_output_crcsell(0),
      ADR3 => tx_output_crcl(1),
      O => tx_output_ncrcbytel_1_FROM
    );
  tx_output_ncrcbyte_1_22 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_CHOICE1369,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1374,
      O => tx_output_ncrcbyte(1)
    );
  tx_output_ncrcbytel_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_ncrcbytel_1_CEMUXNOT
    );
  tx_output_ncrcbytel_1_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_1_FROM,
      O => tx_output_CHOICE1374
    );
  mac_control_Ker521611 : X_LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_bitcnt_109,
      ADR2 => mac_control_sclkdeltall,
      ADR3 => mac_control_N52138,
      O => mac_control_N52163_FROM
    );
  mac_control_Mmux_n0017_Result_15_108_SW0 : X_LUT4
    generic map(
      INIT => X"C4CC"
    )
    port map (
      ADR0 => mac_control_sclkdeltall,
      ADR1 => mac_control_dout(14),
      ADR2 => mac_control_bitcnt_109,
      ADR3 => mac_control_N52138,
      O => mac_control_N52163_GROM
    );
  mac_control_N52163_XUSED : X_BUF
    port map (
      I => mac_control_N52163_FROM,
      O => mac_control_N52163
    );
  mac_control_N52163_YUSED : X_BUF
    port map (
      I => mac_control_N52163_GROM,
      O => mac_control_N82001
    );
  tx_output_ncrcbyte_6_10 : X_LUT4
    generic map(
      INIT => X"0CAE"
    )
    port map (
      ADR0 => tx_output_crcsell(3),
      ADR1 => tx_output_crcsell(2),
      ADR2 => tx_output_crcl(22),
      ADR3 => tx_output_crcl(30),
      O => tx_output_CHOICE1314_FROM
    );
  tx_output_ncrcbyte_2_10 : X_LUT4
    generic map(
      INIT => X"2F22"
    )
    port map (
      ADR0 => tx_output_crcsell(3),
      ADR1 => tx_output_crcl(26),
      ADR2 => tx_output_crcl(18),
      ADR3 => tx_output_crcsell(2),
      O => tx_output_CHOICE1314_GROM
    );
  tx_output_CHOICE1314_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1314_FROM,
      O => tx_output_CHOICE1314
    );
  tx_output_CHOICE1314_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1314_GROM,
      O => tx_output_CHOICE1358
    );
  tx_output_ncrcbyte_2_21 : X_LUT4
    generic map(
      INIT => X"5D0C"
    )
    port map (
      ADR0 => tx_output_crcl(2),
      ADR1 => tx_output_crcsell(1),
      ADR2 => tx_output_crcl(10),
      ADR3 => tx_output_crcsell(0),
      O => tx_output_ncrcbytel_2_FROM
    );
  tx_output_ncrcbyte_2_22 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_CHOICE1363,
      ADR3 => tx_output_CHOICE1358,
      O => tx_output_ncrcbyte(2)
    );
  tx_output_ncrcbytel_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_ncrcbytel_2_CEMUXNOT
    );
  tx_output_ncrcbytel_2_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_2_FROM,
      O => tx_output_CHOICE1363
    );
  tx_output_ncrcbyte_3_21 : X_LUT4
    generic map(
      INIT => X"5D0C"
    )
    port map (
      ADR0 => tx_output_crcl(3),
      ADR1 => tx_output_crcsell(1),
      ADR2 => tx_output_crcl(11),
      ADR3 => tx_output_crcsell(0),
      O => tx_output_ncrcbytel_3_FROM
    );
  tx_output_ncrcbyte_3_22 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_CHOICE1336,
      ADR3 => tx_output_CHOICE1341,
      O => tx_output_ncrcbyte(3)
    );
  tx_output_ncrcbytel_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_ncrcbytel_3_CEMUXNOT
    );
  tx_output_ncrcbytel_3_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_3_FROM,
      O => tx_output_CHOICE1341
    );
  tx_output_ncrcbyte_5_10 : X_LUT4
    generic map(
      INIT => X"7350"
    )
    port map (
      ADR0 => tx_output_crcl(29),
      ADR1 => tx_output_crcl(21),
      ADR2 => tx_output_crcsell(3),
      ADR3 => tx_output_crcsell(2),
      O => tx_output_CHOICE1325_FROM
    );
  tx_output_ncrcbyte_4_10 : X_LUT4
    generic map(
      INIT => X"7350"
    )
    port map (
      ADR0 => tx_output_crcl(20),
      ADR1 => tx_output_crcl(28),
      ADR2 => tx_output_crcsell(2),
      ADR3 => tx_output_crcsell(3),
      O => tx_output_CHOICE1325_GROM
    );
  tx_output_CHOICE1325_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1325_FROM,
      O => tx_output_CHOICE1325
    );
  tx_output_CHOICE1325_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1325_GROM,
      O => tx_output_CHOICE1347
    );
  rx_input_memio_crccomb_Mxor_n0005_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0104(0),
      ADR1 => rx_input_memio_crcl(28),
      ADR2 => rx_input_memio_datal(3),
      ADR3 => rx_input_memio_crccomb_n0122(1),
      O => rx_input_memio_crcl_4_FROM
    );
  rx_input_memio_n0048_4_1 : X_LUT4
    generic map(
      INIT => X"CFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => rx_input_memio_crccomb_Mxor_CO_4_Xo_1_1_2,
      ADR3 => rx_input_memio_crccomb_n0056(2),
      O => rx_input_memio_n0048(4)
    );
  rx_input_memio_crcl_4_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_4_FROM,
      O => rx_input_memio_crccomb_n0056(2)
    );
  tx_output_ncrcbyte_4_21 : X_LUT4
    generic map(
      INIT => X"44F4"
    )
    port map (
      ADR0 => tx_output_crcl(12),
      ADR1 => tx_output_crcsell(1),
      ADR2 => tx_output_crcsell(0),
      ADR3 => tx_output_crcl(4),
      O => tx_output_ncrcbytel_4_FROM
    );
  tx_output_ncrcbyte_4_22 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_CHOICE1347,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1352,
      O => tx_output_ncrcbyte(4)
    );
  tx_output_ncrcbytel_4_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_ncrcbytel_4_CEMUXNOT
    );
  tx_output_ncrcbytel_4_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_4_FROM,
      O => tx_output_CHOICE1352
    );
  rx_input_fifo_fifo_BU329 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N4490,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2483_FFX_RST,
      O => rx_input_fifo_fifo_N2483
    );
  rx_input_fifo_fifo_N2483_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2483_FFX_RST
    );
  tx_output_crc_loigc_Mxor_n0004_Result1 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_crcl(27),
      ADR2 => VCC,
      ADR3 => tx_output_data(4),
      O => tx_output_crcl_25_FROM
    );
  tx_output_n0034_25_1 : X_LUT4
    generic map(
      INIT => X"AFFA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => VCC,
      ADR2 => tx_output_crc_loigc_Mxor_CO_25_Xo_1_1_2,
      ADR3 => tx_output_crc_loigc_n0124(1),
      O => tx_output_n0034(25)
    );
  tx_output_crcl_25_XUSED : X_BUF
    port map (
      I => tx_output_crcl_25_FROM,
      O => tx_output_crc_loigc_n0124(1)
    );
  rx_input_fifo_fifo_BU380 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2404,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2423_FFY_RST,
      O => rx_input_fifo_fifo_N2424
    );
  rx_input_fifo_fifo_N2423_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2423_FFY_RST
    );
  tx_output_ncrcbyte_5_21 : X_LUT4
    generic map(
      INIT => X"5D0C"
    )
    port map (
      ADR0 => tx_output_crcl(13),
      ADR1 => tx_output_crcsell(0),
      ADR2 => tx_output_crcl(5),
      ADR3 => tx_output_crcsell(1),
      O => tx_output_ncrcbytel_5_FROM
    );
  tx_output_ncrcbyte_5_22 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_CHOICE1325,
      ADR3 => tx_output_CHOICE1330,
      O => tx_output_ncrcbyte(5)
    );
  tx_output_ncrcbytel_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_ncrcbytel_5_CEMUXNOT
    );
  tx_output_ncrcbytel_5_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_5_FROM,
      O => tx_output_CHOICE1330
    );
  tx_output_ncrcbyte_6_21 : X_LUT4
    generic map(
      INIT => X"4F44"
    )
    port map (
      ADR0 => tx_output_crcl(14),
      ADR1 => tx_output_crcsell(1),
      ADR2 => tx_output_crcl(6),
      ADR3 => tx_output_crcsell(0),
      O => tx_output_ncrcbytel_6_FROM
    );
  tx_output_ncrcbyte_6_22 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_CHOICE1314,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1319,
      O => tx_output_ncrcbyte(6)
    );
  tx_output_ncrcbytel_6_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_ncrcbytel_6_CEMUXNOT
    );
  tx_output_ncrcbytel_6_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_6_FROM,
      O => tx_output_CHOICE1319
    );
  rx_input_memio_addrchk_n0051_2_103 : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_bcast(4),
      ADR2 => rx_input_memio_addrchk_bcast(0),
      ADR3 => rx_input_memio_addrchk_bcast(5),
      O => rx_input_memio_addrchk_validbcast_FROM
    );
  rx_input_memio_addrchk_n0051_104 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_bcast(3),
      ADR1 => rx_input_memio_addrchk_bcast(2),
      ADR2 => rx_input_memio_addrchk_bcast(1),
      ADR3 => rx_input_memio_addrchk_n0051_2,
      O => rx_input_memio_addrchk_n0051
    );
  rx_input_memio_addrchk_validbcast_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_validbcast_CEMUXNOT
    );
  rx_input_memio_addrchk_validbcast_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_validbcast_FROM,
      O => rx_input_memio_addrchk_n0051_2
    );
  rx_input_fifo_fifo_BU264 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3938,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N9_FFY_RST,
      O => rx_input_fifo_fifo_N8
    );
  rx_input_fifo_fifo_N9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N9_FFY_RST
    );
  tx_output_ncrcbyte_7_21 : X_LUT4
    generic map(
      INIT => X"7350"
    )
    port map (
      ADR0 => tx_output_crcl(7),
      ADR1 => tx_output_crcl(15),
      ADR2 => tx_output_crcsell(0),
      ADR3 => tx_output_crcsell(1),
      O => tx_output_ncrcbytel_7_FROM
    );
  tx_output_ncrcbyte_7_22 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_CHOICE1303,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1308,
      O => tx_output_ncrcbyte(7)
    );
  tx_output_ncrcbytel_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_ncrcbytel_7_CEMUXNOT
    );
  tx_output_ncrcbytel_7_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_7_FROM,
      O => tx_output_CHOICE1308
    );
  rx_input_memio_addrchk_n0052_2_105 : X_LUT4
    generic map(
      INIT => X"8800"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_maceq(4),
      ADR1 => rx_input_memio_addrchk_maceq(0),
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_maceq(5),
      O => rx_input_memio_addrchk_validucast_FROM
    );
  rx_input_memio_addrchk_n0052_106 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_maceq(2),
      ADR1 => rx_input_memio_addrchk_maceq(3),
      ADR2 => rx_input_memio_addrchk_maceq(1),
      ADR3 => rx_input_memio_addrchk_n0052_2,
      O => rx_input_memio_addrchk_n0052
    );
  rx_input_memio_addrchk_validucast_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_validucast_CEMUXNOT
    );
  rx_input_memio_addrchk_validucast_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_validucast_FROM,
      O => rx_input_memio_addrchk_n0052_2
    );
  rx_fifocheck_n000212 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(0),
      ADR1 => rx_fifocheck_diff(3),
      ADR2 => rx_fifocheck_diff(1),
      ADR3 => rx_fifocheck_diff(2),
      O => rx_fifocheck_CHOICE1774_GROM
    );
  rx_fifocheck_CHOICE1774_YUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1774_GROM,
      O => rx_fifocheck_CHOICE1774
    );
  rx_fifocheck_n000225 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(4),
      ADR1 => rx_fifocheck_diff(5),
      ADR2 => rx_fifocheck_diff(6),
      ADR3 => rx_fifocheck_diff(7),
      O => rx_fifocheck_CHOICE1781_GROM
    );
  rx_fifocheck_CHOICE1781_YUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1781_GROM,
      O => rx_fifocheck_CHOICE1781
    );
  rx_fifocheck_n000262 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(15),
      ADR1 => rx_fifocheck_diff(14),
      ADR2 => rx_fifocheck_diff(13),
      ADR3 => rx_fifocheck_diff(12),
      O => rx_fifocheck_CHOICE1796_GROM
    );
  rx_fifocheck_CHOICE1796_YUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1796_GROM,
      O => rx_fifocheck_CHOICE1796
    );
  mac_control_LEDDPX_OBUF_107 : X_TRI
    port map (
      I => LEDDPX_OUTMUX,
      CTL => LEDDPX_ENABLE,
      O => LEDDPX
    );
  LEDDPX_ENABLEINV : X_INV
    port map (
      I => LEDDPX_TORGTS,
      O => LEDDPX_ENABLE
    );
  LEDDPX_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDDPX_TORGTS
    );
  LEDDPX_OUTMUX_108 : X_BUF
    port map (
      I => mac_control_LEDDPX_OBUF,
      O => LEDDPX_OUTMUX
    );
  LEDDPX_OMUX : X_BUF
    port map (
      I => mac_control_phystat(1),
      O => LEDDPX_OD
    );
  rx_input_GMII_RXD_0_IBUF_109 : X_BUF
    port map (
      I => RXD(0),
      O => rx_input_GMII_RXD_0_IBUF
    );
  rx_input_GMII_RXD_1_IBUF_110 : X_BUF
    port map (
      I => RXD(1),
      O => rx_input_GMII_RXD_1_IBUF
    );
  rx_input_GMII_RXD_2_IBUF_111 : X_BUF
    port map (
      I => RXD(2),
      O => rx_input_GMII_RXD_2_IBUF
    );
  rx_input_GMII_RXD_3_IBUF_112 : X_BUF
    port map (
      I => RXD(3),
      O => rx_input_GMII_RXD_3_IBUF
    );
  rx_input_GMII_RXD_4_IBUF_113 : X_BUF
    port map (
      I => RXD(4),
      O => rx_input_GMII_RXD_4_IBUF
    );
  rx_input_GMII_RXD_5_IBUF_114 : X_BUF
    port map (
      I => RXD(5),
      O => rx_input_GMII_RXD_5_IBUF
    );
  rx_input_GMII_RXD_6_IBUF_115 : X_BUF
    port map (
      I => RXD(6),
      O => rx_input_GMII_RXD_6_IBUF
    );
  rx_input_GMII_RXD_7_IBUF_116 : X_BUF
    port map (
      I => RXD(7),
      O => rx_input_GMII_RXD_7_IBUF
    );
  tx_input_DIN_10_IBUF_117 : X_BUF
    port map (
      I => DIN(10),
      O => tx_input_DIN_10_IBUF
    );
  tx_input_DIN_11_IBUF_118 : X_BUF
    port map (
      I => DIN(11),
      O => tx_input_DIN_11_IBUF
    );
  tx_input_DIN_12_IBUF_119 : X_BUF
    port map (
      I => DIN(12),
      O => tx_input_DIN_12_IBUF
    );
  tx_input_DIN_13_IBUF_120 : X_BUF
    port map (
      I => DIN(13),
      O => tx_input_DIN_13_IBUF
    );
  tx_input_DIN_14_IBUF_121 : X_BUF
    port map (
      I => DIN(14),
      O => tx_input_DIN_14_IBUF
    );
  tx_input_DIN_15_IBUF_122 : X_BUF
    port map (
      I => DIN(15),
      O => tx_input_DIN_15_IBUF
    );
  rx_output_DOUT_0_OBUF_123 : X_TRI
    port map (
      I => DOUT_0_OUTMUX,
      CTL => DOUT_0_ENABLE,
      O => DOUT(0)
    );
  DOUT_0_ENABLEINV : X_INV
    port map (
      I => DOUT_0_TORGTS,
      O => DOUT_0_ENABLE
    );
  DOUT_0_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_0_TORGTS
    );
  DOUT_0_OUTMUX_124 : X_BUF
    port map (
      I => rx_output_DOUT_0_OBUF,
      O => DOUT_0_OUTMUX
    );
  DOUT_0_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(0),
      O => DOUT_0_OD
    );
  rx_output_DOUT_1_OBUF_125 : X_TRI
    port map (
      I => DOUT_1_OUTMUX,
      CTL => DOUT_1_ENABLE,
      O => DOUT(1)
    );
  DOUT_1_ENABLEINV : X_INV
    port map (
      I => DOUT_1_TORGTS,
      O => DOUT_1_ENABLE
    );
  DOUT_1_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_1_TORGTS
    );
  DOUT_1_OUTMUX_126 : X_BUF
    port map (
      I => rx_output_DOUT_1_OBUF,
      O => DOUT_1_OUTMUX
    );
  DOUT_1_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(1),
      O => DOUT_1_OD
    );
  rx_input_fifo_fifo_BU178 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3600,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N2397_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2397
    );
  rx_input_fifo_fifo_N2397_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2397_FFX_SET
    );
  rx_output_DOUT_2_OBUF_127 : X_TRI
    port map (
      I => DOUT_2_OUTMUX,
      CTL => DOUT_2_ENABLE,
      O => DOUT(2)
    );
  DOUT_2_ENABLEINV : X_INV
    port map (
      I => DOUT_2_TORGTS,
      O => DOUT_2_ENABLE
    );
  DOUT_2_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_2_TORGTS
    );
  DOUT_2_OUTMUX_128 : X_BUF
    port map (
      I => rx_output_DOUT_2_OBUF,
      O => DOUT_2_OUTMUX
    );
  DOUT_2_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(2),
      O => DOUT_2_OD
    );
  rx_output_DOUT_3_OBUF_129 : X_TRI
    port map (
      I => DOUT_3_OUTMUX,
      CTL => DOUT_3_ENABLE,
      O => DOUT(3)
    );
  DOUT_3_ENABLEINV : X_INV
    port map (
      I => DOUT_3_TORGTS,
      O => DOUT_3_ENABLE
    );
  DOUT_3_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_3_TORGTS
    );
  DOUT_3_OUTMUX_130 : X_BUF
    port map (
      I => rx_output_DOUT_3_OBUF,
      O => DOUT_3_OUTMUX
    );
  DOUT_3_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(3),
      O => DOUT_3_OD
    );
  rx_output_DOUT_4_OBUF_131 : X_TRI
    port map (
      I => DOUT_4_OUTMUX,
      CTL => DOUT_4_ENABLE,
      O => DOUT(4)
    );
  DOUT_4_ENABLEINV : X_INV
    port map (
      I => DOUT_4_TORGTS,
      O => DOUT_4_ENABLE
    );
  DOUT_4_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_4_TORGTS
    );
  DOUT_4_OUTMUX_132 : X_BUF
    port map (
      I => rx_output_DOUT_4_OBUF,
      O => DOUT_4_OUTMUX
    );
  DOUT_4_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(4),
      O => DOUT_4_OD
    );
  rx_output_DOUT_5_OBUF_133 : X_TRI
    port map (
      I => DOUT_5_OUTMUX,
      CTL => DOUT_5_ENABLE,
      O => DOUT(5)
    );
  DOUT_5_ENABLEINV : X_INV
    port map (
      I => DOUT_5_TORGTS,
      O => DOUT_5_ENABLE
    );
  DOUT_5_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_5_TORGTS
    );
  DOUT_5_OUTMUX_134 : X_BUF
    port map (
      I => rx_output_DOUT_5_OBUF,
      O => DOUT_5_OUTMUX
    );
  DOUT_5_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(5),
      O => DOUT_5_OD
    );
  rx_output_DOUT_6_OBUF_135 : X_TRI
    port map (
      I => DOUT_6_OUTMUX,
      CTL => DOUT_6_ENABLE,
      O => DOUT(6)
    );
  DOUT_6_ENABLEINV : X_INV
    port map (
      I => DOUT_6_TORGTS,
      O => DOUT_6_ENABLE
    );
  DOUT_6_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_6_TORGTS
    );
  DOUT_6_OUTMUX_136 : X_BUF
    port map (
      I => rx_output_DOUT_6_OBUF,
      O => DOUT_6_OUTMUX
    );
  DOUT_6_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(6),
      O => DOUT_6_OD
    );
  rx_output_DOUT_7_OBUF_137 : X_TRI
    port map (
      I => DOUT_7_OUTMUX,
      CTL => DOUT_7_ENABLE,
      O => DOUT(7)
    );
  DOUT_7_ENABLEINV : X_INV
    port map (
      I => DOUT_7_TORGTS,
      O => DOUT_7_ENABLE
    );
  DOUT_7_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_7_TORGTS
    );
  DOUT_7_OUTMUX_138 : X_BUF
    port map (
      I => rx_output_DOUT_7_OBUF,
      O => DOUT_7_OUTMUX
    );
  DOUT_7_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(7),
      O => DOUT_7_OD
    );
  rx_output_DOUT_8_OBUF_139 : X_TRI
    port map (
      I => DOUT_8_OUTMUX,
      CTL => DOUT_8_ENABLE,
      O => DOUT(8)
    );
  DOUT_8_ENABLEINV : X_INV
    port map (
      I => DOUT_8_TORGTS,
      O => DOUT_8_ENABLE
    );
  DOUT_8_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_8_TORGTS
    );
  DOUT_8_OUTMUX_140 : X_BUF
    port map (
      I => rx_output_DOUT_8_OBUF,
      O => DOUT_8_OUTMUX
    );
  DOUT_8_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(8),
      O => DOUT_8_OD
    );
  rx_input_fifo_fifo_BU211 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2478,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2499_FFY_RST,
      O => rx_input_fifo_fifo_N2498
    );
  rx_input_fifo_fifo_N2499_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2499_FFY_RST
    );
  rx_output_DOUT_9_OBUF_141 : X_TRI
    port map (
      I => DOUT_9_OUTMUX,
      CTL => DOUT_9_ENABLE,
      O => DOUT(9)
    );
  DOUT_9_ENABLEINV : X_INV
    port map (
      I => DOUT_9_TORGTS,
      O => DOUT_9_ENABLE
    );
  DOUT_9_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_9_TORGTS
    );
  DOUT_9_OUTMUX_142 : X_BUF
    port map (
      I => rx_output_DOUT_9_OBUF,
      O => DOUT_9_OUTMUX
    );
  DOUT_9_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(9),
      O => DOUT_9_OD
    );
  mac_control_SOUT_OBUF_143 : X_TRI
    port map (
      I => SOUT_OUTMUX,
      CTL => SOUT_ENABLE,
      O => SOUT
    );
  SOUT_ENABLEINV : X_INV
    port map (
      I => SOUT_TORGTS,
      O => SOUT_ENABLE
    );
  SOUT_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => SOUT_TORGTS
    );
  SOUT_OUTMUX_144 : X_BUF
    port map (
      I => mac_control_SOUT_OBUF,
      O => SOUT_OUTMUX
    );
  SOUT_OMUX : X_BUF
    port map (
      I => mac_control_dout(31),
      O => SOUT_OD
    );
  mac_control_SCLK_IBUF_145 : X_BUF
    port map (
      I => SCLK,
      O => mac_control_SCLK_IBUF
    );
  mac_control_LEDRX_OBUF_146 : X_TRI
    port map (
      I => LEDRX_OUTMUX,
      CTL => LEDRX_ENABLE,
      O => LEDRX
    );
  LEDRX_ENABLEINV : X_INV
    port map (
      I => LEDRX_TORGTS,
      O => LEDRX_ENABLE
    );
  LEDRX_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDRX_TORGTS
    );
  LEDRX_OUTMUX_147 : X_BUF
    port map (
      I => mac_control_LEDRX_OBUF,
      O => LEDRX_OUTMUX
    );
  LEDRX_OMUX : X_BUF
    port map (
      I => mac_control_n0041,
      O => LEDRX_OD
    );
  mac_control_LEDTX_OBUF_148 : X_TRI
    port map (
      I => LEDTX_OUTMUX,
      CTL => LEDTX_ENABLE,
      O => LEDTX
    );
  LEDTX_ENABLEINV : X_INV
    port map (
      I => LEDTX_TORGTS,
      O => LEDTX_ENABLE
    );
  LEDTX_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDTX_TORGTS
    );
  LEDTX_OUTMUX_149 : X_BUF
    port map (
      I => mac_control_LEDTX_OBUF,
      O => LEDTX_OUTMUX
    );
  LEDTX_OMUX : X_BUF
    port map (
      I => mac_control_n0039,
      O => LEDTX_OD
    );
  tx_input_DIN_0_IBUF_150 : X_BUF
    port map (
      I => DIN(0),
      O => tx_input_DIN_0_IBUF
    );
  tx_input_DIN_1_IBUF_151 : X_BUF
    port map (
      I => DIN(1),
      O => tx_input_DIN_1_IBUF
    );
  tx_input_DIN_2_IBUF_152 : X_BUF
    port map (
      I => DIN(2),
      O => tx_input_DIN_2_IBUF
    );
  tx_input_DIN_3_IBUF_153 : X_BUF
    port map (
      I => DIN(3),
      O => tx_input_DIN_3_IBUF
    );
  tx_input_DIN_4_IBUF_154 : X_BUF
    port map (
      I => DIN(4),
      O => tx_input_DIN_4_IBUF
    );
  tx_input_DIN_5_IBUF_155 : X_BUF
    port map (
      I => DIN(5),
      O => tx_input_DIN_5_IBUF
    );
  tx_input_DIN_6_IBUF_156 : X_BUF
    port map (
      I => DIN(6),
      O => tx_input_DIN_6_IBUF
    );
  rx_input_fifo_fifo_BU164 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3520,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2400_FFY_RST,
      O => rx_input_fifo_fifo_N2399
    );
  rx_input_fifo_fifo_N2400_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2400_FFY_RST
    );
  tx_input_DIN_7_IBUF_157 : X_BUF
    port map (
      I => DIN(7),
      O => tx_input_DIN_7_IBUF
    );
  tx_input_DIN_8_IBUF_158 : X_BUF
    port map (
      I => DIN(8),
      O => tx_input_DIN_8_IBUF
    );
  tx_input_DIN_9_IBUF_159 : X_BUF
    port map (
      I => DIN(9),
      O => tx_input_DIN_9_IBUF
    );
  rx_input_GMII_RX_ER_IBUF_160 : X_BUF
    port map (
      I => RX_ER,
      O => rx_input_GMII_RX_ER_IBUF
    );
  rx_input_GMII_RX_DV_IBUF_161 : X_BUF
    port map (
      I => RX_DV,
      O => rx_input_GMII_RX_DV_IBUF
    );
  memcontroller_MA_10_OBUF : X_TRI
    port map (
      I => MA_10_OUTMUX,
      CTL => MA_10_ENABLE,
      O => MA(10)
    );
  MA_10_ENABLEINV : X_INV
    port map (
      I => MA_10_TORGTS,
      O => MA_10_ENABLE
    );
  MA_10_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_10_TORGTS
    );
  MA_10_OUTMUX_162 : X_BUF
    port map (
      I => memcontroller_ADDREXT(10),
      O => MA_10_OUTMUX
    );
  MA_10_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_10_OCEMUXNOT
    );
  MA_10_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(10),
      O => MA_10_OD
    );
  rx_input_fifo_fifo_BU101 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2813,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N13_FFX_RST,
      O => rx_input_fifo_fifo_N13
    );
  rx_input_fifo_fifo_N13_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N13_FFX_RST
    );
  memcontroller_MA_11_OBUF : X_TRI
    port map (
      I => MA_11_OUTMUX,
      CTL => MA_11_ENABLE,
      O => MA(11)
    );
  MA_11_ENABLEINV : X_INV
    port map (
      I => MA_11_TORGTS,
      O => MA_11_ENABLE
    );
  MA_11_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_11_TORGTS
    );
  MA_11_OUTMUX_163 : X_BUF
    port map (
      I => memcontroller_ADDREXT(11),
      O => MA_11_OUTMUX
    );
  MA_11_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_11_OCEMUXNOT
    );
  MA_11_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(11),
      O => MA_11_OD
    );
  memcontroller_MA_12_OBUF : X_TRI
    port map (
      I => MA_12_OUTMUX,
      CTL => MA_12_ENABLE,
      O => MA(12)
    );
  MA_12_ENABLEINV : X_INV
    port map (
      I => MA_12_TORGTS,
      O => MA_12_ENABLE
    );
  MA_12_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_12_TORGTS
    );
  MA_12_OUTMUX_164 : X_BUF
    port map (
      I => memcontroller_ADDREXT(12),
      O => MA_12_OUTMUX
    );
  MA_12_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_12_OCEMUXNOT
    );
  MA_12_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(12),
      O => MA_12_OD
    );
  mac_control_n00371 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_phystat(3),
      ADR3 => mac_control_phystat(4),
      O => mac_control_n0037_FROM
    );
  mac_control_n00361 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phystat(3),
      ADR2 => mac_control_phystat(4),
      ADR3 => VCC,
      O => mac_control_n0037_GROM
    );
  mac_control_n0037_XUSED : X_BUF
    port map (
      I => mac_control_n0037_FROM,
      O => mac_control_n0037
    );
  mac_control_n0037_YUSED : X_BUF
    port map (
      I => mac_control_n0037_GROM,
      O => mac_control_n0036
    );
  mac_control_n00441 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => mac_control_rxf_rst,
      ADR1 => clkslen,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_n0044_GROM
    );
  mac_control_n0044_YUSED : X_BUF
    port map (
      I => mac_control_n0044_GROM,
      O => mac_control_n0044
    );
  mac_control_n00531 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => rxoferrsr,
      ADR1 => VCC,
      ADR2 => clkslen,
      ADR3 => VCC,
      O => mac_control_n0053_GROM
    );
  mac_control_n0053_YUSED : X_BUF
    port map (
      I => mac_control_n0053_GROM,
      O => mac_control_n0053
    );
  mac_control_n00451 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rxfsr,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => clkslen,
      O => mac_control_n0045_GROM
    );
  mac_control_n0045_YUSED : X_BUF
    port map (
      I => mac_control_n0045_GROM,
      O => mac_control_n0045
    );
  rx_input_fifo_fifo_BU444 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N9,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2473_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2474
    );
  rx_input_fifo_fifo_N2473_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2473_FFY_SET
    );
  mac_control_n00541 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => clkslen,
      ADR3 => mac_control_rxcrcerr_rst,
      O => mac_control_n0054_GROM
    );
  mac_control_n0054_YUSED : X_BUF
    port map (
      I => mac_control_n0054_GROM,
      O => mac_control_n0054
    );
  mac_control_n00461 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_rst,
      ADR2 => clkslen,
      ADR3 => VCC,
      O => mac_control_n0046_GROM
    );
  mac_control_n0046_YUSED : X_BUF
    port map (
      I => mac_control_n0046_GROM,
      O => mac_control_n0046
    );
  mac_control_n00551 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rxcrcerrsr,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => clkslen,
      O => mac_control_n0055_GROM
    );
  mac_control_n0055_YUSED : X_BUF
    port map (
      I => mac_control_n0055_GROM,
      O => mac_control_n0055
    );
  mac_control_n00471 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => clkslen,
      ADR2 => txfifowerrsr,
      ADR3 => VCC,
      O => mac_control_n0047_GROM
    );
  mac_control_n0047_YUSED : X_BUF
    port map (
      I => mac_control_n0047_GROM,
      O => mac_control_n0047
    );
  mac_control_n00481 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_rst,
      ADR1 => VCC,
      ADR2 => clkslen,
      ADR3 => VCC,
      O => mac_control_n0048_GROM
    );
  mac_control_n0048_YUSED : X_BUF
    port map (
      I => mac_control_n0048_GROM,
      O => mac_control_n0048
    );
  mac_control_n00801 : X_LUT4
    generic map(
      INIT => X"0008"
    )
    port map (
      ADR0 => mac_control_addr(4),
      ADR1 => mac_control_N52244,
      ADR2 => mac_control_addr(3),
      ADR3 => mac_control_addr(2),
      O => mac_control_n0080_FROM
    );
  mac_control_Mmux_n0017_Result_3_74 : X_LUT4
    generic map(
      INIT => X"FEFA"
    )
    port map (
      ADR0 => mac_control_CHOICE2801,
      ADR1 => mac_control_txfifowerr_cnt(3),
      ADR2 => mac_control_N81693,
      ADR3 => mac_control_n0080,
      O => mac_control_n0080_GROM
    );
  mac_control_n0080_XUSED : X_BUF
    port map (
      I => mac_control_n0080_FROM,
      O => mac_control_n0080
    );
  mac_control_n0080_YUSED : X_BUF
    port map (
      I => mac_control_n0080_GROM,
      O => mac_control_CHOICE2810
    );
  mac_control_n00491 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => clkslen,
      ADR1 => rxfifowerrsr,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_n0049_GROM
    );
  mac_control_n0049_YUSED : X_BUF
    port map (
      I => mac_control_n0049_GROM,
      O => mac_control_n0049
    );
  mac_control_Ker52151_SW0 : X_LUT4
    generic map(
      INIT => X"0010"
    )
    port map (
      ADR0 => mac_control_addr(4),
      ADR1 => mac_control_addr(2),
      ADR2 => mac_control_din(0),
      ADR3 => mac_control_addr(3),
      O => mac_control_N69420_FROM
    );
  mac_control_n00731 : X_LUT4
    generic map(
      INIT => X"0010"
    )
    port map (
      ADR0 => mac_control_addr(4),
      ADR1 => mac_control_addr(2),
      ADR2 => mac_control_N52228,
      ADR3 => mac_control_addr(3),
      O => mac_control_N69420_GROM
    );
  mac_control_N69420_XUSED : X_BUF
    port map (
      I => mac_control_N69420_FROM,
      O => mac_control_N69420
    );
  mac_control_N69420_YUSED : X_BUF
    port map (
      I => mac_control_N69420_GROM,
      O => mac_control_n0073
    );
  mac_control_n00811 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => mac_control_N52236,
      ADR1 => mac_control_addr(4),
      ADR2 => mac_control_addr(3),
      ADR3 => mac_control_addr(2),
      O => mac_control_n0081_FROM
    );
  mac_control_Mmux_n0017_Result_30_7 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(30),
      ADR1 => mac_control_rxfifowerr_cnt(30),
      ADR2 => mac_control_n0080,
      ADR3 => mac_control_n0081,
      O => mac_control_n0081_GROM
    );
  mac_control_n0081_XUSED : X_BUF
    port map (
      I => mac_control_n0081_FROM,
      O => mac_control_n0081
    );
  mac_control_n0081_YUSED : X_BUF
    port map (
      I => mac_control_n0081_GROM,
      O => mac_control_CHOICE2054
    );
  mac_control_n00851 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_addr(4),
      ADR1 => mac_control_addr(2),
      ADR2 => mac_control_N52220,
      ADR3 => mac_control_addr(3),
      O => mac_control_n0085_FROM
    );
  mac_control_n00741 : X_LUT4
    generic map(
      INIT => X"0010"
    )
    port map (
      ADR0 => mac_control_addr(3),
      ADR1 => mac_control_addr(2),
      ADR2 => mac_control_N52244,
      ADR3 => mac_control_addr(4),
      O => mac_control_n0085_GROM
    );
  mac_control_n0085_XUSED : X_BUF
    port map (
      I => mac_control_n0085_FROM,
      O => mac_control_n0085
    );
  mac_control_n0085_YUSED : X_BUF
    port map (
      I => mac_control_n0085_GROM,
      O => mac_control_n0074
    );
  mac_control_n00581 : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_sclkdeltal,
      ADR2 => mac_control_bitcnt_109,
      ADR3 => mac_control_N52138,
      O => mac_control_txf_rst_FROM
    );
  mac_control_n00621 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_N52236,
      ADR1 => mac_control_din(0),
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_newcmd,
      O => mac_control_n0062
    );
  mac_control_txf_rst_XUSED : X_BUF
    port map (
      I => mac_control_txf_rst_FROM,
      O => mac_control_newcmd
    );
  mac_control_n00821 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => mac_control_addr(3),
      ADR1 => mac_control_addr(4),
      ADR2 => mac_control_N52220,
      ADR3 => mac_control_addr(2),
      O => mac_control_n0082_FROM
    );
  mac_control_Mmux_n0017_Result_9_45 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(9),
      ADR1 => mac_control_n0081,
      ADR2 => mac_control_rxphyerr_cnt(9),
      ADR3 => mac_control_n0082,
      O => mac_control_n0082_GROM
    );
  mac_control_n0082_XUSED : X_BUF
    port map (
      I => mac_control_n0082_FROM,
      O => mac_control_n0082
    );
  mac_control_n0082_YUSED : X_BUF
    port map (
      I => mac_control_n0082_GROM,
      O => mac_control_CHOICE2645
    );
  mac_control_n00831 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => mac_control_addr(4),
      ADR1 => mac_control_addr(3),
      ADR2 => mac_control_addr(2),
      ADR3 => mac_control_N52228,
      O => mac_control_n0083_FROM
    );
  mac_control_Mmux_n0017_Result_3_48 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(3),
      ADR1 => mac_control_rxoferr_cnt(3),
      ADR2 => mac_control_n0082,
      ADR3 => mac_control_n0083,
      O => mac_control_n0083_GROM
    );
  mac_control_n0083_XUSED : X_BUF
    port map (
      I => mac_control_n0083_FROM,
      O => mac_control_n0083
    );
  mac_control_n0083_YUSED : X_BUF
    port map (
      I => mac_control_n0083_GROM,
      O => mac_control_CHOICE2801
    );
  rx_input_fifo_fifo_BU560 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N5343,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2453_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2454
    );
  rx_input_fifo_fifo_N2453_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2453_FFY_SET
    );
  mac_control_n00761 : X_LUT4
    generic map(
      INIT => X"0020"
    )
    port map (
      ADR0 => mac_control_N52220,
      ADR1 => mac_control_addr(4),
      ADR2 => mac_control_addr(3),
      ADR3 => mac_control_addr(2),
      O => mac_control_n0076_FROM
    );
  mac_control_Mmux_n0017_Result_30_29 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0073,
      ADR1 => mac_control_phydi(30),
      ADR2 => mac_control_phystat(30),
      ADR3 => mac_control_n0076,
      O => mac_control_n0076_GROM
    );
  mac_control_n0076_XUSED : X_BUF
    port map (
      I => mac_control_n0076_FROM,
      O => mac_control_n0076
    );
  mac_control_n0076_YUSED : X_BUF
    port map (
      I => mac_control_n0076_GROM,
      O => mac_control_CHOICE2064
    );
  mac_control_n00841 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => mac_control_N52244,
      ADR1 => mac_control_addr(4),
      ADR2 => mac_control_addr(3),
      ADR3 => mac_control_addr(2),
      O => mac_control_n0084_FROM
    );
  mac_control_Mmux_n0017_Result_13_57 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxoferr_cnt(13),
      ADR1 => mac_control_rxcrcerr_cnt(13),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_n0084,
      O => mac_control_n0084_GROM
    );
  mac_control_n0084_XUSED : X_BUF
    port map (
      I => mac_control_n0084_FROM,
      O => mac_control_n0084
    );
  mac_control_n0084_YUSED : X_BUF
    port map (
      I => mac_control_n0084_GROM,
      O => mac_control_CHOICE2711
    );
  mac_control_n00771 : X_LUT4
    generic map(
      INIT => X"0400"
    )
    port map (
      ADR0 => mac_control_addr(4),
      ADR1 => mac_control_N52228,
      ADR2 => mac_control_addr(2),
      ADR3 => mac_control_addr(3),
      O => mac_control_n0077_FROM
    );
  mac_control_Mmux_n0017_Result_3_15 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0076,
      ADR1 => mac_control_phydo(3),
      ADR2 => mac_control_phydi(3),
      ADR3 => mac_control_n0077,
      O => mac_control_n0077_GROM
    );
  mac_control_n0077_XUSED : X_BUF
    port map (
      I => mac_control_n0077_FROM,
      O => mac_control_n0077
    );
  mac_control_n0077_YUSED : X_BUF
    port map (
      I => mac_control_n0077_GROM,
      O => mac_control_CHOICE2790
    );
  mac_control_n00871 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => mac_control_N52143,
      ADR1 => mac_control_addr(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_n0087_FROM
    );
  mac_control_n00861 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N52143,
      ADR2 => mac_control_addr(0),
      ADR3 => VCC,
      O => mac_control_n0087_GROM
    );
  mac_control_n0087_XUSED : X_BUF
    port map (
      I => mac_control_n0087_FROM,
      O => mac_control_n0087
    );
  mac_control_n0087_YUSED : X_BUF
    port map (
      I => mac_control_n0087_GROM,
      O => mac_control_n0086
    );
  mac_control_n00791 : X_LUT4
    generic map(
      INIT => X"0200"
    )
    port map (
      ADR0 => mac_control_addr(4),
      ADR1 => mac_control_addr(3),
      ADR2 => mac_control_addr(2),
      ADR3 => mac_control_N52228,
      O => mac_control_n0079_FROM
    );
  mac_control_Mmux_n0017_Result_3_20 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(3),
      ADR1 => mac_control_n0078,
      ADR2 => mac_control_txf_cnt(3),
      ADR3 => mac_control_n0079,
      O => mac_control_n0079_GROM
    );
  mac_control_n0079_XUSED : X_BUF
    port map (
      I => mac_control_n0079_FROM,
      O => mac_control_n0079
    );
  mac_control_n0079_YUSED : X_BUF
    port map (
      I => mac_control_n0079_GROM,
      O => mac_control_CHOICE2793
    );
  mac_control_Mmux_n0017_Result_4_7 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_lmacaddr(36),
      ADR1 => mac_control_n0087,
      ADR2 => mac_control_n0103,
      ADR3 => mac_control_phyaddr(4),
      O => mac_control_CHOICE2600_FROM
    );
  mac_control_Mmux_n0017_Result_11_30_SW0 : X_LUT4
    generic map(
      INIT => X"FEFA"
    )
    port map (
      ADR0 => mac_control_CHOICE2857,
      ADR1 => mac_control_phyaddr(11),
      ADR2 => mac_control_CHOICE2854,
      ADR3 => mac_control_n0103,
      O => mac_control_CHOICE2600_GROM
    );
  mac_control_CHOICE2600_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2600_FROM,
      O => mac_control_CHOICE2600
    );
  mac_control_CHOICE2600_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2600_GROM,
      O => mac_control_N81785
    );
  rx_input_fifo_fifo_BU468 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2403,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2443_FFX_RST,
      O => rx_input_fifo_fifo_N2443
    );
  rx_input_fifo_fifo_N2443_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2443_FFX_RST
    );
  mac_control_Mmux_n0017_Result_27_103_SW1 : X_LUT4
    generic map(
      INIT => X"0007"
    )
    port map (
      ADR0 => mac_control_N52132,
      ADR1 => mac_control_CHOICE1901,
      ADR2 => mac_control_CHOICE1898,
      ADR3 => mac_control_CHOICE1905,
      O => mac_control_dout_27_FROM
    );
  mac_control_Mmux_n0017_Result_27_103 : X_LUT4
    generic map(
      INIT => X"5072"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_addr(5),
      ADR2 => mac_control_dout(26),
      ADR3 => mac_control_N82086,
      O => mac_control_N74720
    );
  mac_control_dout_27_XUSED : X_BUF
    port map (
      I => mac_control_dout_27_FROM,
      O => mac_control_N82086
    );
  mac_control_Mmux_n0017_Result_19_103_SW1 : X_LUT4
    generic map(
      INIT => X"0103"
    )
    port map (
      ADR0 => mac_control_CHOICE1845,
      ADR1 => mac_control_CHOICE1842,
      ADR2 => mac_control_CHOICE1849,
      ADR3 => mac_control_N52132,
      O => mac_control_dout_19_FROM
    );
  mac_control_Mmux_n0017_Result_19_103 : X_LUT4
    generic map(
      INIT => X"0C5C"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_dout(18),
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_N82078,
      O => mac_control_N74424
    );
  mac_control_dout_19_XUSED : X_BUF
    port map (
      I => mac_control_dout_19_FROM,
      O => mac_control_N82078
    );
  mac_control_PHY_status_MII_Interface_sts28 : X_LUT4
    generic map(
      INIT => X"2237"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR1 => mac_control_PHY_status_miirw,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR3 => mac_control_PHY_status_MII_Interface_N81600,
      O => mac_control_PHY_status_MII_Interface_CHOICE1201_FROM
    );
  mac_control_PHY_status_MII_Interface_sts35 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(5),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE1201,
      O => mac_control_PHY_status_MII_Interface_CHOICE1201_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE1201_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE1201_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE1201
    );
  mac_control_PHY_status_MII_Interface_CHOICE1201_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE1201_GROM,
      O => mac_control_PHY_status_MII_Interface_sts
    );
  mac_control_PHY_status_MII_Interface_n001118 : X_LUT4
    generic map(
      INIT => X"00E0"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd4,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd3,
      ADR2 => clkslen,
      ADR3 => RESET_IBUF,
      O => mac_control_PHY_status_MII_Interface_CHOICE1541_FROM
    );
  mac_control_PHY_status_MII_Interface_n001124 : X_LUT4
    generic map(
      INIT => X"1100"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_n001124_2,
      ADR1 => mac_control_PHY_status_MII_Interface_n001124_SW0_2,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE1541,
      O => mac_control_PHY_status_MII_Interface_CHOICE1541_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE1541_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE1541_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE1541
    );
  mac_control_PHY_status_MII_Interface_CHOICE1541_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE1541_GROM,
      O => mac_control_PHY_status_MII_Interface_N72822
    );
  rx_input_memio_crccomb_Mxor_n0009_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_datal(3),
      ADR3 => rx_input_memio_crcl(28),
      O => rx_input_memio_crcl_30_FROM
    );
  rx_input_memio_n0048_30_1 : X_LUT4
    generic map(
      INIT => X"F3FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crccomb_Mxor_CO_30_Xo_1_1_2,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crccomb_n0115(0),
      O => rx_input_memio_n0048(30)
    );
  rx_input_memio_crcl_30_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_30_FROM,
      O => rx_input_memio_crccomb_n0115(0)
    );
  rx_input_memio_addrchk_n00301 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd3,
      ADR1 => VCC,
      ADR2 => rx_input_RESET_1,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_n0030_GROM
    );
  rx_input_memio_addrchk_n0030_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_n0030_GROM,
      O => rx_input_memio_addrchk_n0030
    );
  rx_input_memio_addrchk_n00311 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_cs_FFd2,
      ADR2 => VCC,
      ADR3 => rx_input_RESET_1,
      O => rx_input_memio_addrchk_n0031_GROM
    );
  rx_input_memio_addrchk_n0031_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_n0031_GROM,
      O => rx_input_memio_addrchk_n0031
    );
  rx_input_memio_addrchk_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"3320"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd1,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => rx_input_memio_brdy,
      ADR3 => rx_input_memio_addrchk_cs_FFd7,
      O => rx_input_memio_addrchk_cs_FFd7_In
    );
  rx_input_memio_addrchk_n00321 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => rx_input_RESET_1,
      ADR1 => VCC,
      ADR2 => rx_input_memio_addrchk_cs_FFd1,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_cs_FFd7_GROM
    );
  rx_input_memio_addrchk_cs_FFd7_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_cs_FFd7_GROM,
      O => rx_input_memio_addrchk_n0032
    );
  rx_input_memio_addrchk_n00414 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(17),
      ADR1 => rx_input_memio_addrchk_datal(16),
      ADR2 => rx_input_memio_addrchk_datal(18),
      ADR3 => rx_input_memio_addrchk_datal(19),
      O => rx_input_memio_addrchk_CHOICE1424_GROM
    );
  rx_input_memio_addrchk_CHOICE1424_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1424_GROM,
      O => rx_input_memio_addrchk_CHOICE1424
    );
  rx_input_memio_addrchk_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"00D8"
    )
    port map (
      ADR0 => rx_input_memio_brdy,
      ADR1 => rx_input_memio_addrchk_cs_FFd6,
      ADR2 => rx_input_memio_addrchk_cs_FFd5,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_addrchk_cs_FFd5_In
    );
  rx_input_memio_addrchk_n00271 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd6,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_RESET_1,
      O => rx_input_memio_addrchk_cs_FFd5_GROM
    );
  rx_input_memio_addrchk_cs_FFd5_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_cs_FFd5_GROM,
      O => rx_input_memio_addrchk_n0027
    );
  tx_output_addrl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_addrl_11_CEMUXNOT
    );
  rx_input_memio_addrchk_n00281 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_cs_FFd5,
      ADR2 => VCC,
      ADR3 => rx_input_RESET_1,
      O => rx_input_memio_addrchk_n0028_GROM
    );
  rx_input_memio_addrchk_n0028_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_n0028_GROM,
      O => rx_input_memio_addrchk_n0028
    );
  tx_output_addrl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_addrl_13_CEMUXNOT
    );
  rx_input_memio_addrchk_n00354 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(1),
      ADR1 => rx_input_memio_addrchk_datal(2),
      ADR2 => rx_input_memio_addrchk_datal(0),
      ADR3 => rx_input_memio_addrchk_datal(3),
      O => rx_input_memio_addrchk_CHOICE1431_GROM
    );
  rx_input_memio_addrchk_CHOICE1431_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1431_GROM,
      O => rx_input_memio_addrchk_CHOICE1431
    );
  rx_input_memio_addrchk_n00291 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_RESET_1,
      ADR3 => rx_input_memio_addrchk_cs_FFd4,
      O => rx_input_memio_addrchk_n0029_GROM
    );
  rx_input_memio_addrchk_n0029_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_n0029_GROM,
      O => rx_input_memio_addrchk_n0029
    );
  rx_input_fifo_fifo_BU446 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N8,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2473_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2473
    );
  rx_input_fifo_fifo_N2473_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2473_FFX_SET
    );
  rx_input_memio_addrchk_n00419 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(22),
      ADR1 => rx_input_memio_addrchk_datal(23),
      ADR2 => rx_input_memio_addrchk_datal(21),
      ADR3 => rx_input_memio_addrchk_datal(20),
      O => rx_input_memio_addrchk_bcast_3_FROM
    );
  rx_input_memio_addrchk_n004110 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_CHOICE1424,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1427,
      O => rx_input_memio_addrchk_lbcast(3)
    );
  rx_input_memio_addrchk_bcast_3_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_bcast_3_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_3_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_3_FROM,
      O => rx_input_memio_addrchk_CHOICE1427
    );
  tx_output_addrl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_addrl_15_CEMUXNOT
    );
  rx_input_memio_addrchk_n00444 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(26),
      ADR1 => rx_input_memio_addrchk_datal(27),
      ADR2 => rx_input_memio_addrchk_datal(24),
      ADR3 => rx_input_memio_addrchk_datal(25),
      O => rx_input_memio_addrchk_CHOICE1417_GROM
    );
  rx_input_memio_addrchk_CHOICE1417_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1417_GROM,
      O => rx_input_memio_addrchk_CHOICE1417
    );
  rx_input_memio_addrchk_n00509 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(46),
      ADR1 => rx_input_memio_addrchk_datal(44),
      ADR2 => rx_input_memio_addrchk_datal(45),
      ADR3 => rx_input_memio_addrchk_datal(47),
      O => rx_input_memio_addrchk_bcast_0_FROM
    );
  rx_input_memio_addrchk_n005010 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_CHOICE1403,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1406,
      O => rx_input_memio_addrchk_lbcast(0)
    );
  rx_input_memio_addrchk_bcast_0_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_bcast_0_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_0_FROM,
      O => rx_input_memio_addrchk_CHOICE1406
    );
  rx_input_memio_addrchk_n00359 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(7),
      ADR1 => rx_input_memio_addrchk_datal(4),
      ADR2 => rx_input_memio_addrchk_datal(5),
      ADR3 => rx_input_memio_addrchk_datal(6),
      O => rx_input_memio_addrchk_bcast_5_FROM
    );
  rx_input_memio_addrchk_n003510 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_CHOICE1431,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1434,
      O => rx_input_memio_addrchk_lbcast(5)
    );
  rx_input_memio_addrchk_bcast_5_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_bcast_5_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_5_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_5_FROM,
      O => rx_input_memio_addrchk_CHOICE1434
    );
  rx_input_memio_addrchk_n00384 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(11),
      ADR1 => rx_input_memio_addrchk_datal(9),
      ADR2 => rx_input_memio_addrchk_datal(10),
      ADR3 => rx_input_memio_addrchk_datal(8),
      O => rx_input_memio_addrchk_CHOICE1438_GROM
    );
  rx_input_memio_addrchk_CHOICE1438_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1438_GROM,
      O => rx_input_memio_addrchk_CHOICE1438
    );
  rx_input_memio_addrchk_n00449 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(29),
      ADR1 => rx_input_memio_addrchk_datal(28),
      ADR2 => rx_input_memio_addrchk_datal(31),
      ADR3 => rx_input_memio_addrchk_datal(30),
      O => rx_input_memio_addrchk_bcast_2_FROM
    );
  rx_input_memio_addrchk_n004410 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_CHOICE1417,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1420,
      O => rx_input_memio_addrchk_lbcast(2)
    );
  rx_input_memio_addrchk_bcast_2_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_bcast_2_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_2_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_2_FROM,
      O => rx_input_memio_addrchk_CHOICE1420
    );
  rx_input_memio_addrchk_n00474 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(32),
      ADR1 => rx_input_memio_addrchk_datal(35),
      ADR2 => rx_input_memio_addrchk_datal(34),
      ADR3 => rx_input_memio_addrchk_datal(33),
      O => rx_input_memio_addrchk_CHOICE1410_GROM
    );
  rx_input_memio_addrchk_CHOICE1410_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1410_GROM,
      O => rx_input_memio_addrchk_CHOICE1410
    );
  rx_input_memio_addrchk_n00389 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(12),
      ADR1 => rx_input_memio_addrchk_datal(15),
      ADR2 => rx_input_memio_addrchk_datal(14),
      ADR3 => rx_input_memio_addrchk_datal(13),
      O => rx_input_memio_addrchk_bcast_4_FROM
    );
  rx_input_memio_addrchk_n003810 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_CHOICE1438,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1441,
      O => rx_input_memio_addrchk_lbcast(4)
    );
  rx_input_memio_addrchk_bcast_4_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_bcast_4_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_4_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_4_FROM,
      O => rx_input_memio_addrchk_CHOICE1441
    );
  mac_control_PHY_status_MII_Interface_n0014_0_1 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(0),
      O => mac_control_PHY_status_MII_Interface_n0014(0)
    );
  mac_control_PHY_status_MII_Interface_n0004_2_165 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(5),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(4),
      O => mac_control_PHY_status_MII_Interface_statecnt_0_GROM
    );
  mac_control_PHY_status_MII_Interface_statecnt_0_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_statecnt_0_GROM,
      O => mac_control_PHY_status_MII_Interface_n0004_2
    );
  rx_input_memio_addrchk_n00479 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(36),
      ADR1 => rx_input_memio_addrchk_datal(37),
      ADR2 => rx_input_memio_addrchk_datal(38),
      ADR3 => rx_input_memio_addrchk_datal(39),
      O => rx_input_memio_addrchk_bcast_1_FROM
    );
  rx_input_memio_addrchk_n004710 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_CHOICE1410,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1413,
      O => rx_input_memio_addrchk_lbcast(1)
    );
  rx_input_memio_addrchk_bcast_1_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_bcast_1_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_1_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_1_FROM,
      O => rx_input_memio_addrchk_CHOICE1413
    );
  memcontroller_n00051 : X_LUT4
    generic map(
      INIT => X"0404"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => memcontroller_clknum(0),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => tx_output_cs_FFd15_FROM
    );
  tx_output_cs_FFd16_In1 : X_LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      ADR0 => tx_output_n0006,
      ADR1 => memcontroller_clknum(1),
      ADR2 => memcontroller_clknum(0),
      ADR3 => tx_output_cs_FFd17,
      O => tx_output_cs_FFd16_In
    );
  tx_output_cs_FFd15_XUSED : X_BUF
    port map (
      I => tx_output_cs_FFd15_FROM,
      O => memcontroller_n0005
    );
  rx_input_memio_crccomb_Mxor_CO_1_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_datal(0),
      ADR1 => rx_input_memio_crccomb_n0122(0),
      ADR2 => rx_input_memio_crc_0_Q,
      ADR3 => rx_input_memio_crcl(31),
      O => rx_input_memio_crcl_1_FROM
    );
  rx_input_memio_n0048_1_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_1_Q,
      O => rx_input_memio_n0048(1)
    );
  rx_input_memio_crcl_1_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_1_FROM,
      O => rx_input_memio_crc_1_Q
    );
  tx_output_ldata_5_18_SW0 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => tx_output_cs_FFd4,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd5,
      ADR3 => VCC,
      O => tx_output_N81617_FROM
    );
  tx_output_ldata_2_18_SW0 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd5,
      ADR2 => VCC,
      ADR3 => tx_output_cs_FFd4,
      O => tx_output_N81617_GROM
    );
  tx_output_N81617_XUSED : X_BUF
    port map (
      I => tx_output_N81617_FROM,
      O => tx_output_N81617
    );
  tx_output_N81617_YUSED : X_BUF
    port map (
      I => tx_output_N81617_GROM,
      O => tx_output_N81613
    );
  tx_output_crc_loigc_Mxor_n0009_Result1 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => tx_output_data(3),
      ADR1 => VCC,
      ADR2 => tx_output_crcl(28),
      ADR3 => VCC,
      O => tx_output_crcl_30_FROM
    );
  tx_output_n0034_30_1 : X_LUT4
    generic map(
      INIT => X"AFFA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => VCC,
      ADR2 => tx_output_crc_loigc_Mxor_CO_30_Xo_1_1_2,
      ADR3 => tx_output_crc_loigc_n0115(0),
      O => tx_output_n0034(30)
    );
  tx_output_crcl_30_XUSED : X_BUF
    port map (
      I => tx_output_crcl_30_FROM,
      O => tx_output_crc_loigc_n0115(0)
    );
  mac_control_Mmux_n0017_Result_7_30_SW0 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => mac_control_phyaddr(7),
      ADR1 => mac_control_CHOICE2822,
      ADR2 => mac_control_n0103,
      ADR3 => mac_control_CHOICE2825,
      O => mac_control_N81817_FROM
    );
  mac_control_Mmux_n0017_Result_21_47_SW0 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_n0103,
      ADR1 => mac_control_phyaddr(21),
      ADR2 => mac_control_CHOICE2159,
      ADR3 => mac_control_CHOICE2162,
      O => mac_control_N81817_GROM
    );
  mac_control_N81817_XUSED : X_BUF
    port map (
      I => mac_control_N81817_FROM,
      O => mac_control_N81817
    );
  mac_control_N81817_YUSED : X_BUF
    port map (
      I => mac_control_N81817_GROM,
      O => mac_control_N81813
    );
  rx_input_memio_n00491 : X_LUT4
    generic map(
      INIT => X"0022"
    )
    port map (
      ADR0 => rx_input_ce,
      ADR1 => rx_input_invalid,
      ADR2 => VCC,
      ADR3 => rx_input_endf,
      O => rx_input_memio_n0049
    );
  rx_input_memio_n01021 : X_LUT4
    generic map(
      INIT => X"AAAE"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => rx_input_ce,
      ADR2 => rx_input_endf,
      ADR3 => rx_input_invalid,
      O => rx_input_memio_crcen_GROM
    );
  rx_input_memio_crcen_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcen_CEMUXNOT
    );
  rx_input_memio_crcen_YUSED : X_BUF
    port map (
      I => rx_input_memio_crcen_GROM,
      O => rx_input_memio_n0102
    );
  rx_input_memio_cs_Out916_2_166 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd5,
      ADR2 => rx_input_memio_cs_FFd2,
      ADR3 => rx_input_memio_cs_FFd3,
      O => rx_input_memio_cs_Out916_2_FROM
    );
  rx_input_memio_n00301 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd2,
      ADR3 => rx_input_RESET_1,
      O => rx_input_memio_cs_Out916_2_GROM
    );
  rx_input_memio_cs_Out916_2_XUSED : X_BUF
    port map (
      I => rx_input_memio_cs_Out916_2_FROM,
      O => rx_input_memio_cs_Out916_2
    );
  rx_input_memio_cs_Out916_2_YUSED : X_BUF
    port map (
      I => rx_input_memio_cs_Out916_2_GROM,
      O => rx_input_memio_n0030
    );
  rx_input_memio_n00311 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => rx_input_memio_bpen,
      ADR1 => rx_input_RESET_1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_n0031_GROM
    );
  rx_input_memio_n0031_YUSED : X_BUF
    port map (
      I => rx_input_memio_n0031_GROM,
      O => rx_input_memio_n0031
    );
  rx_input_memio_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"FF40"
    )
    port map (
      ADR0 => rx_input_invalid,
      ADR1 => rx_input_endf,
      ADR2 => rx_input_memio_cs_FFd10,
      ADR3 => rx_input_memio_cs_FFd9,
      O => rx_input_memio_cs_FFd8_In
    );
  rx_input_memio_n00321 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => rx_input_endf,
      ADR1 => rx_input_RESET_1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_cs_FFd8_GROM
    );
  rx_input_memio_cs_FFd8_YUSED : X_BUF
    port map (
      I => rx_input_memio_cs_FFd8_GROM,
      O => rx_input_memio_n0032
    );
  rx_input_memio_n00331 : X_LUT4
    generic map(
      INIT => X"000A"
    )
    port map (
      ADR0 => rx_input_memio_men,
      ADR1 => VCC,
      ADR2 => rx_input_RESET_1,
      ADR3 => rx_input_memio_menl,
      O => rx_input_memio_n0033_GROM
    );
  rx_input_memio_n0033_YUSED : X_BUF
    port map (
      I => rx_input_memio_n0033_GROM,
      O => rx_input_memio_n0033
    );
  rx_input_memio_n0048_5_1 : X_LUT4
    generic map(
      INIT => X"FF66"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0056(2),
      ADR1 => rx_input_memio_crccomb_Mxor_CO_5_Xo_1_1_2,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crcrst,
      O => rx_input_memio_n0048(5)
    );
  rx_input_memio_n00341 : X_LUT4
    generic map(
      INIT => X"5544"
    )
    port map (
      ADR0 => rx_input_RESET_1,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crcen,
      O => rx_input_memio_crcl_5_GROM
    );
  rx_input_memio_crcl_5_YUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_5_GROM,
      O => rx_input_memio_n0034
    );
  rx_input_fifo_fifo_BU562 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N5344,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2453_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2453
    );
  rx_input_fifo_fifo_N2453_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2453_FFX_SET
    );
  rx_input_memio_n00441 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd14,
      ADR3 => rx_input_RESET_1,
      O => rx_input_memio_n0044_GROM
    );
  rx_input_memio_n0044_YUSED : X_BUF
    port map (
      I => rx_input_memio_n0044_GROM,
      O => rx_input_memio_n0044
    );
  rx_input_memio_n00461 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd10,
      ADR2 => VCC,
      ADR3 => rx_input_RESET_1,
      O => rx_input_memio_n0046_GROM
    );
  rx_input_memio_n0046_YUSED : X_BUF
    port map (
      I => rx_input_memio_n0046_GROM,
      O => rx_input_memio_n0046
    );
  rx_input_memio_n00471 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_RESET_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd12,
      O => rx_input_memio_n0047_GROM
    );
  rx_input_memio_n0047_YUSED : X_BUF
    port map (
      I => rx_input_memio_n0047_GROM,
      O => rx_input_memio_n0047
    );
  rx_input_memio_n00597 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => rx_input_memio_crcll(3),
      ADR1 => rx_input_memio_crcll(2),
      ADR2 => rx_input_memio_crcll(0),
      ADR3 => rx_input_memio_crcll(1),
      O => rx_input_memio_CHOICE2913_GROM
    );
  rx_input_memio_CHOICE2913_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE2913_GROM,
      O => rx_input_memio_CHOICE2913
    );
  mac_control_Mmux_n0017_Result_31_67 : X_LUT4
    generic map(
      INIT => X"C800"
    )
    port map (
      ADR0 => mac_control_phystat(31),
      ADR1 => mac_control_N52125,
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_addr(1),
      O => mac_control_CHOICE1821_FROM
    );
  mac_control_n0238_SW0 : X_LUT4
    generic map(
      INIT => X"F7FF"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => mac_control_N52268,
      ADR2 => mac_control_addr(1),
      ADR3 => clkslen,
      O => mac_control_CHOICE1821_GROM
    );
  mac_control_CHOICE1821_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1821_FROM,
      O => mac_control_CHOICE1821
    );
  mac_control_CHOICE1821_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1821_GROM,
      O => mac_control_N70611
    );
  rx_input_fifo_fifo_BU315 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N4410,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2486_FFY_RST,
      O => rx_input_fifo_fifo_N2485
    );
  rx_input_fifo_fifo_N2486_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2486_FFY_RST
    );
  mac_control_Mmux_n0017_Result_12_7 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0087,
      ADR1 => mac_control_lmacaddr(44),
      ADR2 => mac_control_n0103,
      ADR3 => mac_control_phyaddr(12),
      O => mac_control_CHOICE2662_FROM
    );
  mac_control_Mmux_n0017_Result_15_30_SW0 : X_LUT4
    generic map(
      INIT => X"FEEE"
    )
    port map (
      ADR0 => mac_control_CHOICE2886,
      ADR1 => mac_control_CHOICE2889,
      ADR2 => mac_control_n0103,
      ADR3 => mac_control_phyaddr(15),
      O => mac_control_CHOICE2662_GROM
    );
  mac_control_CHOICE2662_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2662_FROM,
      O => mac_control_CHOICE2662
    );
  mac_control_CHOICE2662_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2662_GROM,
      O => mac_control_N81757
    );
  mac_control_PHY_status_n00111 : X_LUT4
    generic map(
      INIT => X"3000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => mac_control_PHY_status_cs_FFd4,
      ADR3 => clkslen,
      O => mac_control_PHY_status_n0011_FROM
    );
  mac_control_PHY_status_n0019_2_167 : X_LUT4
    generic map(
      INIT => X"FFF5"
    )
    port map (
      ADR0 => clkslen,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_cs_FFd2,
      ADR3 => mac_control_PHY_status_cs_FFd4,
      O => mac_control_PHY_status_n0011_GROM
    );
  mac_control_PHY_status_n0011_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_n0011_FROM,
      O => mac_control_PHY_status_n0011
    );
  mac_control_PHY_status_n0011_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_n0011_GROM,
      O => mac_control_PHY_status_n0019_2
    );
  tx_output_ldata_7_18_SW0 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => tx_output_cs_FFd4,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_cs_FFd5,
      O => tx_output_N81605_FROM
    );
  tx_output_ldata_4_18_SW0 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd5,
      ADR2 => VCC,
      ADR3 => tx_output_cs_FFd4,
      O => tx_output_N81605_GROM
    );
  tx_output_N81605_XUSED : X_BUF
    port map (
      I => tx_output_N81605_FROM,
      O => tx_output_N81605
    );
  tx_output_N81605_YUSED : X_BUF
    port map (
      I => tx_output_N81605_GROM,
      O => tx_output_N81609
    );
  rx_input_fifo_fifo_BU252 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3936,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N11_FFY_RST,
      O => rx_input_fifo_fifo_N10
    );
  rx_input_fifo_fifo_N11_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N11_FFY_RST
    );
  mac_control_Mmux_n0017_Result_0_107_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_N52111,
      ADR1 => mac_control_N52132,
      ADR2 => mac_control_rxfifowerr_cnt(0),
      ADR3 => mac_control_phyaddr(0),
      O => mac_control_N81753_FROM
    );
  mac_control_Mmux_n0017_Result_0_107 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0085,
      ADR1 => mac_control_N52236,
      ADR2 => mac_control_lmacaddr(0),
      ADR3 => mac_control_N81753,
      O => mac_control_N81753_GROM
    );
  mac_control_N81753_XUSED : X_BUF
    port map (
      I => mac_control_N81753_FROM,
      O => mac_control_N81753
    );
  mac_control_N81753_YUSED : X_BUF
    port map (
      I => mac_control_N81753_GROM,
      O => mac_control_CHOICE2223
    );
  tx_output_bcntl_12_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bcntl_12_CEMUXNOT
    );
  tx_output_bcntl_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_14_FFY_RST
    );
  tx_output_bcntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_51,
      CE => tx_output_bcntl_14_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_14_FFY_RST,
      O => tx_output_bcntl(13)
    );
  tx_output_bcntl_14_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bcntl_14_CEMUXNOT
    );
  tx_output_bcntl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_15_FFY_RST
    );
  tx_output_bcntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_53,
      CE => tx_output_bcntl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_15_FFY_RST,
      O => tx_output_bcntl(15)
    );
  tx_output_bcntl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bcntl_15_CEMUXNOT
    );
  rx_output_bpl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_bpl_11_CEMUXNOT
    );
  rx_output_bpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_13_FFY_RST
    );
  rx_output_bpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(12),
      CE => rx_output_bpl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_13_FFY_RST,
      O => rx_output_bpl(12)
    );
  rx_output_bpl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_bpl_13_CEMUXNOT
    );
  rx_output_bpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_15_FFY_RST
    );
  rx_output_bpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(14),
      CE => rx_output_bpl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_15_FFY_RST,
      O => rx_output_bpl(14)
    );
  rx_output_bpl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_bpl_15_CEMUXNOT
    );
  rx_output_fifo_N1546_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1546_FFY_RST
    );
  rx_output_fifo_BU133 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2499,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1546_FFY_RST,
      O => rx_output_fifo_N1547
    );
  rx_output_fifo_BU132 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N11,
      ADR3 => rx_output_fifo_N10,
      O => rx_output_fifo_N2499
    );
  rx_output_fifo_N1610_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1610_FFY_RST
    );
  rx_output_fifo_BU294 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3427,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1610_FFY_RST,
      O => rx_output_fifo_N1611
    );
  rx_output_fifo_BU293 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N2,
      ADR3 => rx_output_fifo_N3,
      O => rx_output_fifo_N3427
    );
  rx_output_fifo_N1563_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1563_FFY_SET
    );
  rx_output_fifo_BU320 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1546,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1563_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1562
    );
  rx_input_fifo_fifo_BU308 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N4370,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2486_FFX_RST,
      O => rx_input_fifo_fifo_N2486
    );
  rx_input_fifo_fifo_N2486_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2486_FFX_RST
    );
  rx_output_fifo_N1567_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1567_FFY_RST
    );
  rx_output_fifo_BU312 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1550,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1567_FFY_RST,
      O => rx_output_fifo_N1566
    );
  rx_output_fifo_N1627_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1627_FFY_SET
    );
  rx_output_fifo_BU170 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1610,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1627_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1626
    );
  rx_output_fifo_BU191 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_ceinll,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_full_0,
      O => rx_output_fifo_N19_FROM
    );
  rx_output_fifo_BU323 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_ceinll,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_full_0,
      O => rx_output_fifo_N19_GROM
    );
  rx_output_fifo_N19_XUSED : X_BUF
    port map (
      I => rx_output_fifo_N19_FROM,
      O => rx_output_fifo_N19
    );
  rx_output_fifo_N19_YUSED : X_BUF
    port map (
      I => rx_output_fifo_N19_GROM,
      O => rx_output_fifo_N3617
    );
  rx_output_fifo_N1565_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1565_FFY_RST
    );
  rx_output_fifo_BU316 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1548,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1565_FFY_RST,
      O => rx_output_fifo_N1564
    );
  rx_output_fifo_N1629_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1629_FFY_RST
    );
  rx_output_fifo_BU164 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1612,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1629_FFY_RST,
      O => rx_output_fifo_N1628
    );
  rx_output_fifo_N1633_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1633_FFY_RST
    );
  rx_output_fifo_BU149 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1616,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1633_FFY_RST,
      O => rx_output_fifo_N1632
    );
  q2_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_21_FFY_RST
    );
  memcontroller_Q2_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(20),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_21_FFY_RST,
      O => q2(20)
    );
  q2_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_13_FFY_RST
    );
  memcontroller_Q2_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(12),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_13_FFY_RST,
      O => q2(12)
    );
  rx_output_fifo_N1631_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1631_FFY_RST
    );
  rx_output_fifo_BU158 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1614,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1631_FFY_RST,
      O => rx_output_fifo_N1630
    );
  rx_output_fifo_N1573_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1573_FFY_RST
    );
  rx_output_fifo_BU343 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1564,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1573_FFY_RST,
      O => rx_output_fifo_N1572
    );
  q2_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_31_FFY_RST
    );
  memcontroller_Q2_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(30),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_31_FFY_RST,
      O => q2(30)
    );
  q2_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_15_FFY_RST
    );
  memcontroller_Q2_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(14),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_15_FFY_RST,
      O => q2(14)
    );
  rx_output_fifo_N1577_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1577_FFY_SET
    );
  rx_output_fifo_BU328 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1568,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1577_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1576
    );
  mac_control_phystat_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_11_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(10),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_11_FFY_RST,
      O => mac_control_phystat(10)
    );
  rx_output_fifo_N1575_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1575_FFY_RST
    );
  rx_output_fifo_BU337 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1566,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1575_FFY_RST,
      O => rx_output_fifo_N1574
    );
  rx_output_fifo_BU185 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_ceinll,
      ADR3 => rx_output_fifo_full_0,
      O => rx_output_fifo_N1517_GROM
    );
  rx_output_fifo_N1517_YUSED : X_BUF
    port map (
      I => rx_output_fifo_N1517_GROM,
      O => rx_output_fifo_N1517
    );
  q2_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_17_FFY_RST
    );
  memcontroller_Q2_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(16),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_17_FFY_RST,
      O => q2(16)
    );
  rx_output_cs_FFd18_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd18_FFY_RST
    );
  rx_output_cs_FFd18_168 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd18_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd18_FFY_RST,
      O => rx_output_cs_FFd18
    );
  memcontroller_n00101 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => memcontroller_clknum(0),
      O => rx_output_cs_FFd18_FROM
    );
  rx_output_cs_FFd18_In_169 : X_LUT4
    generic map(
      INIT => X"D5F5"
    )
    port map (
      ADR0 => rx_output_cs_FFd18_In_2,
      ADR1 => rx_output_n0017,
      ADR2 => rx_output_cs_FFd18,
      ADR3 => clken3,
      O => rx_output_cs_FFd18_In
    );
  rx_output_cs_FFd18_XUSED : X_BUF
    port map (
      I => rx_output_cs_FFd18_FROM,
      O => clken3
    );
  rx_output_fifo_N1609_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1609_FFY_SET
    );
  rx_output_fifo_BU362 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N8,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1609_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1608
    );
  mac_control_phystat_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_21_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(4),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_21_FFY_RST,
      O => mac_control_phystat(20)
    );
  mac_control_phystat_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_13_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(12),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_13_FFY_RST,
      O => mac_control_phystat(12)
    );
  q2_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_27_FFY_RST
    );
  memcontroller_Q2_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(26),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_27_FFY_RST,
      O => q2(26)
    );
  rx_input_fifo_fifo_BU402 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2425,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N2436_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2435
    );
  rx_input_fifo_fifo_N2436_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2436_FFY_SET
    );
  q2_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_19_FFY_RST
    );
  memcontroller_Q2_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(18),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_19_FFY_RST,
      O => q2(18)
    );
  q3_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_11_FFY_RST
    );
  memcontroller_Q3_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(10),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_11_FFY_RST,
      O => q3(10)
    );
  rx_output_fifo_N1585_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1585_FFY_RST
    );
  rx_output_fifo_BU380 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1552,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1585_FFY_RST,
      O => rx_output_fifo_N1584
    );
  mac_control_phystat_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_23_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(6),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_23_FFY_RST,
      O => mac_control_phystat(22)
    );
  rx_input_fifo_fifo_BU246 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3935,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N11_FFX_RST,
      O => rx_input_fifo_fifo_N11
    );
  rx_input_fifo_fifo_N11_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N11_FFX_RST
    );
  mac_control_phystat_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_31_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(14),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_31_FFY_RST,
      O => mac_control_phystat(30)
    );
  rx_output_fifo_N1571_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1571_FFY_SET
    );
  rx_output_fifo_BU349 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1562,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1571_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1570
    );
  rx_input_fifo_fifo_BU376 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2406,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N2425_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2426
    );
  rx_input_fifo_fifo_N2425_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2425_FFY_SET
    );
  q2_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_29_FFY_RST
    );
  memcontroller_Q2_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(28),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_29_FFY_RST,
      O => q2(28)
    );
  q3_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_21_FFY_RST
    );
  memcontroller_Q3_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(20),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_21_FFY_RST,
      O => q3(20)
    );
  q3_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_13_FFY_RST
    );
  memcontroller_Q3_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(12),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_13_FFY_RST,
      O => q3(12)
    );
  rx_output_fifo_N1586_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1586_FFY_SET
    );
  rx_output_fifo_BU468 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3974,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1586_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1587
    );
  rx_output_fifo_BU410 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N1578,
      ADR2 => rx_output_fifo_N1579,
      ADR3 => VCC,
      O => rx_output_fifo_N3974
    );
  rx_output_fifo_N1591_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1591_FFX_SET
    );
  rx_output_fifo_BU460 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3970,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1591_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1591
    );
  rx_output_fifo_BU434 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => rx_output_fifo_N3959,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N1583,
      ADR3 => rx_output_fifo_N1582,
      O => rx_output_fifo_N3970
    );
  rx_output_fifo_BU446 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_output_fifo_N1583,
      ADR1 => rx_output_fifo_N1584,
      ADR2 => rx_output_fifo_N1585,
      ADR3 => rx_output_fifo_N1582,
      O => rx_output_fifo_N1591_GROM
    );
  rx_output_fifo_N1591_YUSED : X_BUF
    port map (
      I => rx_output_fifo_N1591_GROM,
      O => rx_output_fifo_N3958
    );
  rx_output_fifo_N1603_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1603_FFY_SET
    );
  rx_output_fifo_BU374 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N2,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1603_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1602
    );
  rx_output_fifo_N1607_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1607_FFY_SET
    );
  rx_output_fifo_BU366 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N6,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1607_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1606
    );
  mac_control_phystat_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_25_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(8),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_25_FFY_RST,
      O => mac_control_phystat(24)
    );
  mac_control_phystat_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_17_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(0),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_17_FFY_RST,
      O => mac_control_phystat(16)
    );
  q3_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_31_FFY_RST
    );
  memcontroller_Q3_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(30),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_31_FFY_RST,
      O => q3(30)
    );
  q3_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_23_FFY_RST
    );
  memcontroller_Q3_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(22),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_23_FFY_RST,
      O => q3(22)
    );
  q3_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_15_FFY_RST
    );
  memcontroller_Q3_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(14),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_15_FFY_RST,
      O => q3(14)
    );
  rx_output_fifo_N1579_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1579_FFY_SET
    );
  rx_output_fifo_BU392 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1546,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1579_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1578
    );
  mac_control_phystat_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_19_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(2),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_19_FFY_RST,
      O => mac_control_phystat(18)
    );
  q3_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_25_FFY_RST
    );
  memcontroller_Q3_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(24),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_25_FFY_RST,
      O => q3(24)
    );
  q3_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_17_FFY_RST
    );
  memcontroller_Q3_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(16),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_17_FFY_RST,
      O => q3(16)
    );
  memcontroller_n00111 : X_LUT4
    generic map(
      INIT => X"F00F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(0),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_wen
    );
  memcontroller_n00061 : X_LUT4
    generic map(
      INIT => X"0500"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(0),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_oe_GROM
    );
  memcontroller_oe_YUSED : X_BUF
    port map (
      I => memcontroller_oe_GROM,
      O => memcontroller_n0006
    );
  rx_input_fifo_fifo_BU378 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2405,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2425_FFX_RST,
      O => rx_input_fifo_fifo_N2425
    );
  rx_input_fifo_fifo_N2425_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2425_FFX_RST
    );
  q3_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_27_FFY_RST
    );
  memcontroller_Q3_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(26),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_27_FFY_RST,
      O => q3(26)
    );
  q3_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_19_FFY_RST
    );
  memcontroller_Q3_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(18),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_19_FFY_RST,
      O => q3(18)
    );
  rx_output_fifo_N1581_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1581_FFY_RST
    );
  rx_output_fifo_BU388 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1548,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1581_FFY_RST,
      O => rx_output_fifo_N1580
    );
  rx_input_fifo_fifo_BU462 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2406,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2445_FFY_RST,
      O => rx_input_fifo_fifo_N2446
    );
  rx_input_fifo_fifo_N2445_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2445_FFY_RST
    );
  q3_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_29_FFY_RST
    );
  memcontroller_Q3_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(28),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_29_FFY_RST,
      O => q3(28)
    );
  tx_output_cs_FFd17_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => tx_output_cs_FFd17_FFY_SET
    );
  tx_output_cs_FFd17_170 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => tx_output_cs_FFd17_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => tx_output_cs_FFd17_FFY_SET,
      RST => GND,
      O => tx_output_cs_FFd17
    );
  memcontroller_n00091 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => memcontroller_clknum(0),
      O => tx_output_cs_FFd17_FROM
    );
  tx_output_cs_FFd17_In1 : X_LUT4
    generic map(
      INIT => X"EAEE"
    )
    port map (
      ADR0 => tx_output_cs_FFd1,
      ADR1 => tx_output_cs_FFd17,
      ADR2 => tx_output_n0006,
      ADR3 => clken2,
      O => tx_output_cs_FFd17_In
    );
  tx_output_cs_FFd17_XUSED : X_BUF
    port map (
      I => tx_output_cs_FFd17_FROM,
      O => clken2
    );
  rx_output_ceinll_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_ceinll_CEMUXNOT
    );
  mac_control_PHY_status_MII_Interface_n00131 : X_LUT4
    generic map(
      INIT => X"F0E0"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd4,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd3,
      ADR2 => mac_control_PHY_status_MII_Interface_N37245,
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      O => mac_control_PHY_status_MII_Interface_n0013_FROM
    );
  mac_control_PHY_status_MII_Interface_cs_FFd3_In_SW0 : X_LUT4
    generic map(
      INIT => X"55FF"
    )
    port map (
      ADR0 => MDC_OBUF,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd4,
      O => mac_control_PHY_status_MII_Interface_n0013_GROM
    );
  mac_control_PHY_status_MII_Interface_n0013_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0013_FROM,
      O => mac_control_PHY_status_MII_Interface_n0013
    );
  mac_control_PHY_status_MII_Interface_n0013_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0013_GROM,
      O => mac_control_PHY_status_MII_Interface_N69539
    );
  tx_output_crc_loigc_Mxor_CO_10_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(2),
      ADR1 => tx_output_crc_loigc_Mxor_CO_7_Xo(1),
      ADR2 => tx_output_crc_loigc_n0118(1),
      ADR3 => tx_output_crc_loigc_n0118(0),
      O => tx_output_crcl_10_FROM
    );
  tx_output_n0034_10_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16,
      ADR2 => VCC,
      ADR3 => tx_output_crc_10_Q,
      O => tx_output_n0034(10)
    );
  tx_output_crcl_10_XUSED : X_BUF
    port map (
      I => tx_output_crcl_10_FROM,
      O => tx_output_crc_10_Q
    );
  mac_control_PHY_status_MII_Interface_n00161 : X_LUT4
    generic map(
      INIT => X"00C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd2,
      ADR2 => clkslen,
      ADR3 => RESET_IBUF,
      O => mac_control_PHY_status_MII_Interface_n0016_GROM
    );
  mac_control_PHY_status_MII_Interface_n0016_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0016_GROM,
      O => mac_control_PHY_status_MII_Interface_n0016
    );
  tx_output_addrl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_addrl_1_CEMUXNOT
    );
  tx_output_addrl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_3_FFY_RST
    );
  tx_output_addrl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(2),
      CE => tx_output_addrl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_3_FFY_RST,
      O => tx_output_addrl(2)
    );
  tx_output_addrl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_addrl_3_CEMUXNOT
    );
  tx_output_addrl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_5_FFY_RST
    );
  tx_output_addrl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(4),
      CE => tx_output_addrl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_5_FFY_RST,
      O => tx_output_addrl(4)
    );
  tx_output_addrl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_addrl_5_CEMUXNOT
    );
  tx_output_addrl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_7_FFY_RST
    );
  tx_output_addrl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(6),
      CE => tx_output_addrl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_7_FFY_RST,
      O => tx_output_addrl(6)
    );
  tx_output_addrl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_addrl_7_CEMUXNOT
    );
  rx_output_len_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_11_FFY_RST
    );
  rx_output_len_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(10),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_11_FFY_RST,
      O => rx_output_len(10)
    );
  rx_input_fifo_fifo_BU399 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2426,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N2436_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2436
    );
  rx_input_fifo_fifo_N2436_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2436_FFX_SET
    );
  rx_output_mdl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_11_FFY_RST
    );
  rx_output_mdl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(10),
      CE => rx_output_mdl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_11_FFY_RST,
      O => rx_output_mdl(10)
    );
  rx_output_mdl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_11_CEMUXNOT
    );
  tx_output_addrl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_addrl_9_CEMUXNOT
    );
  rx_output_len_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_13_FFY_RST
    );
  rx_output_len_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(12),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_13_FFY_RST,
      O => rx_output_len(12)
    );
  rx_output_mdl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_21_FFY_RST
    );
  rx_output_mdl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(20),
      CE => rx_output_mdl_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_21_FFY_RST,
      O => rx_output_mdl(20)
    );
  rx_output_mdl_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_21_CEMUXNOT
    );
  rx_output_mdl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_13_FFY_RST
    );
  rx_output_mdl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(12),
      CE => rx_output_mdl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_13_FFY_RST,
      O => rx_output_mdl(12)
    );
  rx_output_mdl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_13_CEMUXNOT
    );
  rx_output_mdl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_31_FFY_RST
    );
  rx_output_mdl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(30),
      CE => rx_output_mdl_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_31_FFY_RST,
      O => rx_output_mdl(30)
    );
  rx_output_mdl_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_31_CEMUXNOT
    );
  rx_output_mdl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_23_FFY_RST
    );
  rx_output_mdl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(22),
      CE => rx_output_mdl_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_23_FFY_RST,
      O => rx_output_mdl(22)
    );
  rx_output_mdl_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_23_CEMUXNOT
    );
  rx_output_mdl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_15_FFY_RST
    );
  rx_output_mdl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(14),
      CE => rx_output_mdl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_15_FFY_RST,
      O => rx_output_mdl(14)
    );
  rx_output_mdl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_15_CEMUXNOT
    );
  rx_input_fifo_fifo_BU464 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2405,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2445_FFX_RST,
      O => rx_input_fifo_fifo_N2445
    );
  rx_input_fifo_fifo_N2445_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2445_FFX_RST
    );
  rx_output_mdl_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_25_CEMUXNOT
    );
  rx_output_mdl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_17_FFY_RST
    );
  rx_output_mdl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(16),
      CE => rx_output_mdl_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_17_FFY_RST,
      O => rx_output_mdl(16)
    );
  rx_output_mdl_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_17_CEMUXNOT
    );
  mac_control_Mmux_n0017_Result_13_7 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phyaddr(13),
      ADR1 => mac_control_lmacaddr(45),
      ADR2 => mac_control_n0087,
      ADR3 => mac_control_n0103,
      O => mac_control_CHOICE2693_FROM
    );
  mac_control_Mmux_n0017_Result_16_47_SW0 : X_LUT4
    generic map(
      INIT => X"FEFC"
    )
    port map (
      ADR0 => mac_control_phyaddr(16),
      ADR1 => mac_control_CHOICE2111,
      ADR2 => mac_control_CHOICE2114,
      ADR3 => mac_control_n0103,
      O => mac_control_CHOICE2693_GROM
    );
  mac_control_CHOICE2693_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2693_FROM,
      O => mac_control_CHOICE2693
    );
  mac_control_CHOICE2693_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2693_GROM,
      O => mac_control_N81793
    );
  rx_output_mdl_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_27_CEMUXNOT
    );
  rx_output_mdl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_19_FFY_RST
    );
  rx_output_mdl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(18),
      CE => rx_output_mdl_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_19_FFY_RST,
      O => rx_output_mdl(18)
    );
  rx_output_mdl_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_19_CEMUXNOT
    );
  rx_output_mdl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_29_FFY_RST
    );
  rx_output_mdl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(28),
      CE => rx_output_mdl_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_29_FFY_RST,
      O => rx_output_mdl(28)
    );
  rx_output_mdl_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_29_CEMUXNOT
    );
  rx_output_lmasell_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lmasell_FFY_RST
    );
  rx_output_lmasell_171 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd7,
      CE => rx_output_lmasell_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lmasell_FFY_RST,
      O => rx_output_lmasell
    );
  rx_output_lmasell_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lmasell_CEMUXNOT
    );
  tx_output_n000774 : X_LUT4
    generic map(
      INIT => X"0010"
    )
    port map (
      ADR0 => tx_output_bcnt_39,
      ADR1 => tx_output_bcnt_40,
      ADR2 => tx_output_bcnt_38,
      ADR3 => tx_output_N81677,
      O => tx_output_cs_FFd3_FROM
    );
  tx_output_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd5,
      ADR2 => VCC,
      ADR3 => tx_output_N73488,
      O => tx_output_cs_FFd4_In
    );
  tx_output_cs_FFd3_XUSED : X_BUF
    port map (
      I => tx_output_cs_FFd3_FROM,
      O => tx_output_N73488
    );
  tx_input_enable_LOGIC_ONE_172 : X_ONE
    port map (
      O => tx_input_enable_LOGIC_ONE
    );
  rx_input_memio_crccomb_Mxor_CO_3_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0118(1),
      ADR1 => rx_input_memio_crccomb_n0122(0),
      ADR2 => rx_input_memio_crccomb_n0124(1),
      ADR3 => rx_input_memio_crccomb_n0124(0),
      O => rx_input_memio_crcl_3_FROM
    );
  rx_input_memio_n0048_3_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_3_Q,
      O => rx_input_memio_n0048(3)
    );
  rx_input_memio_crcl_3_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_3_FROM,
      O => rx_input_memio_crc_3_Q
    );
  mac_control_Mmux_n0017_Result_6_107_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(6),
      ADR1 => mac_control_phyaddr(6),
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_N52132,
      O => mac_control_N82125_FROM
    );
  mac_control_Mmux_n0017_Result_1_107_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_N52111,
      ADR1 => mac_control_N52132,
      ADR2 => mac_control_rxfifowerr_cnt(1),
      ADR3 => mac_control_phyaddr(1),
      O => mac_control_N82125_GROM
    );
  mac_control_N82125_XUSED : X_BUF
    port map (
      I => mac_control_N82125_FROM,
      O => mac_control_N82125
    );
  mac_control_N82125_YUSED : X_BUF
    port map (
      I => mac_control_N82125_GROM,
      O => mac_control_N82137
    );
  txfifofull_LOGIC_ONE_173 : X_ONE
    port map (
      O => txfifofull_LOGIC_ONE
    );
  rx_input_fifo_fifo_BU442 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N10,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2475_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2475
    );
  rx_input_fifo_fifo_N2475_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2475_FFX_SET
    );
  mac_control_Mmux_n0017_Result_9_7 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_lmacaddr(41),
      ADR1 => mac_control_n0103,
      ADR2 => mac_control_phyaddr(9),
      ADR3 => mac_control_n0087,
      O => mac_control_CHOICE2631_FROM
    );
  mac_control_Mmux_n0017_Result_17_47_SW0 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_CHOICE2135,
      ADR1 => mac_control_n0103,
      ADR2 => mac_control_phyaddr(17),
      ADR3 => mac_control_CHOICE2138,
      O => mac_control_CHOICE2631_GROM
    );
  mac_control_CHOICE2631_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2631_FROM,
      O => mac_control_CHOICE2631
    );
  mac_control_CHOICE2631_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2631_GROM,
      O => mac_control_N81749
    );
  rx_input_fifo_fifo_BU556 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N5341,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2455_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2456
    );
  rx_input_fifo_fifo_N2455_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2455_FFY_SET
    );
  tx_output_bcntl_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bcntl_2_CEMUXNOT
    );
  tx_output_bcntl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_4_FFY_RST
    );
  tx_output_bcntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_41,
      CE => tx_output_bcntl_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_4_FFY_RST,
      O => tx_output_bcntl(3)
    );
  tx_output_bcntl_4_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bcntl_4_CEMUXNOT
    );
  tx_output_bcntl_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_6_FFY_RST
    );
  tx_output_bcntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_43,
      CE => tx_output_bcntl_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_6_FFY_RST,
      O => tx_output_bcntl(5)
    );
  tx_output_bcntl_6_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bcntl_6_CEMUXNOT
    );
  rx_output_bpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_1_FFY_RST
    );
  rx_output_bpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(0),
      CE => rx_output_bpl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_1_FFY_RST,
      O => rx_output_bpl(0)
    );
  rx_output_bpl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_bpl_1_CEMUXNOT
    );
  tx_output_bcntl_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_8_FFY_RST
    );
  tx_output_bcntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_45,
      CE => tx_output_bcntl_8_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_8_FFY_RST,
      O => tx_output_bcntl(7)
    );
  tx_output_bcntl_8_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bcntl_8_CEMUXNOT
    );
  rx_output_bpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_3_FFY_RST
    );
  rx_output_bpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(2),
      CE => rx_output_bpl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_3_FFY_RST,
      O => rx_output_bpl(2)
    );
  rx_output_bpl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_bpl_3_CEMUXNOT
    );
  tx_output_datal_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_1_FFY_RST
    );
  tx_output_datal_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(0),
      CE => tx_output_datal_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_1_FFY_RST,
      O => tx_output_datal(0)
    );
  tx_output_datal_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_datal_1_CEMUXNOT
    );
  tx_output_bcntl_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_10_FFY_RST
    );
  tx_output_bcntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_47,
      CE => tx_output_bcntl_10_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_10_FFY_RST,
      O => tx_output_bcntl(9)
    );
  tx_output_bcntl_10_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bcntl_10_CEMUXNOT
    );
  rx_output_bpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_5_FFY_RST
    );
  rx_output_bpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(4),
      CE => rx_output_bpl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_5_FFY_RST,
      O => rx_output_bpl(4)
    );
  rx_output_bpl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_bpl_5_CEMUXNOT
    );
  tx_output_datal_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_3_FFY_RST
    );
  tx_output_datal_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(2),
      CE => tx_output_datal_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_3_FFY_RST,
      O => tx_output_datal(2)
    );
  tx_output_datal_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_datal_3_CEMUXNOT
    );
  rx_output_bpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_7_FFY_RST
    );
  rx_output_bpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(6),
      CE => rx_output_bpl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_7_FFY_RST,
      O => rx_output_bpl(6)
    );
  rx_output_bpl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_bpl_7_CEMUXNOT
    );
  tx_output_datal_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_5_FFY_RST
    );
  tx_output_datal_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(4),
      CE => tx_output_datal_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_5_FFY_RST,
      O => tx_output_datal(4)
    );
  tx_output_datal_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_datal_5_CEMUXNOT
    );
  tx_output_crcl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_11_FFY_RST
    );
  tx_output_crcl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(11),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_11_FFY_RST,
      O => tx_output_crcl(11)
    );
  tx_output_crc_loigc_Mxor_CO_11_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_Mxor_CO_23_Xo(0),
      ADR1 => tx_output_crc_loigc_n0124(1),
      ADR2 => tx_output_crc_loigc_n0115(0),
      ADR3 => tx_output_crcl(3),
      O => tx_output_crcl_11_FROM
    );
  tx_output_n0034_11_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_crc_11_Q,
      ADR3 => tx_output_cs_FFd16,
      O => tx_output_n0034(11)
    );
  tx_output_crcl_11_XUSED : X_BUF
    port map (
      I => tx_output_crcl_11_FROM,
      O => tx_output_crc_11_Q
    );
  rx_output_bpl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_bpl_9_CEMUXNOT
    );
  tx_output_datal_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_7_FFY_RST
    );
  tx_output_datal_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(6),
      CE => tx_output_datal_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_7_FFY_RST,
      O => tx_output_datal(6)
    );
  tx_output_datal_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_datal_7_CEMUXNOT
    );
  mac_control_dout_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_1_FFY_RST
    );
  mac_control_dout_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N76543,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_1_FFY_RST,
      O => mac_control_dout(1)
    );
  mac_control_Mmux_n0017_Result_1_149_SW0 : X_LUT4
    generic map(
      INIT => X"0105"
    )
    port map (
      ADR0 => mac_control_CHOICE2259,
      ADR1 => mac_control_lmacaddr(1),
      ADR2 => mac_control_CHOICE2242,
      ADR3 => mac_control_n0085,
      O => mac_control_dout_1_FROM
    );
  mac_control_Mmux_n0017_Result_1_149 : X_LUT4
    generic map(
      INIT => X"444E"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_dout(0),
      ADR2 => mac_control_addr(5),
      ADR3 => mac_control_N81657,
      O => mac_control_N76543
    );
  mac_control_dout_1_XUSED : X_BUF
    port map (
      I => mac_control_dout_1_FROM,
      O => mac_control_N81657
    );
  tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_2_174 : X_LUT4
    generic map(
      INIT => X"C33C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_crc_loigc_n0104(0),
      ADR2 => tx_output_crcl(4),
      ADR3 => tx_output_crc_loigc_n0115(0),
      O => tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_2_GROM
    );
  tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_2_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_2_GROM,
      O => tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_2
    );
  rx_output_mdl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_1_FFY_RST
    );
  rx_output_mdl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(0),
      CE => rx_output_mdl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_1_FFY_RST,
      O => rx_output_mdl(0)
    );
  rx_output_mdl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_1_CEMUXNOT
    );
  rx_output_mdl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_3_FFY_RST
    );
  rx_output_mdl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(2),
      CE => rx_output_mdl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_3_FFY_RST,
      O => rx_output_mdl(2)
    );
  rx_output_mdl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_3_CEMUXNOT
    );
  rx_output_mdl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_5_FFY_RST
    );
  rx_output_mdl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(4),
      CE => rx_output_mdl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_5_FFY_RST,
      O => rx_output_mdl(4)
    );
  rx_output_mdl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_5_CEMUXNOT
    );
  rx_output_mdl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_7_FFY_RST
    );
  rx_output_mdl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(6),
      CE => rx_output_mdl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_7_FFY_RST,
      O => rx_output_mdl(6)
    );
  rx_output_mdl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_7_CEMUXNOT
    );
  rx_input_fifo_fifo_BU558 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N5342,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2455_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2455
    );
  rx_input_fifo_fifo_N2455_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2455_FFX_SET
    );
  rx_output_mdl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_9_FFY_RST
    );
  rx_output_mdl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(8),
      CE => rx_output_mdl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_9_FFY_RST,
      O => rx_output_mdl(8)
    );
  rx_output_mdl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_9_CEMUXNOT
    );
  tx_output_ltxd_0_SW0 : X_LUT4
    generic map(
      INIT => X"EEAA"
    )
    port map (
      ADR0 => tx_output_outselll(1),
      ADR1 => tx_output_datal(0),
      ADR2 => VCC,
      ADR3 => tx_output_outselll(0),
      O => tx_output_N70584_FROM
    );
  tx_output_ltxd_0_Q : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => tx_output_outselll(3),
      ADR1 => tx_output_outselll(2),
      ADR2 => tx_output_ncrcbytel(7),
      ADR3 => tx_output_N70584,
      O => tx_output_N70584_GROM
    );
  tx_output_N70584_XUSED : X_BUF
    port map (
      I => tx_output_N70584_FROM,
      O => tx_output_N70584
    );
  tx_output_N70584_YUSED : X_BUF
    port map (
      I => tx_output_N70584_GROM,
      O => tx_output_ltxd(0)
    );
  rx_input_GMII_ro_LOGIC_ONE_175 : X_ONE
    port map (
      O => rx_input_GMII_ro_LOGIC_ONE
    );
  mac_control_n00561_2_176 : X_LUT4
    generic map(
      INIT => X"8080"
    )
    port map (
      ADR0 => mac_control_addr(7),
      ADR1 => mac_control_N52236,
      ADR2 => mac_control_N52132,
      ADR3 => VCC,
      O => mac_control_n00561_2_FROM
    );
  mac_control_Mmux_n0017_Result_2_107_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_phyaddr(2),
      ADR1 => mac_control_rxfifowerr_cnt(2),
      ADR2 => mac_control_N52132,
      ADR3 => mac_control_N52111,
      O => mac_control_n00561_2_GROM
    );
  mac_control_n00561_2_XUSED : X_BUF
    port map (
      I => mac_control_n00561_2_FROM,
      O => mac_control_n00561_2
    );
  mac_control_n00561_2_YUSED : X_BUF
    port map (
      I => mac_control_n00561_2_GROM,
      O => mac_control_N82113
    );
  tx_output_outselll_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_outselll_1_CEMUXNOT
    );
  tx_output_outselll_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_outselll_3_CEMUXNOT
    );
  tx_output_ltxd_2_SW0 : X_LUT4
    generic map(
      INIT => X"EEAA"
    )
    port map (
      ADR0 => tx_output_outselll(1),
      ADR1 => tx_output_outselll(0),
      ADR2 => VCC,
      ADR3 => tx_output_datal(2),
      O => tx_output_N70557_FROM
    );
  tx_output_ltxd_2_Q : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => tx_output_outselll(2),
      ADR1 => tx_output_ncrcbytel(5),
      ADR2 => tx_output_outselll(3),
      ADR3 => tx_output_N70557,
      O => tx_output_N70557_GROM
    );
  tx_output_N70557_XUSED : X_BUF
    port map (
      I => tx_output_N70557_FROM,
      O => tx_output_N70557
    );
  tx_output_N70557_YUSED : X_BUF
    port map (
      I => tx_output_N70557_GROM,
      O => tx_output_ltxd(2)
    );
  tx_output_ltxd_4_SW0 : X_LUT4
    generic map(
      INIT => X"FAAA"
    )
    port map (
      ADR0 => tx_output_outselll(1),
      ADR1 => VCC,
      ADR2 => tx_output_datal(4),
      ADR3 => tx_output_outselll(0),
      O => tx_output_N70530_FROM
    );
  tx_output_ltxd_4_Q : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => tx_output_outselll(3),
      ADR1 => tx_output_outselll(2),
      ADR2 => tx_output_ncrcbytel(3),
      ADR3 => tx_output_N70530,
      O => tx_output_N70530_GROM
    );
  tx_output_N70530_XUSED : X_BUF
    port map (
      I => tx_output_N70530_FROM,
      O => tx_output_N70530
    );
  tx_output_N70530_YUSED : X_BUF
    port map (
      I => tx_output_N70530_GROM,
      O => tx_output_ltxd(4)
    );
  rx_input_fifo_fifo_BU42 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2724,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_dout_9_FFY_RST,
      O => rx_input_fifo_dout(9)
    );
  rx_input_fifo_dout_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_dout_9_FFY_RST
    );
  tx_output_ldata_0_18 : X_LUT4
    generic map(
      INIT => X"E4A0"
    )
    port map (
      ADR0 => tx_output_cs_FFd6,
      ADR1 => q2(8),
      ADR2 => q2(0),
      ADR3 => tx_output_N81625,
      O => tx_output_data_0_FROM
    );
  tx_output_ldata_0_25 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_CHOICE1289,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1297,
      O => tx_output_ldata(0)
    );
  tx_output_data_0_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_data_0_CEMUXNOT
    );
  tx_output_data_0_XUSED : X_BUF
    port map (
      I => tx_output_data_0_FROM,
      O => tx_output_CHOICE1297
    );
  tx_output_ldata_1_18 : X_LUT4
    generic map(
      INIT => X"CAC0"
    )
    port map (
      ADR0 => tx_output_N81625,
      ADR1 => q2(1),
      ADR2 => tx_output_cs_FFd6,
      ADR3 => q2(9),
      O => tx_output_data_1_FROM
    );
  tx_output_ldata_1_25 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_CHOICE1277,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1285,
      O => tx_output_ldata(1)
    );
  tx_output_data_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_data_1_CEMUXNOT
    );
  tx_output_data_1_XUSED : X_BUF
    port map (
      I => tx_output_data_1_FROM,
      O => tx_output_CHOICE1285
    );
  tx_output_crc_loigc_Mxor_CO_12_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(2),
      ADR1 => tx_output_crc_loigc_Mxor_CO_23_Xo(0),
      ADR2 => tx_output_crcl(29),
      ADR3 => tx_output_crc_loigc_n0118(1),
      O => tx_output_crcl_12_FROM
    );
  tx_output_n0034_12_1 : X_LUT4
    generic map(
      INIT => X"CFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16,
      ADR2 => tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_2,
      ADR3 => tx_output_crc_loigc_Mxor_CO_12_Xo(1),
      O => tx_output_n0034(12)
    );
  tx_output_crcl_12_XUSED : X_BUF
    port map (
      I => tx_output_crcl_12_FROM,
      O => tx_output_crc_loigc_Mxor_CO_12_Xo(1)
    );
  tx_output_ldata_2_18 : X_LUT4
    generic map(
      INIT => X"F088"
    )
    port map (
      ADR0 => q2(10),
      ADR1 => tx_output_N81613,
      ADR2 => q2(2),
      ADR3 => tx_output_cs_FFd6,
      O => tx_output_data_2_FROM
    );
  tx_output_ldata_2_25 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_CHOICE1253,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1261,
      O => tx_output_ldata(2)
    );
  tx_output_data_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_data_2_CEMUXNOT
    );
  tx_output_data_2_XUSED : X_BUF
    port map (
      I => tx_output_data_2_FROM,
      O => tx_output_CHOICE1261
    );
  tx_output_ldata_3_18 : X_LUT4
    generic map(
      INIT => X"EA40"
    )
    port map (
      ADR0 => tx_output_cs_FFd6,
      ADR1 => tx_output_N81625,
      ADR2 => q2(11),
      ADR3 => q2(3),
      O => tx_output_data_3_FROM
    );
  tx_output_ldata_3_25 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_CHOICE1265,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1273,
      O => tx_output_ldata(3)
    );
  tx_output_data_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_data_3_CEMUXNOT
    );
  tx_output_data_3_XUSED : X_BUF
    port map (
      I => tx_output_data_3_FROM,
      O => tx_output_CHOICE1273
    );
  mac_control_Mmux_n0017_Result_2_149_SW0 : X_LUT4
    generic map(
      INIT => X"0015"
    )
    port map (
      ADR0 => mac_control_CHOICE2280,
      ADR1 => mac_control_n0085,
      ADR2 => mac_control_lmacaddr(2),
      ADR3 => mac_control_CHOICE2297,
      O => mac_control_dout_2_FROM
    );
  mac_control_Mmux_n0017_Result_2_149 : X_LUT4
    generic map(
      INIT => X"222E"
    )
    port map (
      ADR0 => mac_control_dout(1),
      ADR1 => mac_control_n0060,
      ADR2 => mac_control_addr(5),
      ADR3 => mac_control_N81645,
      O => mac_control_N76751
    );
  mac_control_dout_2_XUSED : X_BUF
    port map (
      I => mac_control_dout_2_FROM,
      O => mac_control_N81645
    );
  tx_output_ldata_4_18 : X_LUT4
    generic map(
      INIT => X"AAC0"
    )
    port map (
      ADR0 => q2(4),
      ADR1 => q2(12),
      ADR2 => tx_output_N81609,
      ADR3 => tx_output_cs_FFd6,
      O => tx_output_data_4_FROM
    );
  tx_output_ldata_4_25 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_CHOICE1241,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1249,
      O => tx_output_ldata(4)
    );
  tx_output_data_4_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_data_4_CEMUXNOT
    );
  tx_output_data_4_XUSED : X_BUF
    port map (
      I => tx_output_data_4_FROM,
      O => tx_output_CHOICE1249
    );
  tx_output_ltxd_6_SW0 : X_LUT4
    generic map(
      INIT => X"EEAA"
    )
    port map (
      ADR0 => tx_output_outselll(1),
      ADR1 => tx_output_datal(6),
      ADR2 => VCC,
      ADR3 => tx_output_outselll(0),
      O => tx_output_N70503_FROM
    );
  tx_output_ltxd_6_Q : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => tx_output_outselll(2),
      ADR1 => tx_output_ncrcbytel(1),
      ADR2 => tx_output_outselll(3),
      ADR3 => tx_output_N70503,
      O => tx_output_N70503_GROM
    );
  tx_output_N70503_XUSED : X_BUF
    port map (
      I => tx_output_N70503_FROM,
      O => tx_output_N70503
    );
  tx_output_N70503_YUSED : X_BUF
    port map (
      I => tx_output_N70503_GROM,
      O => tx_output_ltxd(6)
    );
  tx_output_ldata_5_18 : X_LUT4
    generic map(
      INIT => X"E2C0"
    )
    port map (
      ADR0 => q2(13),
      ADR1 => tx_output_cs_FFd6,
      ADR2 => q2(5),
      ADR3 => tx_output_N81617,
      O => tx_output_data_5_FROM
    );
  tx_output_ldata_5_25 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_CHOICE1229,
      ADR3 => tx_output_CHOICE1237,
      O => tx_output_ldata(5)
    );
  tx_output_data_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_data_5_CEMUXNOT
    );
  tx_output_data_5_XUSED : X_BUF
    port map (
      I => tx_output_data_5_FROM,
      O => tx_output_CHOICE1237
    );
  tx_output_ldata_6_18 : X_LUT4
    generic map(
      INIT => X"F088"
    )
    port map (
      ADR0 => tx_output_N81625,
      ADR1 => q2(14),
      ADR2 => q2(6),
      ADR3 => tx_output_cs_FFd6,
      O => tx_output_data_6_FROM
    );
  tx_output_ldata_6_25 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_CHOICE1217,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1225,
      O => tx_output_ldata(6)
    );
  tx_output_data_6_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_data_6_CEMUXNOT
    );
  tx_output_data_6_XUSED : X_BUF
    port map (
      I => tx_output_data_6_FROM,
      O => tx_output_CHOICE1225
    );
  tx_output_ldata_7_18 : X_LUT4
    generic map(
      INIT => X"B888"
    )
    port map (
      ADR0 => q2(7),
      ADR1 => tx_output_cs_FFd6,
      ADR2 => q2(15),
      ADR3 => tx_output_N81605,
      O => tx_output_data_7_FROM
    );
  tx_output_ldata_7_25 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_CHOICE1205,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1213,
      O => tx_output_ldata(7)
    );
  tx_output_data_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_data_7_CEMUXNOT
    );
  tx_output_data_7_XUSED : X_BUF
    port map (
      I => tx_output_data_7_FROM,
      O => tx_output_CHOICE1213
    );
  tx_output_cs_Out1160_2_177 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => tx_output_cs_FFd4,
      ADR1 => tx_output_cs_FFd5,
      ADR2 => VCC,
      ADR3 => tx_output_cs_FFd6,
      O => tx_output_cs_Out1160_2_FROM
    );
  tx_output_ldata_0_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => tx_output_cs_FFd4,
      ADR1 => q2(16),
      ADR2 => tx_output_cs_FFd5,
      ADR3 => q2(24),
      O => tx_output_cs_Out1160_2_GROM
    );
  tx_output_cs_Out1160_2_XUSED : X_BUF
    port map (
      I => tx_output_cs_Out1160_2_FROM,
      O => tx_output_cs_Out1160_2
    );
  tx_output_cs_Out1160_2_YUSED : X_BUF
    port map (
      I => tx_output_cs_Out1160_2_GROM,
      O => tx_output_CHOICE1289
    );
  tx_output_ldata_5_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => tx_output_cs_FFd5,
      ADR1 => q2(29),
      ADR2 => tx_output_cs_FFd4,
      ADR3 => q2(21),
      O => tx_output_CHOICE1229_FROM
    );
  tx_output_ldata_1_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => tx_output_cs_FFd4,
      ADR1 => tx_output_cs_FFd5,
      ADR2 => q2(17),
      ADR3 => q2(25),
      O => tx_output_CHOICE1229_GROM
    );
  tx_output_CHOICE1229_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1229_FROM,
      O => tx_output_CHOICE1229
    );
  tx_output_CHOICE1229_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1229_GROM,
      O => tx_output_CHOICE1277
    );
  tx_output_ltxd_7_SW0 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_datal(7),
      ADR2 => VCC,
      ADR3 => tx_output_outselll(0),
      O => tx_output_N69304_FROM
    );
  tx_output_ltxd_7_Q : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => tx_output_outselll(3),
      ADR1 => tx_output_outselll(2),
      ADR2 => tx_output_ncrcbytel(0),
      ADR3 => tx_output_N69304,
      O => tx_output_N69304_GROM
    );
  tx_output_N69304_XUSED : X_BUF
    port map (
      I => tx_output_N69304_FROM,
      O => tx_output_N69304
    );
  tx_output_N69304_YUSED : X_BUF
    port map (
      I => tx_output_N69304_GROM,
      O => tx_output_ltxd(7)
    );
  tx_output_ldata_3_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => q2(19),
      ADR1 => tx_output_cs_FFd4,
      ADR2 => tx_output_cs_FFd5,
      ADR3 => q2(27),
      O => tx_output_CHOICE1265_FROM
    );
  tx_output_ldata_2_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => q2(26),
      ADR1 => tx_output_cs_FFd4,
      ADR2 => q2(18),
      ADR3 => tx_output_cs_FFd5,
      O => tx_output_CHOICE1265_GROM
    );
  tx_output_CHOICE1265_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1265_FROM,
      O => tx_output_CHOICE1265
    );
  tx_output_CHOICE1265_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1265_GROM,
      O => tx_output_CHOICE1253
    );
  tx_output_ldata_7_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => q2(31),
      ADR1 => tx_output_cs_FFd4,
      ADR2 => tx_output_cs_FFd5,
      ADR3 => q2(23),
      O => tx_output_CHOICE1205_FROM
    );
  tx_output_ldata_4_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => q2(20),
      ADR1 => q2(28),
      ADR2 => tx_output_cs_FFd4,
      ADR3 => tx_output_cs_FFd5,
      O => tx_output_CHOICE1205_GROM
    );
  tx_output_CHOICE1205_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1205_FROM,
      O => tx_output_CHOICE1205
    );
  tx_output_CHOICE1205_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1205_GROM,
      O => tx_output_CHOICE1241
    );
  tx_output_ldata_6_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => q2(22),
      ADR1 => q2(30),
      ADR2 => tx_output_cs_FFd5,
      ADR3 => tx_output_cs_FFd4,
      O => tx_output_CHOICE1217_GROM
    );
  tx_output_CHOICE1217_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1217_GROM,
      O => tx_output_CHOICE1217
    );
  RESET_IBUF_1_178 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => RESET_IBUF_1_FROM
    );
  tx_input_n00331 : X_LUT4
    generic map(
      INIT => X"00FE"
    )
    port map (
      ADR0 => tx_input_cs_FFd9,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => tx_input_cs_FFd5,
      ADR3 => RESET_IBUF_1,
      O => RESET_IBUF_1_GROM
    );
  RESET_IBUF_1_XUSED : X_BUF
    port map (
      I => RESET_IBUF_1_FROM,
      O => RESET_IBUF_1
    );
  RESET_IBUF_1_YUSED : X_BUF
    port map (
      I => RESET_IBUF_1_GROM,
      O => tx_input_n0033
    );
  RESET_IBUF_2_179 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => RESET_IBUF_2_FROM
    );
  rx_input_fifo_control_n00081 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => RESET_IBUF_2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_ce,
      O => RESET_IBUF_2_GROM
    );
  RESET_IBUF_2_XUSED : X_BUF
    port map (
      I => RESET_IBUF_2_FROM,
      O => RESET_IBUF_2
    );
  RESET_IBUF_2_YUSED : X_BUF
    port map (
      I => RESET_IBUF_2_GROM,
      O => rx_input_fifo_control_n0008
    );
  mac_control_PHY_status_MII_Interface_iobuffer_OBUFT : X_TRI
    port map (
      I => MDIO_OUTMUX,
      CTL => MDIO_ENABLE,
      O => MDIO
    );
  MDIO_ENABLEINV : X_INV
    port map (
      I => MDIO_TORGTS,
      O => MDIO_ENABLE
    );
  MDIO_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => mac_control_PHY_status_MII_Interface_sts,
      O => MDIO_TORGTS
    );
  MDIO_OUTMUX_180 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_sout,
      O => MDIO_OUTMUX
    );
  mac_control_PHY_status_MII_Interface_iobuffer_IBUF : X_BUF
    port map (
      I => MDIO,
      O => mac_control_PHY_status_MII_Interface_sin
    );
  rx_input_fifo_fifo_BU220 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3647,
      CE => rx_input_fifo_fifo_N3646,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_empty_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_empty
    );
  rx_input_fifo_fifo_empty_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_empty_FFX_SET
    );
  rx_output_DOUT_10_OBUF_181 : X_TRI
    port map (
      I => DOUT_10_OUTMUX,
      CTL => DOUT_10_ENABLE,
      O => DOUT(10)
    );
  DOUT_10_ENABLEINV : X_INV
    port map (
      I => DOUT_10_TORGTS,
      O => DOUT_10_ENABLE
    );
  DOUT_10_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_10_TORGTS
    );
  DOUT_10_OUTMUX_182 : X_BUF
    port map (
      I => rx_output_DOUT_10_OBUF,
      O => DOUT_10_OUTMUX
    );
  DOUT_10_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(10),
      O => DOUT_10_OD
    );
  rx_output_DOUT_11_OBUF_183 : X_TRI
    port map (
      I => DOUT_11_OUTMUX,
      CTL => DOUT_11_ENABLE,
      O => DOUT(11)
    );
  DOUT_11_ENABLEINV : X_INV
    port map (
      I => DOUT_11_TORGTS,
      O => DOUT_11_ENABLE
    );
  DOUT_11_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_11_TORGTS
    );
  DOUT_11_OUTMUX_184 : X_BUF
    port map (
      I => rx_output_DOUT_11_OBUF,
      O => DOUT_11_OUTMUX
    );
  DOUT_11_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(11),
      O => DOUT_11_OD
    );
  rx_output_DOUT_12_OBUF_185 : X_TRI
    port map (
      I => DOUT_12_OUTMUX,
      CTL => DOUT_12_ENABLE,
      O => DOUT(12)
    );
  DOUT_12_ENABLEINV : X_INV
    port map (
      I => DOUT_12_TORGTS,
      O => DOUT_12_ENABLE
    );
  DOUT_12_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_12_TORGTS
    );
  DOUT_12_OUTMUX_186 : X_BUF
    port map (
      I => rx_output_DOUT_12_OBUF,
      O => DOUT_12_OUTMUX
    );
  DOUT_12_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(12),
      O => DOUT_12_OD
    );
  rx_output_DOUT_13_OBUF_187 : X_TRI
    port map (
      I => DOUT_13_OUTMUX,
      CTL => DOUT_13_ENABLE,
      O => DOUT(13)
    );
  DOUT_13_ENABLEINV : X_INV
    port map (
      I => DOUT_13_TORGTS,
      O => DOUT_13_ENABLE
    );
  DOUT_13_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_13_TORGTS
    );
  DOUT_13_OUTMUX_188 : X_BUF
    port map (
      I => rx_output_DOUT_13_OBUF,
      O => DOUT_13_OUTMUX
    );
  DOUT_13_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(13),
      O => DOUT_13_OD
    );
  rx_output_DOUT_14_OBUF_189 : X_TRI
    port map (
      I => DOUT_14_OUTMUX,
      CTL => DOUT_14_ENABLE,
      O => DOUT(14)
    );
  DOUT_14_ENABLEINV : X_INV
    port map (
      I => DOUT_14_TORGTS,
      O => DOUT_14_ENABLE
    );
  DOUT_14_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_14_TORGTS
    );
  DOUT_14_OUTMUX_190 : X_BUF
    port map (
      I => rx_output_DOUT_14_OBUF,
      O => DOUT_14_OUTMUX
    );
  DOUT_14_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(14),
      O => DOUT_14_OD
    );
  rx_output_DOUT_15_OBUF_191 : X_TRI
    port map (
      I => DOUT_15_OUTMUX,
      CTL => DOUT_15_ENABLE,
      O => DOUT(15)
    );
  DOUT_15_ENABLEINV : X_INV
    port map (
      I => DOUT_15_TORGTS,
      O => DOUT_15_ENABLE
    );
  DOUT_15_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_15_TORGTS
    );
  DOUT_15_OUTMUX_192 : X_BUF
    port map (
      I => rx_output_DOUT_15_OBUF,
      O => DOUT_15_OUTMUX
    );
  DOUT_15_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(15),
      O => DOUT_15_OD
    );
  rx_input_fifo_fifo_BU214 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2477,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2497_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2497
    );
  rx_input_fifo_fifo_N2497_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2497_FFY_SET
    );
  MDC_OBUF_193 : X_TRI
    port map (
      I => MDC_OUTMUX,
      CTL => MDC_ENABLE,
      O => MDC
    );
  MDC_ENABLEINV : X_INV
    port map (
      I => MDC_TORGTS,
      O => MDC_ENABLE
    );
  MDC_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MDC_TORGTS
    );
  MDC_OUTMUX_194 : X_BUF
    port map (
      I => MDC_OBUF,
      O => MDC_OUTMUX
    );
  SCS_IMUX : X_BUF
    port map (
      I => SCS_IBUF_1,
      O => SCS_IBUF
    );
  SCS_IBUF_195 : X_BUF
    port map (
      I => SCS,
      O => SCS_IBUF_1
    );
  SIN_IMUX : X_BUF
    port map (
      I => SIN_IBUF_2,
      O => SIN_IBUF
    );
  SIN_IBUF_196 : X_BUF
    port map (
      I => SIN,
      O => SIN_IBUF_2
    );
  mac_control_LED100_OBUF_197 : X_TRI
    port map (
      I => LED100_OUTMUX,
      CTL => LED100_ENABLE,
      O => LED100
    );
  LED100_ENABLEINV : X_INV
    port map (
      I => LED100_TORGTS,
      O => LED100_ENABLE
    );
  LED100_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LED100_TORGTS
    );
  LED100_OUTMUX_198 : X_BUF
    port map (
      I => mac_control_LED100_OBUF,
      O => LED100_OUTMUX
    );
  LED100_OMUX : X_BUF
    port map (
      I => mac_control_n0037,
      O => LED100_OD
    );
  rx_input_fifo_fifo_BU171 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3560,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2397_FFY_RST,
      O => rx_input_fifo_fifo_N2398
    );
  rx_input_fifo_fifo_N2397_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2397_FFY_RST
    );
  MCLK_OBUF_199 : X_TRI
    port map (
      I => MCLK_OUTMUX,
      CTL => MCLK_ENABLE,
      O => MCLK
    );
  MCLK_ENABLEINV : X_INV
    port map (
      I => MCLK_TORGTS,
      O => MCLK_ENABLE
    );
  MCLK_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MCLK_TORGTS
    );
  MCLK_OUTMUX_200 : X_BUF
    port map (
      I => MCLK_OBUF,
      O => MCLK_OUTMUX
    );
  tx_input_NEWFRAME_IBUF_201 : X_BUF
    port map (
      I => NEWFRAME,
      O => tx_input_NEWFRAME_IBUF
    );
  mac_control_LED1000_OBUF_202 : X_TRI
    port map (
      I => LED1000_OUTMUX,
      CTL => LED1000_ENABLE,
      O => LED1000
    );
  LED1000_ENABLEINV : X_INV
    port map (
      I => LED1000_TORGTS,
      O => LED1000_ENABLE
    );
  LED1000_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LED1000_TORGTS
    );
  LED1000_OUTMUX_203 : X_BUF
    port map (
      I => mac_control_LED1000_OBUF,
      O => LED1000_OUTMUX
    );
  LED1000_OMUX : X_BUF
    port map (
      I => mac_control_n0036,
      O => LED1000_OD
    );
  tx_output_TX_EN_OBUF : X_TRI
    port map (
      I => TX_EN_OUTMUX,
      CTL => TX_EN_ENABLE,
      O => TX_EN
    );
  TX_EN_ENABLEINV : X_INV
    port map (
      I => TX_EN_TORGTS,
      O => TX_EN_ENABLE
    );
  TX_EN_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TX_EN_TORGTS
    );
  TX_EN_OUTMUX_204 : X_BUF
    port map (
      I => tx_output_TXEN,
      O => TX_EN_OUTMUX
    );
  TX_EN_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => TX_EN_OCEMUXNOT
    );
  TX_EN_OMUX : X_BUF
    port map (
      I => tx_output_ltxen3,
      O => TX_EN_OD
    );
  rx_output_DOUTEN_OBUF_205 : X_TRI
    port map (
      I => DOUTEN_OUTMUX,
      CTL => DOUTEN_ENABLE,
      O => DOUTEN
    );
  DOUTEN_ENABLEINV : X_INV
    port map (
      I => DOUTEN_TORGTS,
      O => DOUTEN_ENABLE
    );
  DOUTEN_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUTEN_TORGTS
    );
  DOUTEN_OUTMUX_206 : X_BUF
    port map (
      I => rx_output_DOUTEN_OBUF,
      O => DOUTEN_OUTMUX
    );
  DOUTEN_OMUX : X_BUF
    port map (
      I => rx_output_ldouten2,
      O => DOUTEN_OD
    );
  memcontroller_MWE_OBUF : X_TRI
    port map (
      I => MWE_OUTMUX,
      CTL => MWE_ENABLE,
      O => MWE
    );
  MWE_ENABLEINV : X_INV
    port map (
      I => MWE_TORGTS,
      O => MWE_ENABLE
    );
  MWE_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MWE_TORGTS
    );
  MWE_OUTMUX_207 : X_BUF
    port map (
      I => memcontroller_WEEXT,
      O => MWE_OUTMUX
    );
  MWE_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MWE_OCEMUXNOT
    );
  MWE_OMUX : X_BUF
    port map (
      I => memcontroller_n0116,
      O => MWE_OD
    );
  RESET_IMUX : X_BUF
    port map (
      I => RESET_IBUF_3,
      O => RESET_IBUF
    );
  RESET_IBUF_208 : X_BUF
    port map (
      I => RESET,
      O => RESET_IBUF_3
    );
  rx_output_NEXTFRAME_IBUF_209 : X_BUF
    port map (
      I => NEXTFRAME,
      O => rx_output_NEXTFRAME_IBUF
    );
  mac_control_LEDACT_OBUF_210 : X_TRI
    port map (
      I => LEDACT_OUTMUX,
      CTL => LEDACT_ENABLE,
      O => LEDACT
    );
  LEDACT_ENABLEINV : X_INV
    port map (
      I => LEDACT_TORGTS,
      O => LEDACT_ENABLE
    );
  LEDACT_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDACT_TORGTS
    );
  LEDACT_OUTMUX_211 : X_BUF
    port map (
      I => mac_control_LEDACT_OBUF,
      O => LEDACT_OUTMUX
    );
  LEDACT_OMUX : X_BUF
    port map (
      I => mac_control_phystat(2),
      O => LEDACT_OD
    );
  tx_output_TXD_0_OBUF_212 : X_TRI
    port map (
      I => TXD_0_OUTMUX,
      CTL => TXD_0_ENABLE,
      O => TXD(0)
    );
  TXD_0_ENABLEINV : X_INV
    port map (
      I => TXD_0_TORGTS,
      O => TXD_0_ENABLE
    );
  TXD_0_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_0_TORGTS
    );
  TXD_0_OUTMUX_213 : X_BUF
    port map (
      I => tx_output_TXD_0_OBUF,
      O => TXD_0_OUTMUX
    );
  TXD_0_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => TXD_0_OCEMUXNOT
    );
  TXD_0_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(0),
      O => TXD_0_OD
    );
  tx_output_TXD_1_OBUF_214 : X_TRI
    port map (
      I => TXD_1_OUTMUX,
      CTL => TXD_1_ENABLE,
      O => TXD(1)
    );
  TXD_1_ENABLEINV : X_INV
    port map (
      I => TXD_1_TORGTS,
      O => TXD_1_ENABLE
    );
  TXD_1_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_1_TORGTS
    );
  TXD_1_OUTMUX_215 : X_BUF
    port map (
      I => tx_output_TXD_1_OBUF,
      O => TXD_1_OUTMUX
    );
  TXD_1_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => TXD_1_OCEMUXNOT
    );
  TXD_1_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(1),
      O => TXD_1_OD
    );
  tx_output_TXD_2_OBUF_216 : X_TRI
    port map (
      I => TXD_2_OUTMUX,
      CTL => TXD_2_ENABLE,
      O => TXD(2)
    );
  TXD_2_ENABLEINV : X_INV
    port map (
      I => TXD_2_TORGTS,
      O => TXD_2_ENABLE
    );
  TXD_2_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_2_TORGTS
    );
  TXD_2_OUTMUX_217 : X_BUF
    port map (
      I => tx_output_TXD_2_OBUF,
      O => TXD_2_OUTMUX
    );
  TXD_2_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => TXD_2_OCEMUXNOT
    );
  TXD_2_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(2),
      O => TXD_2_OD
    );
  tx_output_TXD_3_OBUF_218 : X_TRI
    port map (
      I => TXD_3_OUTMUX,
      CTL => TXD_3_ENABLE,
      O => TXD(3)
    );
  TXD_3_ENABLEINV : X_INV
    port map (
      I => TXD_3_TORGTS,
      O => TXD_3_ENABLE
    );
  TXD_3_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_3_TORGTS
    );
  TXD_3_OUTMUX_219 : X_BUF
    port map (
      I => tx_output_TXD_3_OBUF,
      O => TXD_3_OUTMUX
    );
  TXD_3_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => TXD_3_OCEMUXNOT
    );
  TXD_3_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(3),
      O => TXD_3_OD
    );
  tx_output_TXD_4_OBUF_220 : X_TRI
    port map (
      I => TXD_4_OUTMUX,
      CTL => TXD_4_ENABLE,
      O => TXD(4)
    );
  TXD_4_ENABLEINV : X_INV
    port map (
      I => TXD_4_TORGTS,
      O => TXD_4_ENABLE
    );
  TXD_4_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_4_TORGTS
    );
  TXD_4_OUTMUX_221 : X_BUF
    port map (
      I => tx_output_TXD_4_OBUF,
      O => TXD_4_OUTMUX
    );
  TXD_4_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => TXD_4_OCEMUXNOT
    );
  TXD_4_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(4),
      O => TXD_4_OD
    );
  tx_output_TXD_5_OBUF_222 : X_TRI
    port map (
      I => TXD_5_OUTMUX,
      CTL => TXD_5_ENABLE,
      O => TXD(5)
    );
  TXD_5_ENABLEINV : X_INV
    port map (
      I => TXD_5_TORGTS,
      O => TXD_5_ENABLE
    );
  TXD_5_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_5_TORGTS
    );
  TXD_5_OUTMUX_223 : X_BUF
    port map (
      I => tx_output_TXD_5_OBUF,
      O => TXD_5_OUTMUX
    );
  TXD_5_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => TXD_5_OCEMUXNOT
    );
  TXD_5_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(5),
      O => TXD_5_OD
    );
  rx_input_fifo_fifo_BU106 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2814,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N13_FFY_RST,
      O => rx_input_fifo_fifo_N12
    );
  rx_input_fifo_fifo_N13_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N13_FFY_RST
    );
  tx_output_TXD_6_OBUF_224 : X_TRI
    port map (
      I => TXD_6_OUTMUX,
      CTL => TXD_6_ENABLE,
      O => TXD(6)
    );
  TXD_6_ENABLEINV : X_INV
    port map (
      I => TXD_6_TORGTS,
      O => TXD_6_ENABLE
    );
  TXD_6_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_6_TORGTS
    );
  TXD_6_OUTMUX_225 : X_BUF
    port map (
      I => tx_output_TXD_6_OBUF,
      O => TXD_6_OUTMUX
    );
  TXD_6_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => TXD_6_OCEMUXNOT
    );
  TXD_6_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(6),
      O => TXD_6_OD
    );
  tx_output_TXD_7_OBUF_226 : X_TRI
    port map (
      I => TXD_7_OUTMUX,
      CTL => TXD_7_ENABLE,
      O => TXD(7)
    );
  TXD_7_ENABLEINV : X_INV
    port map (
      I => TXD_7_TORGTS,
      O => TXD_7_ENABLE
    );
  TXD_7_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_7_TORGTS
    );
  TXD_7_OUTMUX_227 : X_BUF
    port map (
      I => tx_output_TXD_7_OBUF,
      O => TXD_7_OUTMUX
    );
  TXD_7_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => TXD_7_OCEMUXNOT
    );
  TXD_7_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(7),
      O => TXD_7_OD
    );
  tx_output_crc_loigc_Mxor_CO_23_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(25),
      ADR1 => tx_output_data(6),
      ADR2 => tx_output_data(7),
      ADR3 => tx_output_crcl(24),
      O => tx_output_crcl_23_FROM
    );
  tx_output_n0034_23_1 : X_LUT4
    generic map(
      INIT => X"F3FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_crc_loigc_Mxor_CO_23_Xo_2_1_2,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crc_loigc_Mxor_CO_23_Xo(0),
      O => tx_output_n0034(23)
    );
  tx_output_crcl_23_XUSED : X_BUF
    port map (
      I => tx_output_crcl_23_FROM,
      O => tx_output_crc_loigc_Mxor_CO_23_Xo(0)
    );
  tx_output_crc_loigc_Mxor_CO_15_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_Mxor_CO_13_Xo(2),
      ADR1 => tx_output_crc_loigc_n0118(0),
      ADR2 => tx_output_crc_loigc_n0115(0),
      ADR3 => tx_output_crcl(7),
      O => tx_output_crcl_15_FROM
    );
  tx_output_n0034_15_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crc_15_Q,
      O => tx_output_n0034(15)
    );
  tx_output_crcl_15_XUSED : X_BUF
    port map (
      I => tx_output_crcl_15_FROM,
      O => tx_output_crc_15_Q
    );
  mac_control_Mmux_n0017_Result_5_149_SW0 : X_LUT4
    generic map(
      INIT => X"0103"
    )
    port map (
      ADR0 => mac_control_n0085,
      ADR1 => mac_control_CHOICE2373,
      ADR2 => mac_control_CHOICE2356,
      ADR3 => mac_control_lmacaddr(5),
      O => mac_control_dout_5_FROM
    );
  mac_control_Mmux_n0017_Result_5_149 : X_LUT4
    generic map(
      INIT => X"5072"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_addr(5),
      ADR2 => mac_control_dout(4),
      ADR3 => mac_control_N81649,
      O => mac_control_N77167
    );
  mac_control_dout_5_XUSED : X_BUF
    port map (
      I => mac_control_dout_5_FROM,
      O => mac_control_N81649
    );
  rx_input_memio_crccomb_Mxor_CO_10_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_Mxor_CO_7_Xo(1),
      ADR1 => rx_input_memio_crccomb_n0118(0),
      ADR2 => rx_input_memio_crcl(2),
      ADR3 => rx_input_memio_crccomb_n0118(1),
      O => rx_input_memio_crcl_10_FROM
    );
  rx_input_memio_n0048_10_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_10_Q,
      O => rx_input_memio_n0048(10)
    );
  rx_input_memio_crcl_10_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_10_FROM,
      O => rx_input_memio_crc_10_Q
    );
  mac_control_lmacaddr_47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_47_FFX_RST,
      O => mac_control_lmacaddr(47)
    );
  mac_control_lmacaddr_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_47_FFX_RST
    );
  mac_control_phydo_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_3_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(2),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_3_FFY_RST,
      O => mac_control_phydo(2)
    );
  rx_input_memio_crccomb_Mxor_CO_8_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0115(0),
      ADR1 => rx_input_memio_crccomb_Mxor_CO_7_Xo(1),
      ADR2 => rx_input_memio_crccomb_n0122(0),
      ADR3 => rx_input_memio_crcl(0),
      O => rx_input_memio_crcl_8_FROM
    );
  rx_input_memio_n0048_8_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_8_Q,
      O => rx_input_memio_n0048(8)
    );
  rx_input_memio_crcl_8_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_8_FROM,
      O => rx_input_memio_crc_8_Q
    );
  mac_control_Mmux_n0017_Result_8_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_N52132,
      ADR1 => mac_control_phystat(8),
      ADR2 => mac_control_phydo(8),
      ADR3 => mac_control_N52125,
      O => mac_control_CHOICE2382_FROM
    );
  mac_control_Mmux_n0017_Result_0_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phystat(0),
      ADR1 => mac_control_N52132,
      ADR2 => mac_control_phydo(0),
      ADR3 => mac_control_N52125,
      O => mac_control_CHOICE2382_GROM
    );
  mac_control_CHOICE2382_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2382_FROM,
      O => mac_control_CHOICE2382
    );
  mac_control_CHOICE2382_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2382_GROM,
      O => mac_control_CHOICE2194
    );
  mac_control_Mmux_n0017_Result_14_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_N52125,
      ADR1 => mac_control_N52132,
      ADR2 => mac_control_phystat(14),
      ADR3 => mac_control_phydo(14),
      O => mac_control_CHOICE2458_FROM
    );
  mac_control_Mmux_n0017_Result_1_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_N52132,
      ADR1 => mac_control_N52125,
      ADR2 => mac_control_phydo(1),
      ADR3 => mac_control_phystat(1),
      O => mac_control_CHOICE2458_GROM
    );
  mac_control_CHOICE2458_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2458_FROM,
      O => mac_control_CHOICE2458
    );
  mac_control_CHOICE2458_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2458_GROM,
      O => mac_control_CHOICE2230
    );
  mac_control_Mmux_n0017_Result_6_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_N52132,
      ADR1 => mac_control_phydo(6),
      ADR2 => mac_control_phystat(6),
      ADR3 => mac_control_N52125,
      O => mac_control_CHOICE2306_FROM
    );
  mac_control_Mmux_n0017_Result_2_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_N52132,
      ADR1 => mac_control_phydo(2),
      ADR2 => mac_control_phystat(2),
      ADR3 => mac_control_N52125,
      O => mac_control_CHOICE2306_GROM
    );
  mac_control_CHOICE2306_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2306_FROM,
      O => mac_control_CHOICE2306
    );
  mac_control_CHOICE2306_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2306_GROM,
      O => mac_control_CHOICE2268
    );
  mac_control_Mmux_n0017_Result_10_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_N52125,
      ADR1 => mac_control_phydo(10),
      ADR2 => mac_control_phystat(10),
      ADR3 => mac_control_N52132,
      O => mac_control_CHOICE2420_FROM
    );
  mac_control_Mmux_n0017_Result_5_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phydo(5),
      ADR1 => mac_control_N52125,
      ADR2 => mac_control_phystat(5),
      ADR3 => mac_control_N52132,
      O => mac_control_CHOICE2420_GROM
    );
  mac_control_CHOICE2420_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2420_FROM,
      O => mac_control_CHOICE2420
    );
  mac_control_CHOICE2420_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2420_GROM,
      O => mac_control_CHOICE2344
    );
  memcontroller_dnl2_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_11_CEMUXNOT
    );
  memcontroller_dnl2_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_21_CEMUXNOT
    );
  rx_input_memio_BPOUT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_11_58,
      CE => rxbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_11_FFX_RST,
      O => rxbp(11)
    );
  rxbp_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_11_FFX_RST
    );
  memcontroller_dnl2_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_13_CEMUXNOT
    );
  memcontroller_dnl2_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_31_CEMUXNOT
    );
  memcontroller_dnl2_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_23_CEMUXNOT
    );
  memcontroller_dnl2_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_15_CEMUXNOT
    );
  memcontroller_dnl2_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_25_CEMUXNOT
    );
  memcontroller_dnl2_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_17_CEMUXNOT
    );
  memcontroller_dnl2_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_27_CEMUXNOT
    );
  memcontroller_dnl2_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_19_CEMUXNOT
    );
  memcontroller_dnl2_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_29_CEMUXNOT
    );
  rx_input_memio_datal_1_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_datal_1_CEMUXNOT
    );
  rx_input_memio_datal_3_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_datal_3_CEMUXNOT
    );
  rx_input_memio_BPOUT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_14_55,
      CE => rxbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_15_FFY_RST,
      O => rxbp(14)
    );
  rxbp_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_15_FFY_RST
    );
  rx_input_memio_datal_5_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_datal_5_CEMUXNOT
    );
  rx_input_memio_datal_7_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_datal_7_CEMUXNOT
    );
  rx_input_memio_BPOUT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_13_56,
      CE => rxbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_13_FFX_RST,
      O => rxbp(13)
    );
  rxbp_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_13_FFX_RST
    );
  rx_input_memio_addrchk_lmaceq_0_rt_228 : X_XOR2
    port map (
      I0 => rx_input_memio_addrchk_maceq_0_CYINIT,
      I1 => rx_input_memio_addrchk_maceq_0_FROM,
      O => rx_input_memio_addrchk_lmaceq_0_rt
    );
  rx_input_memio_addrchk_maceq_0_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_maceq_0_FROM
    );
  rx_input_memio_addrchk_maceq_0_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_maceq_0_CEMUXNOT
    );
  rx_input_memio_addrchk_maceq_0_CYINIT_229 : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq(0),
      O => rx_input_memio_addrchk_maceq_0_CYINIT
    );
  rx_input_memio_addrchk_lmaceq_2_rt_230 : X_XOR2
    port map (
      I0 => rx_input_memio_addrchk_maceq_2_CYINIT,
      I1 => rx_input_memio_addrchk_maceq_2_FROM,
      O => rx_input_memio_addrchk_lmaceq_2_rt
    );
  rx_input_memio_addrchk_maceq_2_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_maceq_2_FROM
    );
  rx_input_memio_addrchk_maceq_2_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_maceq_2_CEMUXNOT
    );
  rx_input_memio_addrchk_maceq_2_CYINIT_231 : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq(2),
      O => rx_input_memio_addrchk_maceq_2_CYINIT
    );
  rx_input_memio_addrchk_lmaceq_4_rt_232 : X_XOR2
    port map (
      I0 => rx_input_memio_addrchk_maceq_4_CYINIT,
      I1 => rx_input_memio_addrchk_maceq_4_FROM,
      O => rx_input_memio_addrchk_lmaceq_4_rt
    );
  rx_input_memio_addrchk_maceq_4_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_maceq_4_FROM
    );
  rx_input_memio_addrchk_maceq_4_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_maceq_4_CEMUXNOT
    );
  rx_input_memio_addrchk_maceq_4_CYINIT_233 : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq(4),
      O => rx_input_memio_addrchk_maceq_4_CYINIT
    );
  tx_output_crc_loigc_Mxor_CO_24_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(16),
      ADR1 => tx_output_crc_loigc_n0118(1),
      ADR2 => tx_output_crc_loigc_n0124(0),
      ADR3 => tx_output_crc_loigc_n0122(0),
      O => tx_output_crcl_24_FROM
    );
  tx_output_n0034_24_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16,
      ADR2 => VCC,
      ADR3 => tx_output_crc_24_Q,
      O => tx_output_n0034(24)
    );
  tx_output_crcl_24_XUSED : X_BUF
    port map (
      I => tx_output_crcl_24_FROM,
      O => tx_output_crc_24_Q
    );
  tx_output_crc_loigc_Mxor_CO_16_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0115(0),
      ADR1 => tx_output_crc_loigc_n0118(0),
      ADR2 => tx_output_crc_loigc_n0122(1),
      ADR3 => tx_output_crcl(8),
      O => tx_output_crcl_16_FROM
    );
  tx_output_n0034_16_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crc_16_Q,
      O => tx_output_n0034(16)
    );
  tx_output_crcl_16_XUSED : X_BUF
    port map (
      I => tx_output_crcl_16_FROM,
      O => tx_output_crc_16_Q
    );
  mac_control_Mmux_n0017_Result_6_149_SW0 : X_LUT4
    generic map(
      INIT => X"0007"
    )
    port map (
      ADR0 => mac_control_lmacaddr(6),
      ADR1 => mac_control_n0085,
      ADR2 => mac_control_CHOICE2335,
      ADR3 => mac_control_CHOICE2318,
      O => mac_control_dout_6_FROM
    );
  mac_control_Mmux_n0017_Result_6_149 : X_LUT4
    generic map(
      INIT => X"5072"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_addr(5),
      ADR2 => mac_control_dout(5),
      ADR3 => mac_control_N81661,
      O => mac_control_N76959
    );
  mac_control_dout_6_XUSED : X_BUF
    port map (
      I => mac_control_dout_6_FROM,
      O => mac_control_N81661
    );
  rx_input_memio_crccomb_Mxor_CO_11_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0115(0),
      ADR1 => rx_input_memio_crccomb_Mxor_CO_23_Xo(0),
      ADR2 => rx_input_memio_crcl(3),
      ADR3 => rx_input_memio_crccomb_n0124(1),
      O => rx_input_memio_crcl_11_FROM
    );
  rx_input_memio_n0048_11_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_11_Q,
      O => rx_input_memio_n0048(11)
    );
  rx_input_memio_crcl_11_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_11_FROM,
      O => rx_input_memio_crc_11_Q
    );
  mac_control_n0238_234 : X_LUT4
    generic map(
      INIT => X"0040"
    )
    port map (
      ADR0 => mac_control_addr(2),
      ADR1 => mac_control_newcmd,
      ADR2 => mac_control_addr(7),
      ADR3 => mac_control_N70611,
      O => mac_control_n0238_FROM
    );
  mac_control_PHY_status_n00151 : X_LUT4
    generic map(
      INIT => X"3320"
    )
    port map (
      ADR0 => mac_control_n00561_2,
      ADR1 => mac_control_PHY_status_n00151_1,
      ADR2 => mac_control_newcmd,
      ADR3 => mac_control_PHY_status_cs_FFd1,
      O => mac_control_n0238_GROM
    );
  mac_control_n0238_XUSED : X_BUF
    port map (
      I => mac_control_n0238_FROM,
      O => mac_control_n0238
    );
  mac_control_n0238_YUSED : X_BUF
    port map (
      I => mac_control_n0238_GROM,
      O => mac_control_PHY_status_n0015
    );
  rx_input_memio_crccomb_Mxor_CO_9_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0118(1),
      ADR1 => rx_input_memio_crcl(1),
      ADR2 => rx_input_memio_crccomb_Mxor_CO_9_Xo(0),
      ADR3 => rx_input_memio_crccomb_n0118(0),
      O => rx_input_memio_crcl_9_FROM
    );
  rx_input_memio_n0048_9_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_9_Q,
      O => rx_input_memio_n0048(9)
    );
  rx_input_memio_crcl_9_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_9_FROM,
      O => rx_input_memio_crc_9_Q
    );
  memcontroller_MA_13_OBUF : X_TRI
    port map (
      I => MA_13_OUTMUX,
      CTL => MA_13_ENABLE,
      O => MA(13)
    );
  MA_13_ENABLEINV : X_INV
    port map (
      I => MA_13_TORGTS,
      O => MA_13_ENABLE
    );
  MA_13_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_13_TORGTS
    );
  MA_13_OUTMUX_235 : X_BUF
    port map (
      I => memcontroller_ADDREXT(13),
      O => MA_13_OUTMUX
    );
  MA_13_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_13_OCEMUXNOT
    );
  MA_13_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(13),
      O => MA_13_OD
    );
  memcontroller_MA_14_OBUF : X_TRI
    port map (
      I => MA_14_OUTMUX,
      CTL => MA_14_ENABLE,
      O => MA(14)
    );
  MA_14_ENABLEINV : X_INV
    port map (
      I => MA_14_TORGTS,
      O => MA_14_ENABLE
    );
  MA_14_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_14_TORGTS
    );
  MA_14_OUTMUX_236 : X_BUF
    port map (
      I => memcontroller_ADDREXT(14),
      O => MA_14_OUTMUX
    );
  MA_14_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_14_OCEMUXNOT
    );
  MA_14_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(14),
      O => MA_14_OD
    );
  memcontroller_MA_15_OBUF : X_TRI
    port map (
      I => MA_15_OUTMUX,
      CTL => MA_15_ENABLE,
      O => MA(15)
    );
  MA_15_ENABLEINV : X_INV
    port map (
      I => MA_15_TORGTS,
      O => MA_15_ENABLE
    );
  MA_15_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_15_TORGTS
    );
  MA_15_OUTMUX_237 : X_BUF
    port map (
      I => memcontroller_ADDREXT(15),
      O => MA_15_OUTMUX
    );
  MA_15_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_15_OCEMUXNOT
    );
  MA_15_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(15),
      O => MA_15_OD
    );
  memcontroller_MA_16_OBUF : X_TRI
    port map (
      I => MA_16_OUTMUX,
      CTL => MA_16_ENABLE,
      O => MA(16)
    );
  MA_16_ENABLEINV : X_INV
    port map (
      I => MA_16_TORGTS,
      O => MA_16_ENABLE
    );
  MA_16_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_16_TORGTS
    );
  MA_16_OUTMUX_238 : X_BUF
    port map (
      I => memcontroller_ADDREXT(16),
      O => MA_16_OUTMUX
    );
  MA_16_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_16_OCEMUXNOT
    );
  MA_16_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(16),
      O => MA_16_OD
    );
  memcontroller_qdout10_OBUFT : X_TRI
    port map (
      I => MD_10_OUTMUX,
      CTL => MD_10_ENABLE,
      O => MD(10)
    );
  MD_10_ENABLEINV : X_INV
    port map (
      I => MD_10_TORGTS,
      O => MD_10_ENABLE
    );
  MD_10_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(10),
      O => MD_10_TORGTS
    );
  MD_10_OUTMUX_239 : X_BUF
    port map (
      I => memcontroller_dnout(10),
      O => MD_10_OUTMUX
    );
  MD_10_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(10),
      O => MD_10_OD
    );
  memcontroller_qdout10_IBUF : X_BUF
    port map (
      I => MD(10),
      O => memcontroller_q(10)
    );
  memcontroller_qdout11_OBUFT : X_TRI
    port map (
      I => MD_11_OUTMUX,
      CTL => MD_11_ENABLE,
      O => MD(11)
    );
  MD_11_ENABLEINV : X_INV
    port map (
      I => MD_11_TORGTS,
      O => MD_11_ENABLE
    );
  MD_11_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(11),
      O => MD_11_TORGTS
    );
  MD_11_OUTMUX_240 : X_BUF
    port map (
      I => memcontroller_dnout(11),
      O => MD_11_OUTMUX
    );
  MD_11_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(11),
      O => MD_11_OD
    );
  memcontroller_qdout11_IBUF : X_BUF
    port map (
      I => MD(11),
      O => memcontroller_q(11)
    );
  memcontroller_qdout20_OBUFT : X_TRI
    port map (
      I => MD_20_OUTMUX,
      CTL => MD_20_ENABLE,
      O => MD(20)
    );
  MD_20_ENABLEINV : X_INV
    port map (
      I => MD_20_TORGTS,
      O => MD_20_ENABLE
    );
  MD_20_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(20),
      O => MD_20_TORGTS
    );
  MD_20_OUTMUX_241 : X_BUF
    port map (
      I => memcontroller_dnout(20),
      O => MD_20_OUTMUX
    );
  MD_20_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(20),
      O => MD_20_OD
    );
  memcontroller_qdout20_IBUF : X_BUF
    port map (
      I => MD(20),
      O => memcontroller_q(20)
    );
  memcontroller_qdout12_OBUFT : X_TRI
    port map (
      I => MD_12_OUTMUX,
      CTL => MD_12_ENABLE,
      O => MD(12)
    );
  MD_12_ENABLEINV : X_INV
    port map (
      I => MD_12_TORGTS,
      O => MD_12_ENABLE
    );
  MD_12_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(12),
      O => MD_12_TORGTS
    );
  MD_12_OUTMUX_242 : X_BUF
    port map (
      I => memcontroller_dnout(12),
      O => MD_12_OUTMUX
    );
  MD_12_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(12),
      O => MD_12_OD
    );
  memcontroller_qdout12_IBUF : X_BUF
    port map (
      I => MD(12),
      O => memcontroller_q(12)
    );
  memcontroller_qdout21_OBUFT : X_TRI
    port map (
      I => MD_21_OUTMUX,
      CTL => MD_21_ENABLE,
      O => MD(21)
    );
  MD_21_ENABLEINV : X_INV
    port map (
      I => MD_21_TORGTS,
      O => MD_21_ENABLE
    );
  MD_21_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(21),
      O => MD_21_TORGTS
    );
  MD_21_OUTMUX_243 : X_BUF
    port map (
      I => memcontroller_dnout(21),
      O => MD_21_OUTMUX
    );
  MD_21_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(21),
      O => MD_21_OD
    );
  memcontroller_qdout21_IBUF : X_BUF
    port map (
      I => MD(21),
      O => memcontroller_q(21)
    );
  memcontroller_qdout13_OBUFT : X_TRI
    port map (
      I => MD_13_OUTMUX,
      CTL => MD_13_ENABLE,
      O => MD(13)
    );
  MD_13_ENABLEINV : X_INV
    port map (
      I => MD_13_TORGTS,
      O => MD_13_ENABLE
    );
  MD_13_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(13),
      O => MD_13_TORGTS
    );
  MD_13_OUTMUX_244 : X_BUF
    port map (
      I => memcontroller_dnout(13),
      O => MD_13_OUTMUX
    );
  MD_13_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(13),
      O => MD_13_OD
    );
  memcontroller_qdout13_IBUF : X_BUF
    port map (
      I => MD(13),
      O => memcontroller_q(13)
    );
  memcontroller_qdout22_OBUFT : X_TRI
    port map (
      I => MD_22_OUTMUX,
      CTL => MD_22_ENABLE,
      O => MD(22)
    );
  MD_22_ENABLEINV : X_INV
    port map (
      I => MD_22_TORGTS,
      O => MD_22_ENABLE
    );
  MD_22_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(22),
      O => MD_22_TORGTS
    );
  MD_22_OUTMUX_245 : X_BUF
    port map (
      I => memcontroller_dnout(22),
      O => MD_22_OUTMUX
    );
  MD_22_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(22),
      O => MD_22_OD
    );
  memcontroller_qdout22_IBUF : X_BUF
    port map (
      I => MD(22),
      O => memcontroller_q(22)
    );
  memcontroller_qdout14_OBUFT : X_TRI
    port map (
      I => MD_14_OUTMUX,
      CTL => MD_14_ENABLE,
      O => MD(14)
    );
  MD_14_ENABLEINV : X_INV
    port map (
      I => MD_14_TORGTS,
      O => MD_14_ENABLE
    );
  MD_14_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(14),
      O => MD_14_TORGTS
    );
  MD_14_OUTMUX_246 : X_BUF
    port map (
      I => memcontroller_dnout(14),
      O => MD_14_OUTMUX
    );
  MD_14_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(14),
      O => MD_14_OD
    );
  memcontroller_qdout14_IBUF : X_BUF
    port map (
      I => MD(14),
      O => memcontroller_q(14)
    );
  memcontroller_qdout30_OBUFT : X_TRI
    port map (
      I => MD_30_OUTMUX,
      CTL => MD_30_ENABLE,
      O => MD(30)
    );
  MD_30_ENABLEINV : X_INV
    port map (
      I => MD_30_TORGTS,
      O => MD_30_ENABLE
    );
  MD_30_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(30),
      O => MD_30_TORGTS
    );
  MD_30_OUTMUX_247 : X_BUF
    port map (
      I => memcontroller_dnout(30),
      O => MD_30_OUTMUX
    );
  MD_30_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(30),
      O => MD_30_OD
    );
  memcontroller_qdout30_IBUF : X_BUF
    port map (
      I => MD(30),
      O => memcontroller_q(30)
    );
  memcontroller_qdout23_OBUFT : X_TRI
    port map (
      I => MD_23_OUTMUX,
      CTL => MD_23_ENABLE,
      O => MD(23)
    );
  MD_23_ENABLEINV : X_INV
    port map (
      I => MD_23_TORGTS,
      O => MD_23_ENABLE
    );
  MD_23_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(23),
      O => MD_23_TORGTS
    );
  MD_23_OUTMUX_248 : X_BUF
    port map (
      I => memcontroller_dnout(23),
      O => MD_23_OUTMUX
    );
  MD_23_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(23),
      O => MD_23_OD
    );
  memcontroller_qdout23_IBUF : X_BUF
    port map (
      I => MD(23),
      O => memcontroller_q(23)
    );
  memcontroller_qdout15_OBUFT : X_TRI
    port map (
      I => MD_15_OUTMUX,
      CTL => MD_15_ENABLE,
      O => MD(15)
    );
  MD_15_ENABLEINV : X_INV
    port map (
      I => MD_15_TORGTS,
      O => MD_15_ENABLE
    );
  MD_15_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(15),
      O => MD_15_TORGTS
    );
  MD_15_OUTMUX_249 : X_BUF
    port map (
      I => memcontroller_dnout(15),
      O => MD_15_OUTMUX
    );
  MD_15_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(15),
      O => MD_15_OD
    );
  memcontroller_qdout15_IBUF : X_BUF
    port map (
      I => MD(15),
      O => memcontroller_q(15)
    );
  MD_31_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_31_TFF_RST
    );
  memcontroller_ts_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_31_TFF_RST,
      O => memcontroller_ts(31)
    );
  MD_31_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_31_OFF_RST
    );
  memcontroller_dnout_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_31_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_31_OFF_RST,
      O => memcontroller_dnout(31)
    );
  memcontroller_qdout31_OBUFT : X_TRI
    port map (
      I => MD_31_OUTMUX,
      CTL => MD_31_ENABLE,
      O => MD(31)
    );
  MD_31_ENABLEINV : X_INV
    port map (
      I => MD_31_TORGTS,
      O => MD_31_ENABLE
    );
  MD_31_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(31),
      O => MD_31_TORGTS
    );
  MD_31_OUTMUX_250 : X_BUF
    port map (
      I => memcontroller_dnout(31),
      O => MD_31_OUTMUX
    );
  MD_31_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(31),
      O => MD_31_OD
    );
  memcontroller_qdout31_IBUF : X_BUF
    port map (
      I => MD(31),
      O => memcontroller_q(31)
    );
  MD_24_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_24_TFF_RST
    );
  memcontroller_ts_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_24_TFF_RST,
      O => memcontroller_ts(24)
    );
  MD_24_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_24_OFF_RST
    );
  memcontroller_dnout_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_24_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_24_OFF_RST,
      O => memcontroller_dnout(24)
    );
  MD_24_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_24_IFF_RST
    );
  memcontroller_qn_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(24),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_24_IFF_RST,
      O => memcontroller_qn(24)
    );
  memcontroller_qdout24_OBUFT : X_TRI
    port map (
      I => MD_24_OUTMUX,
      CTL => MD_24_ENABLE,
      O => MD(24)
    );
  MD_24_ENABLEINV : X_INV
    port map (
      I => MD_24_TORGTS,
      O => MD_24_ENABLE
    );
  MD_24_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(24),
      O => MD_24_TORGTS
    );
  MD_24_OUTMUX_251 : X_BUF
    port map (
      I => memcontroller_dnout(24),
      O => MD_24_OUTMUX
    );
  MD_24_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(24),
      O => MD_24_OD
    );
  memcontroller_qdout24_IBUF : X_BUF
    port map (
      I => MD(24),
      O => memcontroller_q(24)
    );
  MD_16_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_16_TFF_RST
    );
  memcontroller_ts_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_16_TFF_RST,
      O => memcontroller_ts(16)
    );
  MD_16_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_16_OFF_RST
    );
  memcontroller_dnout_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_16_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_16_OFF_RST,
      O => memcontroller_dnout(16)
    );
  MD_16_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_16_IFF_RST
    );
  memcontroller_qn_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(16),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_16_IFF_RST,
      O => memcontroller_qn(16)
    );
  memcontroller_qdout16_OBUFT : X_TRI
    port map (
      I => MD_16_OUTMUX,
      CTL => MD_16_ENABLE,
      O => MD(16)
    );
  MD_16_ENABLEINV : X_INV
    port map (
      I => MD_16_TORGTS,
      O => MD_16_ENABLE
    );
  MD_16_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(16),
      O => MD_16_TORGTS
    );
  MD_16_OUTMUX_252 : X_BUF
    port map (
      I => memcontroller_dnout(16),
      O => MD_16_OUTMUX
    );
  MD_16_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(16),
      O => MD_16_OD
    );
  memcontroller_qdout16_IBUF : X_BUF
    port map (
      I => MD(16),
      O => memcontroller_q(16)
    );
  rx_input_fifo_fifo_BU157 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3480,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2400_FFX_RST,
      O => rx_input_fifo_fifo_N2400
    );
  rx_input_fifo_fifo_N2400_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2400_FFX_RST
    );
  MD_17_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_17_TFF_RST
    );
  memcontroller_ts_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_17_TFF_RST,
      O => memcontroller_ts(17)
    );
  MD_17_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_17_OFF_RST
    );
  memcontroller_dnout_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_17_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_17_OFF_RST,
      O => memcontroller_dnout(17)
    );
  MD_17_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_17_IFF_RST
    );
  memcontroller_qn_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(17),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_17_IFF_RST,
      O => memcontroller_qn(17)
    );
  memcontroller_qdout17_OBUFT : X_TRI
    port map (
      I => MD_17_OUTMUX,
      CTL => MD_17_ENABLE,
      O => MD(17)
    );
  MD_17_ENABLEINV : X_INV
    port map (
      I => MD_17_TORGTS,
      O => MD_17_ENABLE
    );
  MD_17_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(17),
      O => MD_17_TORGTS
    );
  MD_17_OUTMUX_253 : X_BUF
    port map (
      I => memcontroller_dnout(17),
      O => MD_17_OUTMUX
    );
  MD_17_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(17),
      O => MD_17_OD
    );
  memcontroller_qdout17_IBUF : X_BUF
    port map (
      I => MD(17),
      O => memcontroller_q(17)
    );
  MD_25_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_25_TFF_RST
    );
  memcontroller_ts_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_25_TFF_RST,
      O => memcontroller_ts(25)
    );
  MD_25_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_25_OFF_RST
    );
  memcontroller_dnout_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_25_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_25_OFF_RST,
      O => memcontroller_dnout(25)
    );
  MD_25_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_25_IFF_RST
    );
  memcontroller_qn_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(25),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_25_IFF_RST,
      O => memcontroller_qn(25)
    );
  memcontroller_qdout25_OBUFT : X_TRI
    port map (
      I => MD_25_OUTMUX,
      CTL => MD_25_ENABLE,
      O => MD(25)
    );
  MD_25_ENABLEINV : X_INV
    port map (
      I => MD_25_TORGTS,
      O => MD_25_ENABLE
    );
  MD_25_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(25),
      O => MD_25_TORGTS
    );
  MD_25_OUTMUX_254 : X_BUF
    port map (
      I => memcontroller_dnout(25),
      O => MD_25_OUTMUX
    );
  MD_25_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(25),
      O => MD_25_OD
    );
  memcontroller_qdout25_IBUF : X_BUF
    port map (
      I => MD(25),
      O => memcontroller_q(25)
    );
  MD_18_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_18_TFF_RST
    );
  memcontroller_ts_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_18_TFF_RST,
      O => memcontroller_ts(18)
    );
  MD_18_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_18_OFF_RST
    );
  memcontroller_dnout_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_18_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_18_OFF_RST,
      O => memcontroller_dnout(18)
    );
  MD_18_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_18_IFF_RST
    );
  memcontroller_qn_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(18),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_18_IFF_RST,
      O => memcontroller_qn(18)
    );
  memcontroller_qdout18_OBUFT : X_TRI
    port map (
      I => MD_18_OUTMUX,
      CTL => MD_18_ENABLE,
      O => MD(18)
    );
  MD_18_ENABLEINV : X_INV
    port map (
      I => MD_18_TORGTS,
      O => MD_18_ENABLE
    );
  MD_18_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(18),
      O => MD_18_TORGTS
    );
  MD_18_OUTMUX_255 : X_BUF
    port map (
      I => memcontroller_dnout(18),
      O => MD_18_OUTMUX
    );
  MD_18_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(18),
      O => MD_18_OD
    );
  memcontroller_qdout18_IBUF : X_BUF
    port map (
      I => MD(18),
      O => memcontroller_q(18)
    );
  MD_26_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_26_IFF_RST
    );
  memcontroller_qn_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(26),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_26_IFF_RST,
      O => memcontroller_qn(26)
    );
  memcontroller_qdout26_OBUFT : X_TRI
    port map (
      I => MD_26_OUTMUX,
      CTL => MD_26_ENABLE,
      O => MD(26)
    );
  MD_26_ENABLEINV : X_INV
    port map (
      I => MD_26_TORGTS,
      O => MD_26_ENABLE
    );
  MD_26_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(26),
      O => MD_26_TORGTS
    );
  MD_26_OUTMUX_256 : X_BUF
    port map (
      I => memcontroller_dnout(26),
      O => MD_26_OUTMUX
    );
  MD_26_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(26),
      O => MD_26_OD
    );
  memcontroller_qdout26_IBUF : X_BUF
    port map (
      I => MD(26),
      O => memcontroller_q(26)
    );
  rx_input_fifo_fifo_BU202 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2481,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2500_FFY_RST,
      O => rx_input_fifo_fifo_N2501
    );
  rx_input_fifo_fifo_N2500_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2500_FFY_RST
    );
  memcontroller_qdout19_OBUFT : X_TRI
    port map (
      I => MD_19_OUTMUX,
      CTL => MD_19_ENABLE,
      O => MD(19)
    );
  MD_19_ENABLEINV : X_INV
    port map (
      I => MD_19_TORGTS,
      O => MD_19_ENABLE
    );
  MD_19_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(19),
      O => MD_19_TORGTS
    );
  MD_19_OUTMUX_257 : X_BUF
    port map (
      I => memcontroller_dnout(19),
      O => MD_19_OUTMUX
    );
  MD_19_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(19),
      O => MD_19_OD
    );
  memcontroller_qdout19_IBUF : X_BUF
    port map (
      I => MD(19),
      O => memcontroller_q(19)
    );
  memcontroller_qdout27_OBUFT : X_TRI
    port map (
      I => MD_27_OUTMUX,
      CTL => MD_27_ENABLE,
      O => MD(27)
    );
  MD_27_ENABLEINV : X_INV
    port map (
      I => MD_27_TORGTS,
      O => MD_27_ENABLE
    );
  MD_27_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(27),
      O => MD_27_TORGTS
    );
  MD_27_OUTMUX_258 : X_BUF
    port map (
      I => memcontroller_dnout(27),
      O => MD_27_OUTMUX
    );
  MD_27_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(27),
      O => MD_27_OD
    );
  memcontroller_qdout27_IBUF : X_BUF
    port map (
      I => MD(27),
      O => memcontroller_q(27)
    );
  memcontroller_qdout28_OBUFT : X_TRI
    port map (
      I => MD_28_OUTMUX,
      CTL => MD_28_ENABLE,
      O => MD(28)
    );
  MD_28_ENABLEINV : X_INV
    port map (
      I => MD_28_TORGTS,
      O => MD_28_ENABLE
    );
  MD_28_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(28),
      O => MD_28_TORGTS
    );
  MD_28_OUTMUX_259 : X_BUF
    port map (
      I => memcontroller_dnout(28),
      O => MD_28_OUTMUX
    );
  MD_28_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(28),
      O => MD_28_OD
    );
  memcontroller_qdout28_IBUF : X_BUF
    port map (
      I => MD(28),
      O => memcontroller_q(28)
    );
  memcontroller_qdout29_OBUFT : X_TRI
    port map (
      I => MD_29_OUTMUX,
      CTL => MD_29_ENABLE,
      O => MD(29)
    );
  MD_29_ENABLEINV : X_INV
    port map (
      I => MD_29_TORGTS,
      O => MD_29_ENABLE
    );
  MD_29_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(29),
      O => MD_29_TORGTS
    );
  MD_29_OUTMUX_260 : X_BUF
    port map (
      I => memcontroller_dnout(29),
      O => MD_29_OUTMUX
    );
  MD_29_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(29),
      O => MD_29_OD
    );
  memcontroller_qdout29_IBUF : X_BUF
    port map (
      I => MD(29),
      O => memcontroller_q(29)
    );
  LEDPOWER_LOGIC_ONE_261 : X_ONE
    port map (
      O => LEDPOWER_LOGIC_ONE
    );
  LEDPOWER_OBUF : X_TRI
    port map (
      I => LEDPOWER_OUTMUX,
      CTL => LEDPOWER_ENABLE,
      O => LEDPOWER
    );
  LEDPOWER_ENABLEINV : X_INV
    port map (
      I => LEDPOWER_TORGTS,
      O => LEDPOWER_ENABLE
    );
  LEDPOWER_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDPOWER_TORGTS
    );
  LEDPOWER_OUTMUX_262 : X_BUF
    port map (
      I => LEDPOWER_LOGIC_ONE,
      O => LEDPOWER_OUTMUX
    );
  memcontroller_MA_0_OBUF : X_TRI
    port map (
      I => MA_0_OUTMUX,
      CTL => MA_0_ENABLE,
      O => MA(0)
    );
  MA_0_ENABLEINV : X_INV
    port map (
      I => MA_0_TORGTS,
      O => MA_0_ENABLE
    );
  MA_0_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_0_TORGTS
    );
  MA_0_OUTMUX_263 : X_BUF
    port map (
      I => memcontroller_ADDREXT(0),
      O => MA_0_OUTMUX
    );
  MA_0_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_0_OCEMUXNOT
    );
  MA_0_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(0),
      O => MA_0_OD
    );
  memcontroller_MA_1_OBUF : X_TRI
    port map (
      I => MA_1_OUTMUX,
      CTL => MA_1_ENABLE,
      O => MA(1)
    );
  MA_1_ENABLEINV : X_INV
    port map (
      I => MA_1_TORGTS,
      O => MA_1_ENABLE
    );
  MA_1_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_1_TORGTS
    );
  MA_1_OUTMUX_264 : X_BUF
    port map (
      I => memcontroller_ADDREXT(1),
      O => MA_1_OUTMUX
    );
  MA_1_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_1_OCEMUXNOT
    );
  MA_1_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(1),
      O => MA_1_OD
    );
  memcontroller_MA_2_OBUF : X_TRI
    port map (
      I => MA_2_OUTMUX,
      CTL => MA_2_ENABLE,
      O => MA(2)
    );
  MA_2_ENABLEINV : X_INV
    port map (
      I => MA_2_TORGTS,
      O => MA_2_ENABLE
    );
  MA_2_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_2_TORGTS
    );
  MA_2_OUTMUX_265 : X_BUF
    port map (
      I => memcontroller_ADDREXT(2),
      O => MA_2_OUTMUX
    );
  MA_2_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_2_OCEMUXNOT
    );
  MA_2_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(2),
      O => MA_2_OD
    );
  rx_input_fifo_fifo_BU208 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2479,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2499_FFX_RST,
      O => rx_input_fifo_fifo_N2499
    );
  rx_input_fifo_fifo_N2499_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2499_FFX_RST
    );
  memcontroller_MA_3_OBUF : X_TRI
    port map (
      I => MA_3_OUTMUX,
      CTL => MA_3_ENABLE,
      O => MA(3)
    );
  MA_3_ENABLEINV : X_INV
    port map (
      I => MA_3_TORGTS,
      O => MA_3_ENABLE
    );
  MA_3_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_3_TORGTS
    );
  MA_3_OUTMUX_266 : X_BUF
    port map (
      I => memcontroller_ADDREXT(3),
      O => MA_3_OUTMUX
    );
  MA_3_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_3_OCEMUXNOT
    );
  MA_3_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(3),
      O => MA_3_OD
    );
  memcontroller_MA_4_OBUF : X_TRI
    port map (
      I => MA_4_OUTMUX,
      CTL => MA_4_ENABLE,
      O => MA(4)
    );
  MA_4_ENABLEINV : X_INV
    port map (
      I => MA_4_TORGTS,
      O => MA_4_ENABLE
    );
  MA_4_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_4_TORGTS
    );
  MA_4_OUTMUX_267 : X_BUF
    port map (
      I => memcontroller_ADDREXT(4),
      O => MA_4_OUTMUX
    );
  MA_4_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_4_OCEMUXNOT
    );
  MA_4_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(4),
      O => MA_4_OD
    );
  memcontroller_MA_5_OBUF : X_TRI
    port map (
      I => MA_5_OUTMUX,
      CTL => MA_5_ENABLE,
      O => MA(5)
    );
  MA_5_ENABLEINV : X_INV
    port map (
      I => MA_5_TORGTS,
      O => MA_5_ENABLE
    );
  MA_5_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_5_TORGTS
    );
  MA_5_OUTMUX_268 : X_BUF
    port map (
      I => memcontroller_ADDREXT(5),
      O => MA_5_OUTMUX
    );
  MA_5_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_5_OCEMUXNOT
    );
  MA_5_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(5),
      O => MA_5_OD
    );
  memcontroller_MA_6_OBUF : X_TRI
    port map (
      I => MA_6_OUTMUX,
      CTL => MA_6_ENABLE,
      O => MA(6)
    );
  MA_6_ENABLEINV : X_INV
    port map (
      I => MA_6_TORGTS,
      O => MA_6_ENABLE
    );
  MA_6_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_6_TORGTS
    );
  MA_6_OUTMUX_269 : X_BUF
    port map (
      I => memcontroller_ADDREXT(6),
      O => MA_6_OUTMUX
    );
  MA_6_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_6_OCEMUXNOT
    );
  MA_6_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(6),
      O => MA_6_OD
    );
  memcontroller_MA_7_OBUF : X_TRI
    port map (
      I => MA_7_OUTMUX,
      CTL => MA_7_ENABLE,
      O => MA(7)
    );
  MA_7_ENABLEINV : X_INV
    port map (
      I => MA_7_TORGTS,
      O => MA_7_ENABLE
    );
  MA_7_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_7_TORGTS
    );
  MA_7_OUTMUX_270 : X_BUF
    port map (
      I => memcontroller_ADDREXT(7),
      O => MA_7_OUTMUX
    );
  MA_7_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_7_OCEMUXNOT
    );
  MA_7_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(7),
      O => MA_7_OD
    );
  memcontroller_MA_8_OBUF : X_TRI
    port map (
      I => MA_8_OUTMUX,
      CTL => MA_8_ENABLE,
      O => MA(8)
    );
  MA_8_ENABLEINV : X_INV
    port map (
      I => MA_8_TORGTS,
      O => MA_8_ENABLE
    );
  MA_8_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_8_TORGTS
    );
  MA_8_OUTMUX_271 : X_BUF
    port map (
      I => memcontroller_ADDREXT(8),
      O => MA_8_OUTMUX
    );
  MA_8_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_8_OCEMUXNOT
    );
  MA_8_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(8),
      O => MA_8_OD
    );
  memcontroller_MA_9_OBUF : X_TRI
    port map (
      I => MA_9_OUTMUX,
      CTL => MA_9_ENABLE,
      O => MA(9)
    );
  MA_9_ENABLEINV : X_INV
    port map (
      I => MA_9_TORGTS,
      O => MA_9_ENABLE
    );
  MA_9_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_9_TORGTS
    );
  MA_9_OUTMUX_272 : X_BUF
    port map (
      I => memcontroller_ADDREXT(9),
      O => MA_9_OUTMUX
    );
  MA_9_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_9_OCEMUXNOT
    );
  MA_9_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(9),
      O => MA_9_OD
    );
  mac_control_PHYRESET_OBUF_273 : X_TRI
    port map (
      I => PHYRESET_OUTMUX,
      CTL => PHYRESET_ENABLE,
      O => PHYRESET
    );
  PHYRESET_ENABLEINV : X_INV
    port map (
      I => PHYRESET_TORGTS,
      O => PHYRESET_ENABLE
    );
  PHYRESET_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => PHYRESET_TORGTS
    );
  PHYRESET_OUTMUX_274 : X_BUF
    port map (
      I => mac_control_PHYRESET_OBUF,
      O => PHYRESET_OUTMUX
    );
  PHYRESET_OMUX : X_BUF
    port map (
      I => mac_control_N79380,
      O => PHYRESET_OD
    );
  memcontroller_qdout0_OBUFT : X_TRI
    port map (
      I => MD_0_OUTMUX,
      CTL => MD_0_ENABLE,
      O => MD(0)
    );
  MD_0_ENABLEINV : X_INV
    port map (
      I => MD_0_TORGTS,
      O => MD_0_ENABLE
    );
  MD_0_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_0_TORGTS
    );
  MD_0_OUTMUX_275 : X_BUF
    port map (
      I => memcontroller_dnout(0),
      O => MD_0_OUTMUX
    );
  MD_0_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(0),
      O => MD_0_OD
    );
  memcontroller_qdout0_IBUF : X_BUF
    port map (
      I => MD(0),
      O => memcontroller_q(0)
    );
  rx_input_fifo_fifo_BU95 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2812,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N15_FFY_RST,
      O => rx_input_fifo_fifo_N14
    );
  rx_input_fifo_fifo_N15_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N15_FFY_RST
    );
  memcontroller_qdout1_OBUFT : X_TRI
    port map (
      I => MD_1_OUTMUX,
      CTL => MD_1_ENABLE,
      O => MD(1)
    );
  MD_1_ENABLEINV : X_INV
    port map (
      I => MD_1_TORGTS,
      O => MD_1_ENABLE
    );
  MD_1_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(1),
      O => MD_1_TORGTS
    );
  MD_1_OUTMUX_276 : X_BUF
    port map (
      I => memcontroller_dnout(1),
      O => MD_1_OUTMUX
    );
  MD_1_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(1),
      O => MD_1_OD
    );
  memcontroller_qdout1_IBUF : X_BUF
    port map (
      I => MD(1),
      O => memcontroller_q(1)
    );
  memcontroller_qdout2_OBUFT : X_TRI
    port map (
      I => MD_2_OUTMUX,
      CTL => MD_2_ENABLE,
      O => MD(2)
    );
  MD_2_ENABLEINV : X_INV
    port map (
      I => MD_2_TORGTS,
      O => MD_2_ENABLE
    );
  MD_2_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(2),
      O => MD_2_TORGTS
    );
  MD_2_OUTMUX_277 : X_BUF
    port map (
      I => memcontroller_dnout(2),
      O => MD_2_OUTMUX
    );
  MD_2_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(2),
      O => MD_2_OD
    );
  memcontroller_qdout2_IBUF : X_BUF
    port map (
      I => MD(2),
      O => memcontroller_q(2)
    );
  memcontroller_qdout3_OBUFT : X_TRI
    port map (
      I => MD_3_OUTMUX,
      CTL => MD_3_ENABLE,
      O => MD(3)
    );
  MD_3_ENABLEINV : X_INV
    port map (
      I => MD_3_TORGTS,
      O => MD_3_ENABLE
    );
  MD_3_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(3),
      O => MD_3_TORGTS
    );
  MD_3_OUTMUX_278 : X_BUF
    port map (
      I => memcontroller_dnout(3),
      O => MD_3_OUTMUX
    );
  MD_3_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(3),
      O => MD_3_OD
    );
  memcontroller_qdout3_IBUF : X_BUF
    port map (
      I => MD(3),
      O => memcontroller_q(3)
    );
  memcontroller_qdout4_OBUFT : X_TRI
    port map (
      I => MD_4_OUTMUX,
      CTL => MD_4_ENABLE,
      O => MD(4)
    );
  MD_4_ENABLEINV : X_INV
    port map (
      I => MD_4_TORGTS,
      O => MD_4_ENABLE
    );
  MD_4_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(4),
      O => MD_4_TORGTS
    );
  MD_4_OUTMUX_279 : X_BUF
    port map (
      I => memcontroller_dnout(4),
      O => MD_4_OUTMUX
    );
  MD_4_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(4),
      O => MD_4_OD
    );
  memcontroller_qdout4_IBUF : X_BUF
    port map (
      I => MD(4),
      O => memcontroller_q(4)
    );
  memcontroller_qdout5_OBUFT : X_TRI
    port map (
      I => MD_5_OUTMUX,
      CTL => MD_5_ENABLE,
      O => MD(5)
    );
  MD_5_ENABLEINV : X_INV
    port map (
      I => MD_5_TORGTS,
      O => MD_5_ENABLE
    );
  MD_5_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(5),
      O => MD_5_TORGTS
    );
  MD_5_OUTMUX_280 : X_BUF
    port map (
      I => memcontroller_dnout(5),
      O => MD_5_OUTMUX
    );
  MD_5_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(5),
      O => MD_5_OD
    );
  memcontroller_qdout5_IBUF : X_BUF
    port map (
      I => MD(5),
      O => memcontroller_q(5)
    );
  rx_input_fifo_control_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_control_cs_FFd3,
      ADR2 => VCC,
      ADR3 => rx_input_ce,
      O => rx_input_fifo_control_cs_FFd2_In
    );
  rx_input_fifo_control_cs_FFd1_In1 : X_LUT4
    generic map(
      INIT => X"FC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_control_cs_FFd1,
      ADR2 => rx_input_fifo_control_cs_FFd2,
      ADR3 => rx_input_ce,
      O => rx_input_fifo_control_cs_FFd1_In
    );
  rx_input_fifo_control_cs_FFd4_In_281 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_ce,
      ADR3 => rx_input_fifo_control_cs_FFd4_In_2,
      O => rx_input_fifo_control_cs_FFd4_In
    );
  rx_input_fifo_control_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd4,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_ce,
      O => rx_input_fifo_control_cs_FFd3_In
    );
  rx_output_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => rx_output_cs_FFd3,
      ADR1 => rx_output_nf,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_cs_FFd2_In
    );
  rx_output_cs_FFd1_In1 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_nf,
      ADR2 => rx_output_cs_FFd2,
      ADR3 => VCC,
      O => rx_output_cs_FFd1_In
    );
  mac_control_lmacaddr_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_23_FFX_RST,
      O => mac_control_lmacaddr(23)
    );
  mac_control_lmacaddr_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_23_FFX_RST
    );
  rx_output_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"C888"
    )
    port map (
      ADR0 => rx_output_cs_FFd4,
      ADR1 => rx_output_nf,
      ADR2 => rx_output_cs_FFd5,
      ADR3 => rx_output_n0018,
      O => rx_output_cs_FFd4_In
    );
  rx_output_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => rx_output_nf,
      ADR1 => rx_output_fifo_nearfull,
      ADR2 => rx_output_cs_FFd6,
      ADR3 => clken3,
      O => rx_output_cs_FFd3_In
    );
  rx_output_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => rx_output_nf,
      ADR1 => VCC,
      ADR2 => rx_output_cs_FFd9,
      ADR3 => VCC,
      O => rx_output_cs_FFd8_In
    );
  rx_output_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => rx_output_nf,
      ADR1 => VCC,
      ADR2 => rx_output_cs_FFd8,
      ADR3 => VCC,
      O => rx_output_cs_FFd7_In
    );
  tx_input_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_fifofulll,
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd5,
      O => tx_input_cs_FFd2_In
    );
  tx_input_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => tx_input_fifofulll,
      ADR1 => VCC,
      ADR2 => tx_input_cs_FFd5,
      ADR3 => VCC,
      O => tx_input_cs_FFd3_In
    );
  tx_input_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"CCC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_cs_FFd9,
      ADR2 => tx_input_N81681,
      ADR3 => tx_input_Ker34480137_2,
      O => tx_input_cs_FFd8_In
    );
  tx_input_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"4F44"
    )
    port map (
      ADR0 => tx_input_N73800,
      ADR1 => tx_input_cs_FFd9,
      ADR2 => tx_input_den,
      ADR3 => tx_input_cs_FFd7,
      O => tx_input_cs_FFd7_In
    );
  tx_input_cs_FFd9_In1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_den,
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd10,
      O => tx_input_cs_FFd9_In
    );
  rx_input_memio_Mshreg_lbpout4_10_srl_5 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_54,
      A1 => GLOBAL_LOGIC1_4,
      A2 => GLOBAL_LOGIC0_54,
      A3 => GLOBAL_LOGIC0_51,
      D => rx_input_memio_bp(10),
      CE => rx_input_memio_Mshreg_lbpout4_10_59_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_10_net14
    );
  rx_input_memio_Mshreg_lbpout4_10_59_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_10_59_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_10_59_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_10_59_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_11_srl_4 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_43,
      A1 => GLOBAL_LOGIC1_11,
      A2 => GLOBAL_LOGIC0_43,
      A3 => GLOBAL_LOGIC0_43,
      D => rx_input_memio_bp(11),
      CE => rx_input_memio_Mshreg_lbpout4_11_58_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_11_net12
    );
  rx_input_memio_Mshreg_lbpout4_11_58_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_11_58_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_11_58_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_11_58_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_12_srl_3 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_47,
      A1 => GLOBAL_LOGIC1_7,
      A2 => GLOBAL_LOGIC0_47,
      A3 => GLOBAL_LOGIC0_47,
      D => rx_input_memio_bp(12),
      CE => rx_input_memio_Mshreg_lbpout4_12_57_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_12_net10
    );
  rx_input_memio_Mshreg_lbpout4_12_57_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_12_57_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_12_57_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_12_57_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_13_srl_2 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_32,
      A1 => GLOBAL_LOGIC1_17,
      A2 => GLOBAL_LOGIC0_33,
      A3 => GLOBAL_LOGIC0_33,
      D => rx_input_memio_bp(13),
      CE => rx_input_memio_Mshreg_lbpout4_13_56_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_13_net8
    );
  rx_input_memio_Mshreg_lbpout4_13_56_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_13_56_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_13_56_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_13_56_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_14_srl_1 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_36,
      A1 => GLOBAL_LOGIC1_13,
      A2 => GLOBAL_LOGIC0_41,
      A3 => GLOBAL_LOGIC0_41,
      D => rx_input_memio_bp(14),
      CE => rx_input_memio_Mshreg_lbpout4_14_55_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_14_net6
    );
  rx_input_memio_Mshreg_lbpout4_14_55_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_14_55_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_14_55_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_14_55_SRMUX_OUTPUTNOT
    );
  mac_control_lmacaddr_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_31_FFX_RST,
      O => mac_control_lmacaddr(31)
    );
  mac_control_lmacaddr_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_31_FFX_RST
    );
  rx_input_memio_Mshreg_lbpout4_15_srl_0 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_36,
      A1 => GLOBAL_LOGIC1_16,
      A2 => GLOBAL_LOGIC0_36,
      A3 => GLOBAL_LOGIC0_36,
      D => rx_input_memio_bp(15),
      CE => rx_input_memio_Mshreg_lbpout4_15_54_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_15_net4
    );
  rx_input_memio_Mshreg_lbpout4_15_54_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_15_54_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_15_54_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_15_54_SRMUX_OUTPUTNOT
    );
  mac_control_Mshreg_sinlll_srl_16 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_27,
      A1 => GLOBAL_LOGIC0_3,
      A2 => GLOBAL_LOGIC0_3,
      A3 => GLOBAL_LOGIC0_3,
      D => SIN_IBUF,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      Q => mac_control_Mshreg_sinlll_net185
    );
  mac_control_n00571 : X_LUT4
    generic map(
      INIT => X"F7FF"
    )
    port map (
      ADR0 => mac_control_N52132,
      ADR1 => mac_control_N52236,
      ADR2 => mac_control_addr(7),
      ADR3 => mac_control_newcmd,
      O => mac_control_phyaddr_31_FROM
    );
  mac_control_PHY_status_n00171 : X_LUT4
    generic map(
      INIT => X"4050"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => mac_control_PHY_status_cs_FFd1,
      ADR2 => clkslen,
      ADR3 => mac_control_PHY_status_n0018,
      O => mac_control_phyaddr_31_GROM
    );
  mac_control_phyaddr_31_XUSED : X_BUF
    port map (
      I => mac_control_phyaddr_31_FROM,
      O => mac_control_PHY_status_n0018
    );
  mac_control_phyaddr_31_YUSED : X_BUF
    port map (
      I => mac_control_phyaddr_31_GROM,
      O => mac_control_PHY_status_n0017
    );
  rx_output_fifo_N1551_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1551_FFY_RST
    );
  rx_output_fifo_BU112 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2379,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1551_FFY_RST,
      O => rx_output_fifo_N1550
    );
  rx_output_fifo_BU104 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_fifo_N15,
      ADR1 => rx_output_fifo_N14,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N2339
    );
  rx_output_fifo_BU111 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_fifo_N14,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N13,
      O => rx_output_fifo_N2379
    );
  rx_output_fifo_BU118 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_fifo_N13,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N12,
      O => rx_output_fifo_N2419
    );
  rx_output_fifo_BU125 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_fifo_N11,
      ADR1 => rx_output_fifo_N12,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N2459
    );
  rx_output_fifo_BU265 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_fifo_N6,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N7,
      ADR3 => VCC,
      O => rx_output_fifo_N3267
    );
  rx_output_fifo_BU272 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_fifo_N6,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N5,
      ADR3 => VCC,
      O => rx_output_fifo_N3307
    );
  rx_output_fifo_BU251 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_fifo_N9,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N8,
      O => rx_output_fifo_N3187
    );
  rx_output_fifo_BU258 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N8,
      ADR2 => rx_output_fifo_N7,
      ADR3 => VCC,
      O => rx_output_fifo_N3227
    );
  rx_output_fifo_BU279 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_fifo_N5,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N4,
      ADR3 => VCC,
      O => rx_output_fifo_N3347
    );
  rx_output_fifo_BU286 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_fifo_N4,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N3,
      ADR3 => VCC,
      O => rx_output_fifo_N3387
    );
  rx_output_fifo_BU422 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_output_fifo_N1581,
      ADR1 => rx_output_fifo_N1579,
      ADR2 => rx_output_fifo_N1578,
      ADR3 => rx_output_fifo_N1580,
      O => rx_output_fifo_N1589_FROM
    );
  rx_output_fifo_BU428 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N1582,
      ADR3 => rx_output_fifo_N3959,
      O => rx_output_fifo_N3971
    );
  rx_output_fifo_N1589_XUSED : X_BUF
    port map (
      I => rx_output_fifo_N1589_FROM,
      O => rx_output_fifo_N3959
    );
  rx_output_fifo_BU416 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => rx_output_fifo_N1578,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N1580,
      ADR3 => rx_output_fifo_N1579,
      O => rx_output_fifo_N3973
    );
  rx_output_fifo_BU452 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_fifo_N3959,
      ADR1 => rx_output_fifo_N3958,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N3968
    );
  rx_output_fifo_BU440 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_output_fifo_N1583,
      ADR1 => rx_output_fifo_N3959,
      ADR2 => rx_output_fifo_N1582,
      ADR3 => rx_output_fifo_N1584,
      O => rx_output_fifo_N3969
    );
  mac_control_lmacaddr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_15_FFX_RST,
      O => mac_control_lmacaddr(15)
    );
  mac_control_lmacaddr_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_15_FFX_RST
    );
  tx_output_cs_FFd6_In1 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => tx_output_N73488,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_cs_FFd8,
      O => tx_output_cs_FFd6_In
    );
  tx_output_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => tx_output_N73488,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd6,
      ADR3 => VCC,
      O => tx_output_cs_FFd5_In
    );
  tx_output_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"AAEE"
    )
    port map (
      ADR0 => tx_output_cs_FFd9,
      ADR1 => tx_output_cs_FFd4,
      ADR2 => VCC,
      ADR3 => tx_output_N73488,
      O => tx_output_cs_FFd8_In
    );
  tx_output_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_decbcnt,
      ADR3 => tx_output_N73488,
      O => tx_output_cs_FFd7_In
    );
  rx_input_memio_Mshreg_lbpout4_0_srl_15 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_40,
      A1 => GLOBAL_LOGIC1_14,
      A2 => GLOBAL_LOGIC0_40,
      A3 => GLOBAL_LOGIC0_40,
      D => rx_input_memio_bp(0),
      CE => rx_input_memio_Mshreg_lbpout4_0_69_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_0_net34
    );
  rx_input_memio_Mshreg_lbpout4_0_69_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_0_69_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_0_69_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_0_69_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_1_srl_14 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_52,
      A1 => GLOBAL_LOGIC1_5,
      A2 => GLOBAL_LOGIC0_53,
      A3 => GLOBAL_LOGIC0_53,
      D => rx_input_memio_bp(1),
      CE => rx_input_memio_Mshreg_lbpout4_1_68_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_1_net32
    );
  rx_input_memio_Mshreg_lbpout4_1_68_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_1_68_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_1_68_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_1_68_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_2_srl_13 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_6,
      A1 => GLOBAL_LOGIC1_2,
      A2 => GLOBAL_LOGIC0,
      A3 => GLOBAL_LOGIC0_55,
      D => rx_input_memio_bp(2),
      CE => rx_input_memio_Mshreg_lbpout4_2_67_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_2_net30
    );
  rx_input_memio_Mshreg_lbpout4_2_67_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_2_67_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_2_67_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_2_67_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_3_srl_12 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_44,
      A1 => GLOBAL_LOGIC1_10,
      A2 => GLOBAL_LOGIC0_48,
      A3 => GLOBAL_LOGIC0_48,
      D => rx_input_memio_bp(3),
      CE => rx_input_memio_Mshreg_lbpout4_3_66_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_3_net28
    );
  rx_input_memio_Mshreg_lbpout4_3_66_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_3_66_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_3_66_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_3_66_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_4_srl_11 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_45,
      A1 => GLOBAL_LOGIC1_9,
      A2 => GLOBAL_LOGIC0_49,
      A3 => GLOBAL_LOGIC0_49,
      D => rx_input_memio_bp(4),
      CE => rx_input_memio_Mshreg_lbpout4_4_65_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_4_net26
    );
  rx_input_memio_Mshreg_lbpout4_4_65_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_4_65_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_4_65_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_4_65_SRMUX_OUTPUTNOT
    );
  memcontroller_qdout6_OBUFT : X_TRI
    port map (
      I => MD_6_OUTMUX,
      CTL => MD_6_ENABLE,
      O => MD(6)
    );
  MD_6_ENABLEINV : X_INV
    port map (
      I => MD_6_TORGTS,
      O => MD_6_ENABLE
    );
  MD_6_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(6),
      O => MD_6_TORGTS
    );
  MD_6_OUTMUX_282 : X_BUF
    port map (
      I => memcontroller_dnout(6),
      O => MD_6_OUTMUX
    );
  MD_6_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(6),
      O => MD_6_OD
    );
  memcontroller_qdout6_IBUF : X_BUF
    port map (
      I => MD(6),
      O => memcontroller_q(6)
    );
  memcontroller_qdout7_OBUFT : X_TRI
    port map (
      I => MD_7_OUTMUX,
      CTL => MD_7_ENABLE,
      O => MD(7)
    );
  MD_7_ENABLEINV : X_INV
    port map (
      I => MD_7_TORGTS,
      O => MD_7_ENABLE
    );
  MD_7_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(7),
      O => MD_7_TORGTS
    );
  MD_7_OUTMUX_283 : X_BUF
    port map (
      I => memcontroller_dnout(7),
      O => MD_7_OUTMUX
    );
  MD_7_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(7),
      O => MD_7_OD
    );
  memcontroller_qdout7_IBUF : X_BUF
    port map (
      I => MD(7),
      O => memcontroller_q(7)
    );
  memcontroller_qdout8_OBUFT : X_TRI
    port map (
      I => MD_8_OUTMUX,
      CTL => MD_8_ENABLE,
      O => MD(8)
    );
  MD_8_ENABLEINV : X_INV
    port map (
      I => MD_8_TORGTS,
      O => MD_8_ENABLE
    );
  MD_8_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(8),
      O => MD_8_TORGTS
    );
  MD_8_OUTMUX_284 : X_BUF
    port map (
      I => memcontroller_dnout(8),
      O => MD_8_OUTMUX
    );
  MD_8_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(8),
      O => MD_8_OD
    );
  memcontroller_qdout8_IBUF : X_BUF
    port map (
      I => MD(8),
      O => memcontroller_q(8)
    );
  memcontroller_qdout9_OBUFT : X_TRI
    port map (
      I => MD_9_OUTMUX,
      CTL => MD_9_ENABLE,
      O => MD(9)
    );
  MD_9_ENABLEINV : X_INV
    port map (
      I => MD_9_TORGTS,
      O => MD_9_ENABLE
    );
  MD_9_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(9),
      O => MD_9_TORGTS
    );
  MD_9_OUTMUX_285 : X_BUF
    port map (
      I => memcontroller_dnout(9),
      O => MD_9_OUTMUX
    );
  MD_9_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(9),
      O => MD_9_OD
    );
  memcontroller_qdout9_IBUF : X_BUF
    port map (
      I => MD(9),
      O => memcontroller_q(9)
    );
  GTX_CLK_OBUF_286 : X_TRI
    port map (
      I => GTX_CLK_OUTMUX,
      CTL => GTX_CLK_ENABLE,
      O => GTX_CLK
    );
  GTX_CLK_ENABLEINV : X_INV
    port map (
      I => GTX_CLK_TORGTS,
      O => GTX_CLK_ENABLE
    );
  GTX_CLK_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => GTX_CLK_TORGTS
    );
  GTX_CLK_OUTMUX_287 : X_BUF
    port map (
      I => GTX_CLK_OBUF,
      O => GTX_CLK_OUTMUX
    );
  clkio_dll : X_CLKDLLE
    generic map(
      CLKDV_DIVIDE => 2.0,
      DUTY_CYCLE_CORRECTION => TRUE,
      MAXPERCLKIN => 40000 ps
    )
    port map (
      CLKIN => CLKIOIN_IBUFG,
      CLKFB => clkio,
      RST => RESET_IBUF,
      CLK0 => clkio_to_bufg,
      CLK90 => clkio_dll_CLK90,
      CLK180 => clkio_dll_CLK180,
      CLK270 => clkio_dll_CLK270,
      CLK2X => clkio_dll_CLK2X,
      CLK2X180 => clkio_dll_CLK2X180,
      CLKDV => clkio_dll_CLKDV,
      LOCKED => clkio_dll_LOCKED
    );
  clk_dll : X_CLKDLLE
    generic map(
      CLKDV_DIVIDE => 2.0,
      DUTY_CYCLE_CORRECTION => TRUE,
      MAXPERCLKIN => 40000 ps
    )
    port map (
      CLKIN => CLKIN_IBUFG,
      CLKFB => GTX_CLK_OBUF,
      RST => RESET_IBUF,
      CLK0 => clk_to_bufg,
      CLK90 => MCLK_OBUF,
      CLK180 => clk_dll_CLK180,
      CLK270 => clk_dll_CLK270,
      CLK2X => clk_dll_CLK2X,
      CLK2X180 => clk_dll_CLK2X180,
      CLKDV => clk_dll_CLKDV,
      LOCKED => clk_dll_LOCKED
    );
  clkrx_dll : X_CLKDLLE
    generic map(
      CLKDV_DIVIDE => 2.0,
      DUTY_CYCLE_CORRECTION => TRUE,
      MAXPERCLKIN => 40000 ps
    )
    port map (
      CLKIN => RX_CLK_IBUFG,
      CLKFB => clkrx,
      RST => RESET_IBUF,
      CLK0 => clkrx_to_bufg,
      CLK90 => clkrx_dll_CLK90,
      CLK180 => clkrx_dll_CLK180,
      CLK270 => clkrx_dll_CLK270,
      CLK2X => clkrx_dll_CLK2X,
      CLK2X180 => clkrx_dll_CLK2X180,
      CLKDV => clkrx_dll_CLKDV,
      LOCKED => clkrx_dll_LOCKED
    );
  rx_input_fifo_fifo_B11_LOGIC_ONE_288 : X_ONE
    port map (
      O => rx_input_fifo_fifo_B11_LOGIC_ONE
    );
  rx_input_fifo_fifo_B11_LOGIC_ZERO_289 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_B11_LOGIC_ZERO
    );
  rx_input_fifo_fifo_B11 : X_RAMB4_S4_S4
    generic map(
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      SETUP_ALL => 3025 ps,
      XON => FALSE
    )
    port map (
      CLKA => clkrx,
      CLKB => GTX_CLK_OBUF,
      ENA => rx_input_fifo_fifo_B11_LOGIC_ONE,
      ENB => rx_input_fifo_fifo_N22,
      RSTA => rx_input_fifo_fifo_B11_LOGIC_ZERO,
      RSTB => rx_input_fifo_fifo_B11_LOGIC_ZERO,
      WEA => rx_input_fifo_fifo_N23,
      WEB => rx_input_fifo_fifo_B11_LOGIC_ZERO,
      GSR => GSR,
      ADDRA(9) => rx_input_fifo_fifo_N2,
      ADDRA(8) => rx_input_fifo_fifo_N3,
      ADDRA(7) => rx_input_fifo_fifo_N4,
      ADDRA(6) => rx_input_fifo_fifo_N5,
      ADDRA(5) => rx_input_fifo_fifo_N6,
      ADDRA(4) => rx_input_fifo_fifo_N7,
      ADDRA(3) => rx_input_fifo_fifo_N8,
      ADDRA(2) => rx_input_fifo_fifo_N9,
      ADDRA(1) => rx_input_fifo_fifo_N10,
      ADDRA(0) => rx_input_fifo_fifo_N11,
      ADDRB(9) => rx_input_fifo_fifo_N12,
      ADDRB(8) => rx_input_fifo_fifo_N13,
      ADDRB(7) => rx_input_fifo_fifo_N14,
      ADDRB(6) => rx_input_fifo_fifo_N15,
      ADDRB(5) => rx_input_fifo_fifo_N16,
      ADDRB(4) => rx_input_fifo_fifo_N17,
      ADDRB(3) => rx_input_fifo_fifo_N18,
      ADDRB(2) => rx_input_fifo_fifo_N19,
      ADDRB(1) => rx_input_fifo_fifo_N20,
      ADDRB(0) => rx_input_fifo_fifo_N21,
      DIA(3) => rx_input_fifoin(7),
      DIA(2) => rx_input_fifoin(6),
      DIA(1) => rx_input_fifoin(5),
      DIA(0) => rx_input_fifoin(4),
      DIB(3) => GLOBAL_LOGIC0_9,
      DIB(2) => GLOBAL_LOGIC0_9,
      DIB(1) => GLOBAL_LOGIC0_9,
      DIB(0) => GLOBAL_LOGIC0_9,
      DOA(3) => rx_input_fifo_fifo_B11_DOA3,
      DOA(2) => rx_input_fifo_fifo_B11_DOA2,
      DOA(1) => rx_input_fifo_fifo_B11_DOA1,
      DOA(0) => rx_input_fifo_fifo_B11_DOA0,
      DOB(3) => rx_input_fifo_fifodout(7),
      DOB(2) => rx_input_fifo_fifodout(6),
      DOB(1) => rx_input_fifo_fifodout(5),
      DOB(0) => rx_input_fifo_fifodout(4)
    );
  rx_input_fifo_fifo_B15_LOGIC_ONE_290 : X_ONE
    port map (
      O => rx_input_fifo_fifo_B15_LOGIC_ONE
    );
  rx_input_fifo_fifo_B15_LOGIC_ZERO_291 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_B15_LOGIC_ZERO
    );
  rx_input_fifo_fifo_B15 : X_RAMB4_S4_S4
    generic map(
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      SETUP_ALL => 3025 ps,
      XON => FALSE
    )
    port map (
      CLKA => clkrx,
      CLKB => GTX_CLK_OBUF,
      ENA => rx_input_fifo_fifo_B15_LOGIC_ONE,
      ENB => rx_input_fifo_fifo_N22,
      RSTA => rx_input_fifo_fifo_B15_LOGIC_ZERO,
      RSTB => rx_input_fifo_fifo_B15_LOGIC_ZERO,
      WEA => rx_input_fifo_fifo_N23,
      WEB => rx_input_fifo_fifo_B15_LOGIC_ZERO,
      GSR => GSR,
      ADDRA(9) => rx_input_fifo_fifo_N2,
      ADDRA(8) => rx_input_fifo_fifo_N3,
      ADDRA(7) => rx_input_fifo_fifo_N4,
      ADDRA(6) => rx_input_fifo_fifo_N5,
      ADDRA(5) => rx_input_fifo_fifo_N6,
      ADDRA(4) => rx_input_fifo_fifo_N7,
      ADDRA(3) => rx_input_fifo_fifo_N8,
      ADDRA(2) => rx_input_fifo_fifo_N9,
      ADDRA(1) => rx_input_fifo_fifo_N10,
      ADDRA(0) => rx_input_fifo_fifo_N11,
      ADDRB(9) => rx_input_fifo_fifo_N12,
      ADDRB(8) => rx_input_fifo_fifo_N13,
      ADDRB(7) => rx_input_fifo_fifo_N14,
      ADDRB(6) => rx_input_fifo_fifo_N15,
      ADDRB(5) => rx_input_fifo_fifo_N16,
      ADDRB(4) => rx_input_fifo_fifo_N17,
      ADDRB(3) => rx_input_fifo_fifo_N18,
      ADDRB(2) => rx_input_fifo_fifo_N19,
      ADDRB(1) => rx_input_fifo_fifo_N20,
      ADDRB(0) => rx_input_fifo_fifo_N21,
      DIA(3) => GLOBAL_LOGIC0_13,
      DIA(2) => GLOBAL_LOGIC0_11,
      DIA(1) => GLOBAL_LOGIC0_13,
      DIA(0) => rx_input_endfin,
      DIB(3) => GLOBAL_LOGIC0_13,
      DIB(2) => GLOBAL_LOGIC0_12,
      DIB(1) => GLOBAL_LOGIC0_13,
      DIB(0) => GLOBAL_LOGIC0_12,
      DOA(3) => rx_input_fifo_fifo_B15_DOA3,
      DOA(2) => rx_input_fifo_fifo_B15_DOA2,
      DOA(1) => rx_input_fifo_fifo_B15_DOA1,
      DOA(0) => rx_input_fifo_fifo_B15_DOA0,
      DOB(3) => rx_input_fifo_fifo_B15_DOB3,
      DOB(2) => rx_input_fifo_fifo_B15_DOB2,
      DOB(1) => rx_input_fifo_fifo_B15_DOB1,
      DOB(0) => rx_input_fifo_fifodout(8)
    );
  rx_input_fifo_fifo_B7_LOGIC_ONE_292 : X_ONE
    port map (
      O => rx_input_fifo_fifo_B7_LOGIC_ONE
    );
  rx_input_fifo_fifo_B7_LOGIC_ZERO_293 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_B7_LOGIC_ZERO
    );
  rx_input_fifo_fifo_B7 : X_RAMB4_S4_S4
    generic map(
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      SETUP_ALL => 3025 ps,
      XON => FALSE
    )
    port map (
      CLKA => clkrx,
      CLKB => GTX_CLK_OBUF,
      ENA => rx_input_fifo_fifo_B7_LOGIC_ONE,
      ENB => rx_input_fifo_fifo_N22,
      RSTA => rx_input_fifo_fifo_B7_LOGIC_ZERO,
      RSTB => rx_input_fifo_fifo_B7_LOGIC_ZERO,
      WEA => rx_input_fifo_fifo_N23,
      WEB => rx_input_fifo_fifo_B7_LOGIC_ZERO,
      GSR => GSR,
      ADDRA(9) => rx_input_fifo_fifo_N2,
      ADDRA(8) => rx_input_fifo_fifo_N3,
      ADDRA(7) => rx_input_fifo_fifo_N4,
      ADDRA(6) => rx_input_fifo_fifo_N5,
      ADDRA(5) => rx_input_fifo_fifo_N6,
      ADDRA(4) => rx_input_fifo_fifo_N7,
      ADDRA(3) => rx_input_fifo_fifo_N8,
      ADDRA(2) => rx_input_fifo_fifo_N9,
      ADDRA(1) => rx_input_fifo_fifo_N10,
      ADDRA(0) => rx_input_fifo_fifo_N11,
      ADDRB(9) => rx_input_fifo_fifo_N12,
      ADDRB(8) => rx_input_fifo_fifo_N13,
      ADDRB(7) => rx_input_fifo_fifo_N14,
      ADDRB(6) => rx_input_fifo_fifo_N15,
      ADDRB(5) => rx_input_fifo_fifo_N16,
      ADDRB(4) => rx_input_fifo_fifo_N17,
      ADDRB(3) => rx_input_fifo_fifo_N18,
      ADDRB(2) => rx_input_fifo_fifo_N19,
      ADDRB(1) => rx_input_fifo_fifo_N20,
      ADDRB(0) => rx_input_fifo_fifo_N21,
      DIA(3) => rx_input_fifoin(3),
      DIA(2) => rx_input_fifoin(2),
      DIA(1) => rx_input_fifoin(1),
      DIA(0) => rx_input_fifoin(0),
      DIB(3) => GLOBAL_LOGIC0_12,
      DIB(2) => GLOBAL_LOGIC0_12,
      DIB(1) => GLOBAL_LOGIC0_12,
      DIB(0) => GLOBAL_LOGIC0_12,
      DOA(3) => rx_input_fifo_fifo_B7_DOA3,
      DOA(2) => rx_input_fifo_fifo_B7_DOA2,
      DOA(1) => rx_input_fifo_fifo_B7_DOA1,
      DOA(0) => rx_input_fifo_fifo_B7_DOA0,
      DOB(3) => rx_input_fifo_fifodout(3),
      DOB(2) => rx_input_fifo_fifodout(2),
      DOB(1) => rx_input_fifo_fifodout(1),
      DOB(0) => rx_input_fifo_fifodout(0)
    );
  rx_output_fifo_B7_LOGIC_ONE_294 : X_ONE
    port map (
      O => rx_output_fifo_B7_LOGIC_ONE
    );
  rx_output_fifo_B7_LOGIC_ZERO_295 : X_ZERO
    port map (
      O => rx_output_fifo_B7_LOGIC_ZERO
    );
  rx_output_fifo_B7 : X_RAMB4_S16_S16
    generic map(
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      SETUP_ALL => 3025 ps,
      XON => FALSE
    )
    port map (
      CLKA => GTX_CLK_OBUF,
      CLKB => clkio,
      ENA => rx_output_fifo_B7_LOGIC_ONE,
      ENB => rx_output_fifo_N18,
      RSTA => rx_output_fifo_B7_LOGIC_ZERO,
      RSTB => rx_output_fifo_B7_LOGIC_ZERO,
      WEA => rx_output_fifo_N19,
      WEB => rx_output_fifo_B7_LOGIC_ZERO,
      GSR => GSR,
      ADDRA(7) => rx_output_fifo_N2,
      ADDRA(6) => rx_output_fifo_N3,
      ADDRA(5) => rx_output_fifo_N4,
      ADDRA(4) => rx_output_fifo_N5,
      ADDRA(3) => rx_output_fifo_N6,
      ADDRA(2) => rx_output_fifo_N7,
      ADDRA(1) => rx_output_fifo_N8,
      ADDRA(0) => rx_output_fifo_N9,
      ADDRB(7) => rx_output_fifo_N10,
      ADDRB(6) => rx_output_fifo_N11,
      ADDRB(5) => rx_output_fifo_N12,
      ADDRB(4) => rx_output_fifo_N13,
      ADDRB(3) => rx_output_fifo_N14,
      ADDRB(2) => rx_output_fifo_N15,
      ADDRB(1) => rx_output_fifo_N16,
      ADDRB(0) => rx_output_fifo_N17,
      DIA(15) => rx_output_fifodin(15),
      DIA(14) => rx_output_fifodin(14),
      DIA(13) => rx_output_fifodin(13),
      DIA(12) => rx_output_fifodin(12),
      DIA(11) => rx_output_fifodin(11),
      DIA(10) => rx_output_fifodin(10),
      DIA(9) => rx_output_fifodin(9),
      DIA(8) => rx_output_fifodin(8),
      DIA(7) => rx_output_fifodin(7),
      DIA(6) => rx_output_fifodin(6),
      DIA(5) => rx_output_fifodin(5),
      DIA(4) => rx_output_fifodin(4),
      DIA(3) => rx_output_fifodin(3),
      DIA(2) => rx_output_fifodin(2),
      DIA(1) => rx_output_fifodin(1),
      DIA(0) => rx_output_fifodin(0),
      DIB(15) => GLOBAL_LOGIC0_14,
      DIB(14) => GLOBAL_LOGIC0_14,
      DIB(13) => GLOBAL_LOGIC0_14,
      DIB(12) => GLOBAL_LOGIC0_14,
      DIB(11) => GLOBAL_LOGIC0_14,
      DIB(10) => GLOBAL_LOGIC0_14,
      DIB(9) => GLOBAL_LOGIC0_14,
      DIB(8) => GLOBAL_LOGIC0_14,
      DIB(7) => GLOBAL_LOGIC0_14,
      DIB(6) => GLOBAL_LOGIC0_14,
      DIB(5) => GLOBAL_LOGIC0_14,
      DIB(4) => GLOBAL_LOGIC0_14,
      DIB(3) => GLOBAL_LOGIC0_14,
      DIB(2) => GLOBAL_LOGIC0_14,
      DIB(1) => GLOBAL_LOGIC0_14,
      DIB(0) => GLOBAL_LOGIC0_14,
      DOA(15) => rx_output_fifo_B7_DOA15,
      DOA(14) => rx_output_fifo_B7_DOA14,
      DOA(13) => rx_output_fifo_B7_DOA13,
      DOA(12) => rx_output_fifo_B7_DOA12,
      DOA(11) => rx_output_fifo_B7_DOA11,
      DOA(10) => rx_output_fifo_B7_DOA10,
      DOA(9) => rx_output_fifo_B7_DOA9,
      DOA(8) => rx_output_fifo_B7_DOA8,
      DOA(7) => rx_output_fifo_B7_DOA7,
      DOA(6) => rx_output_fifo_B7_DOA6,
      DOA(5) => rx_output_fifo_B7_DOA5,
      DOA(4) => rx_output_fifo_B7_DOA4,
      DOA(3) => rx_output_fifo_B7_DOA3,
      DOA(2) => rx_output_fifo_B7_DOA2,
      DOA(1) => rx_output_fifo_B7_DOA1,
      DOA(0) => rx_output_fifo_B7_DOA0,
      DOB(15) => rx_output_fifodout(15),
      DOB(14) => rx_output_fifodout(14),
      DOB(13) => rx_output_fifodout(13),
      DOB(12) => rx_output_fifodout(12),
      DOB(11) => rx_output_fifodout(11),
      DOB(10) => rx_output_fifodout(10),
      DOB(9) => rx_output_fifodout(9),
      DOB(8) => rx_output_fifodout(8),
      DOB(7) => rx_output_fifodout(7),
      DOB(6) => rx_output_fifodout(6),
      DOB(5) => rx_output_fifodout(5),
      DOB(4) => rx_output_fifodout(4),
      DOB(3) => rx_output_fifodout(3),
      DOB(2) => rx_output_fifodout(2),
      DOB(1) => rx_output_fifodout(1),
      DOB(0) => rx_output_fifodout(0)
    );
  mac_control_Mmux_n0017_Result_31_38 : X_MUX2
    port map (
      IA => mac_control_N82509,
      IB => mac_control_N82511,
      SEL => mac_control_addr(1),
      O => mac_control_CHOICE1813_F5MUX
    );
  mac_control_Mmux_n0017_Result_31_38_G : X_LUT4
    generic map(
      INIT => X"8A80"
    )
    port map (
      ADR0 => mac_control_N52118,
      ADR1 => mac_control_txfifowerr_cnt(31),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_rxf_cnt(31),
      O => mac_control_N82511
    );
  mac_control_Mmux_n0017_Result_31_38_F : X_LUT4
    generic map(
      INIT => X"A000"
    )
    port map (
      ADR0 => mac_control_txf_cnt(31),
      ADR1 => VCC,
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_N52118,
      O => mac_control_N82509
    );
  mac_control_CHOICE1813_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1813_F5MUX,
      O => mac_control_CHOICE1813
    );
  mac_control_Mmux_n0017_Result_23_38 : X_MUX2
    port map (
      IA => mac_control_N82499,
      IB => mac_control_N82501,
      SEL => mac_control_addr(1),
      O => mac_control_CHOICE1869_F5MUX
    );
  mac_control_Mmux_n0017_Result_23_38_G : X_LUT4
    generic map(
      INIT => X"B080"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(23),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_rxf_cnt(23),
      O => mac_control_N82501
    );
  mac_control_Mmux_n0017_Result_23_38_F : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(23),
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_addr(0),
      O => mac_control_N82499
    );
  mac_control_CHOICE1869_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1869_F5MUX,
      O => mac_control_CHOICE1869
    );
  mac_control_Mmux_n0017_Result_19_38 : X_MUX2
    port map (
      IA => mac_control_N82504,
      IB => mac_control_N82506,
      SEL => mac_control_addr(1),
      O => mac_control_CHOICE1841_F5MUX
    );
  mac_control_Mmux_n0017_Result_19_38_G : X_LUT4
    generic map(
      INIT => X"E200"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(19),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_txfifowerr_cnt(19),
      ADR3 => mac_control_N52118,
      O => mac_control_N82506
    );
  mac_control_Mmux_n0017_Result_19_38_F : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_txf_cnt(19),
      ADR3 => mac_control_N52118,
      O => mac_control_N82504
    );
  mac_control_CHOICE1841_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1841_F5MUX,
      O => mac_control_CHOICE1841
    );
  mac_control_Mmux_n0017_Result_27_38 : X_MUX2
    port map (
      IA => mac_control_N82494,
      IB => mac_control_N82496,
      SEL => mac_control_addr(1),
      O => mac_control_CHOICE1897_F5MUX
    );
  mac_control_Mmux_n0017_Result_27_38_G : X_LUT4
    generic map(
      INIT => X"C0A0"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(27),
      ADR1 => mac_control_txfifowerr_cnt(27),
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_addr(0),
      O => mac_control_N82496
    );
  mac_control_Mmux_n0017_Result_27_38_F : X_LUT4
    generic map(
      INIT => X"A000"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(27),
      ADR3 => mac_control_N52118,
      O => mac_control_N82494
    );
  mac_control_CHOICE1897_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1897_F5MUX,
      O => mac_control_CHOICE1897
    );
  mac_control_PHY_status_MII_Interface_sout414 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_N82489,
      IB => mac_control_PHY_status_MII_Interface_N82491,
      SEL => mac_control_PHY_status_MII_Interface_statecnt(2),
      O => mac_control_PHY_status_MII_Interface_CHOICE2588_F5MUX
    );
  mac_control_PHY_status_MII_Interface_sout414_G : X_LUT4
    generic map(
      INIT => X"3000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR2 => mac_control_PHY_status_din(9),
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(4),
      O => mac_control_PHY_status_MII_Interface_N82491
    );
  mac_control_PHY_status_MII_Interface_sout414_F : X_LUT4
    generic map(
      INIT => X"0D01"
    )
    port map (
      ADR0 => mac_control_PHY_status_miirw,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR3 => mac_control_PHY_status_din(13),
      O => mac_control_PHY_status_MII_Interface_N82489
    );
  mac_control_PHY_status_MII_Interface_CHOICE2588_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2588_F5MUX,
      O => mac_control_PHY_status_MII_Interface_CHOICE2588
    );
  memcontroller_Mmux_addrn_inst_mux_f5_10111 : X_MUX2
    port map (
      IA => memcontroller_N82419,
      IB => memcontroller_N82421,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_10_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_10111_G : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(10),
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr4ext(10),
      O => memcontroller_N82421
    );
  memcontroller_Mmux_addrn_inst_mux_f5_10111_F : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => addr3ext(10),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr1ext(10),
      O => memcontroller_N82419
    );
  memcontroller_addrn_10_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_10_F5MUX,
      O => memcontroller_addrn(10)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_11111 : X_MUX2
    port map (
      IA => memcontroller_N82424,
      IB => memcontroller_N82426,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_11_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_11111_G : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(11),
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr4ext(11),
      O => memcontroller_N82426
    );
  memcontroller_Mmux_addrn_inst_mux_f5_11111_F : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => addr3ext(11),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr1ext(11),
      O => memcontroller_N82424
    );
  memcontroller_addrn_11_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_11_F5MUX,
      O => memcontroller_addrn(11)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_12111 : X_MUX2
    port map (
      IA => memcontroller_N82429,
      IB => memcontroller_N82431,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_12_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_12111_G : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => addr4ext(12),
      ADR1 => addr2ext(12),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82431
    );
  memcontroller_Mmux_addrn_inst_mux_f5_12111_F : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => addr1ext(12),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr3ext(12),
      O => memcontroller_N82429
    );
  memcontroller_addrn_12_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_12_F5MUX,
      O => memcontroller_addrn(12)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_13111 : X_MUX2
    port map (
      IA => memcontroller_N82434,
      IB => memcontroller_N82436,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_13_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_13111_G : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr4ext(13),
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr2ext(13),
      O => memcontroller_N82436
    );
  memcontroller_Mmux_addrn_inst_mux_f5_13111_F : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => addr3ext(13),
      ADR1 => addr1ext(13),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82434
    );
  memcontroller_addrn_13_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_13_F5MUX,
      O => memcontroller_addrn(13)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_14111 : X_MUX2
    port map (
      IA => memcontroller_N82439,
      IB => memcontroller_N82441,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_14_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_14111_G : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => addr4ext(14),
      ADR1 => addr2ext(14),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82441
    );
  memcontroller_Mmux_addrn_inst_mux_f5_14111_F : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(14),
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr1ext(14),
      O => memcontroller_N82439
    );
  memcontroller_addrn_14_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_14_F5MUX,
      O => memcontroller_addrn(14)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_15111 : X_MUX2
    port map (
      IA => memcontroller_N82444,
      IB => memcontroller_N82446,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_15_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_15111_G : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => addr4ext(15),
      ADR1 => addr2ext(15),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82446
    );
  memcontroller_Mmux_addrn_inst_mux_f5_15111_F : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => addr1ext(15),
      ADR1 => addr3ext(15),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82444
    );
  memcontroller_addrn_15_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_15_F5MUX,
      O => memcontroller_addrn(15)
    );
  rx_input_fifo_fifo_BU143 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3400,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2401_FFY_RST,
      O => rx_input_fifo_fifo_N2402
    );
  rx_input_fifo_fifo_N2401_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2401_FFY_RST
    );
  memcontroller_Mmux_addrn_inst_mux_f5_16111 : X_MUX2
    port map (
      IA => memcontroller_addrn_16_GROM,
      IB => memcontroller_addrn_16_FROM,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_16_F5MUX
    );
  memcontroller_addrn_16_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_addrn_16_FROM
    );
  memcontroller_addrn_16_G : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_addrn_16_GROM
    );
  memcontroller_addrn_16_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_16_F5MUX,
      O => memcontroller_addrn(16)
    );
  rx_input_fifo_fifo_BU89 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2811,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N15_FFX_RST,
      O => rx_input_fifo_fifo_N15
    );
  rx_input_fifo_fifo_N15_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N15_FFX_RST
    );
  memcontroller_Mmux_dn_inst_mux_f5_20111 : X_MUX2
    port map (
      IA => memcontroller_N82469,
      IB => memcontroller_N82471,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(3)
    );
  memcontroller_Mmux_dn_inst_mux_f5_20111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82471
    );
  memcontroller_Mmux_dn_inst_mux_f5_20111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => d1(3),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82469
    );
  memcontroller_dnl1_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_3_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_21111 : X_MUX2
    port map (
      IA => memcontroller_N82474,
      IB => memcontroller_N82476,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(4)
    );
  memcontroller_Mmux_dn_inst_mux_f5_21111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82476
    );
  memcontroller_Mmux_dn_inst_mux_f5_21111_F : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => d1(4),
      O => memcontroller_N82474
    );
  memcontroller_dnl1_4_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_4_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_22111 : X_MUX2
    port map (
      IA => memcontroller_N82479,
      IB => memcontroller_N82481,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(5)
    );
  memcontroller_Mmux_dn_inst_mux_f5_22111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82481
    );
  memcontroller_Mmux_dn_inst_mux_f5_22111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(5),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82479
    );
  memcontroller_dnl1_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_5_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_30111 : X_MUX2
    port map (
      IA => memcontroller_N82329,
      IB => memcontroller_N82331,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(13)
    );
  memcontroller_Mmux_dn_inst_mux_f5_30111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82331
    );
  memcontroller_Mmux_dn_inst_mux_f5_30111_F : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => d1(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82329
    );
  memcontroller_dnl1_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_13_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_31111 : X_MUX2
    port map (
      IA => memcontroller_N82324,
      IB => memcontroller_N82326,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(14)
    );
  memcontroller_Mmux_dn_inst_mux_f5_31111_G : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(14),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82326
    );
  memcontroller_Mmux_dn_inst_mux_f5_31111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(14),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82324
    );
  memcontroller_dnl1_14_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_14_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_23111 : X_MUX2
    port map (
      IA => memcontroller_N82484,
      IB => memcontroller_N82486,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(6)
    );
  memcontroller_Mmux_dn_inst_mux_f5_23111_G : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(6),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82486
    );
  memcontroller_Mmux_dn_inst_mux_f5_23111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => d1(6),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82484
    );
  memcontroller_dnl1_6_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_6_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_24111 : X_MUX2
    port map (
      IA => memcontroller_N82359,
      IB => memcontroller_N82361,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(7)
    );
  memcontroller_Mmux_dn_inst_mux_f5_24111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => d4(7),
      O => memcontroller_N82361
    );
  memcontroller_Mmux_dn_inst_mux_f5_24111_F : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(7),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82359
    );
  memcontroller_dnl1_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_7_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_32111 : X_MUX2
    port map (
      IA => memcontroller_N82319,
      IB => memcontroller_N82321,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(15)
    );
  memcontroller_Mmux_dn_inst_mux_f5_32111_G : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum(1),
      ADR2 => VCC,
      ADR3 => d4(15),
      O => memcontroller_N82321
    );
  memcontroller_Mmux_dn_inst_mux_f5_32111_F : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(15),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82319
    );
  memcontroller_dnl1_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_15_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_40111 : X_MUX2
    port map (
      IA => memcontroller_N82279,
      IB => memcontroller_N82281,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(23)
    );
  memcontroller_Mmux_dn_inst_mux_f5_40111_G : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(23),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82281
    );
  memcontroller_Mmux_dn_inst_mux_f5_40111_F : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(23),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82279
    );
  memcontroller_dnl1_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_23_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_17111 : X_MUX2
    port map (
      IA => memcontroller_N82454,
      IB => memcontroller_N82456,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(0)
    );
  memcontroller_Mmux_dn_inst_mux_f5_17111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82456
    );
  memcontroller_Mmux_dn_inst_mux_f5_17111_F : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(0),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82454
    );
  memcontroller_dnl1_0_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_0_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_25111 : X_MUX2
    port map (
      IA => memcontroller_N82354,
      IB => memcontroller_N82356,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(8)
    );
  memcontroller_Mmux_dn_inst_mux_f5_25111_G : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => d4(8),
      ADR1 => memcontroller_clknum(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N82356
    );
  memcontroller_Mmux_dn_inst_mux_f5_25111_F : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(8),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82354
    );
  memcontroller_dnl1_8_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_8_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_33111 : X_MUX2
    port map (
      IA => memcontroller_N82314,
      IB => memcontroller_N82316,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(16)
    );
  memcontroller_Mmux_dn_inst_mux_f5_33111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d4(16),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82316
    );
  memcontroller_Mmux_dn_inst_mux_f5_33111_F : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(16),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82314
    );
  memcontroller_dnl1_16_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_16_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_41111 : X_MUX2
    port map (
      IA => memcontroller_N82274,
      IB => memcontroller_N82276,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(24)
    );
  memcontroller_Mmux_dn_inst_mux_f5_41111_G : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => d4(24),
      ADR1 => memcontroller_clknum(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N82276
    );
  memcontroller_Mmux_dn_inst_mux_f5_41111_F : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum(1),
      ADR2 => d1(24),
      ADR3 => VCC,
      O => memcontroller_N82274
    );
  memcontroller_dnl1_24_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_24_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_18111 : X_MUX2
    port map (
      IA => memcontroller_N82459,
      IB => memcontroller_N82461,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(1)
    );
  memcontroller_Mmux_dn_inst_mux_f5_18111_G : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(1),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82461
    );
  memcontroller_Mmux_dn_inst_mux_f5_18111_F : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => d1(1),
      O => memcontroller_N82459
    );
  memcontroller_dnl1_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_1_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_26111 : X_MUX2
    port map (
      IA => memcontroller_N82349,
      IB => memcontroller_N82351,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(9)
    );
  memcontroller_Mmux_dn_inst_mux_f5_26111_G : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(9),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82351
    );
  memcontroller_Mmux_dn_inst_mux_f5_26111_F : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(9),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82349
    );
  memcontroller_dnl1_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_9_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_34111 : X_MUX2
    port map (
      IA => memcontroller_N82309,
      IB => memcontroller_N82311,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(17)
    );
  memcontroller_Mmux_dn_inst_mux_f5_34111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(17),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82311
    );
  memcontroller_Mmux_dn_inst_mux_f5_34111_F : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => d1(17),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82309
    );
  memcontroller_dnl1_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_17_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_42111 : X_MUX2
    port map (
      IA => memcontroller_N82269,
      IB => memcontroller_N82271,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(25)
    );
  memcontroller_Mmux_dn_inst_mux_f5_42111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => d4(25),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82271
    );
  memcontroller_Mmux_dn_inst_mux_f5_42111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(25),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82269
    );
  memcontroller_dnl1_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_25_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_19111 : X_MUX2
    port map (
      IA => memcontroller_N82464,
      IB => memcontroller_N82466,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(2)
    );
  memcontroller_Mmux_dn_inst_mux_f5_19111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => d4(2),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82466
    );
  memcontroller_Mmux_dn_inst_mux_f5_19111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => d1(2),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82464
    );
  memcontroller_dnl1_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_2_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_27111 : X_MUX2
    port map (
      IA => memcontroller_N82344,
      IB => memcontroller_N82346,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(10)
    );
  memcontroller_Mmux_dn_inst_mux_f5_27111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => d4(10),
      O => memcontroller_N82346
    );
  memcontroller_Mmux_dn_inst_mux_f5_27111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(10),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82344
    );
  memcontroller_dnl1_10_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_10_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_35111 : X_MUX2
    port map (
      IA => memcontroller_N82304,
      IB => memcontroller_N82306,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(18)
    );
  memcontroller_Mmux_dn_inst_mux_f5_35111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(18),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82306
    );
  memcontroller_Mmux_dn_inst_mux_f5_35111_F : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(18),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82304
    );
  memcontroller_dnl1_18_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_18_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_43111 : X_MUX2
    port map (
      IA => memcontroller_N82264,
      IB => memcontroller_N82266,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(26)
    );
  memcontroller_Mmux_dn_inst_mux_f5_43111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => d4(26),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82266
    );
  memcontroller_Mmux_dn_inst_mux_f5_43111_F : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(26),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82264
    );
  memcontroller_dnl1_26_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_26_CEMUXNOT
    );
  rx_input_fifo_fifo_BU83 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2810,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N17_FFY_RST,
      O => rx_input_fifo_fifo_N16
    );
  rx_input_fifo_fifo_N17_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N17_FFY_RST
    );
  memcontroller_Mmux_dn_inst_mux_f5_28111 : X_MUX2
    port map (
      IA => memcontroller_N82339,
      IB => memcontroller_N82341,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(11)
    );
  memcontroller_Mmux_dn_inst_mux_f5_28111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => d4(11),
      O => memcontroller_N82341
    );
  memcontroller_Mmux_dn_inst_mux_f5_28111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => d1(11),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82339
    );
  memcontroller_dnl1_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_11_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_36111 : X_MUX2
    port map (
      IA => memcontroller_N82299,
      IB => memcontroller_N82301,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(19)
    );
  memcontroller_Mmux_dn_inst_mux_f5_36111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => d4(19),
      O => memcontroller_N82301
    );
  memcontroller_Mmux_dn_inst_mux_f5_36111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => d1(19),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82299
    );
  memcontroller_dnl1_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_19_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_44111 : X_MUX2
    port map (
      IA => memcontroller_N82259,
      IB => memcontroller_N82261,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(27)
    );
  memcontroller_Mmux_dn_inst_mux_f5_44111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => d4(27),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82261
    );
  memcontroller_Mmux_dn_inst_mux_f5_44111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => d1(27),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82259
    );
  memcontroller_dnl1_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_27_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_29111 : X_MUX2
    port map (
      IA => memcontroller_N82334,
      IB => memcontroller_N82336,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(12)
    );
  memcontroller_Mmux_dn_inst_mux_f5_29111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(12),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82336
    );
  memcontroller_Mmux_dn_inst_mux_f5_29111_F : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => d1(12),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82334
    );
  memcontroller_dnl1_12_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_12_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_37111 : X_MUX2
    port map (
      IA => memcontroller_N82294,
      IB => memcontroller_N82296,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(20)
    );
  memcontroller_Mmux_dn_inst_mux_f5_37111_G : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(20),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82296
    );
  memcontroller_Mmux_dn_inst_mux_f5_37111_F : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => d1(20),
      O => memcontroller_N82294
    );
  memcontroller_dnl1_20_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_20_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_45111 : X_MUX2
    port map (
      IA => memcontroller_N82249,
      IB => memcontroller_N82251,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(28)
    );
  memcontroller_Mmux_dn_inst_mux_f5_45111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => d4(28),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82251
    );
  memcontroller_Mmux_dn_inst_mux_f5_45111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => d1(28),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82249
    );
  memcontroller_dnl1_28_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_28_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_38111 : X_MUX2
    port map (
      IA => memcontroller_N82289,
      IB => memcontroller_N82291,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(21)
    );
  memcontroller_Mmux_dn_inst_mux_f5_38111_G : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => d4(21),
      ADR1 => memcontroller_clknum(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N82291
    );
  memcontroller_Mmux_dn_inst_mux_f5_38111_F : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => memcontroller_clknum(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(21),
      O => memcontroller_N82289
    );
  memcontroller_dnl1_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_21_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_46111 : X_MUX2
    port map (
      IA => memcontroller_N82244,
      IB => memcontroller_N82246,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(29)
    );
  memcontroller_Mmux_dn_inst_mux_f5_46111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => d4(29),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82246
    );
  memcontroller_Mmux_dn_inst_mux_f5_46111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => d1(29),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82244
    );
  memcontroller_dnl1_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_29_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_39111 : X_MUX2
    port map (
      IA => memcontroller_N82284,
      IB => memcontroller_N82286,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(22)
    );
  memcontroller_Mmux_dn_inst_mux_f5_39111_G : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(22),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82286
    );
  memcontroller_Mmux_dn_inst_mux_f5_39111_F : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(22),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82284
    );
  memcontroller_dnl1_22_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_22_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_47111 : X_MUX2
    port map (
      IA => memcontroller_N82254,
      IB => memcontroller_N82256,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(30)
    );
  memcontroller_Mmux_dn_inst_mux_f5_47111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d4(30),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82256
    );
  memcontroller_Mmux_dn_inst_mux_f5_47111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => d1(30),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82254
    );
  memcontroller_dnl1_30_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_30_CEMUXNOT
    );
  rx_input_fifo_fifo_BU205 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2480,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2500_FFX_RST,
      O => rx_input_fifo_fifo_N2500
    );
  rx_input_fifo_fifo_N2500_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2500_FFX_RST
    );
  memcontroller_Mmux_dn_inst_mux_f5_48111 : X_MUX2
    port map (
      IA => memcontroller_N82449,
      IB => memcontroller_N82451,
      SEL => memcontroller_clknum(0),
      O => memcontroller_dn(31)
    );
  memcontroller_Mmux_dn_inst_mux_f5_48111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => d4(31),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82451
    );
  memcontroller_Mmux_dn_inst_mux_f5_48111_F : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => d1(31),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82449
    );
  memcontroller_dnl1_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_31_CEMUXNOT
    );
  memcontroller_Mmux_addrn_inst_mux_f5_0111 : X_MUX2
    port map (
      IA => memcontroller_N82369,
      IB => memcontroller_N82371,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_0_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_0111_G : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => addr4ext(0),
      ADR1 => addr2ext(0),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82371
    );
  memcontroller_Mmux_addrn_inst_mux_f5_0111_F : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => addr1ext(0),
      ADR1 => VCC,
      ADR2 => addr3ext(0),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82369
    );
  memcontroller_addrn_0_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_0_F5MUX,
      O => memcontroller_addrn(0)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_2111 : X_MUX2
    port map (
      IA => memcontroller_N82379,
      IB => memcontroller_N82381,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_2_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_2111_G : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => addr4ext(2),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr2ext(2),
      O => memcontroller_N82381
    );
  memcontroller_Mmux_addrn_inst_mux_f5_2111_F : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => addr1ext(2),
      ADR1 => addr3ext(2),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82379
    );
  memcontroller_addrn_2_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_2_F5MUX,
      O => memcontroller_addrn(2)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_3111 : X_MUX2
    port map (
      IA => memcontroller_N82384,
      IB => memcontroller_N82386,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_3_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_3111_G : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => addr4ext(3),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr2ext(3),
      O => memcontroller_N82386
    );
  memcontroller_Mmux_addrn_inst_mux_f5_3111_F : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => addr1ext(3),
      ADR1 => addr3ext(3),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82384
    );
  memcontroller_addrn_3_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_3_F5MUX,
      O => memcontroller_addrn(3)
    );
  rx_input_fifo_fifo_BU150 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3440,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2401_FFX_RST,
      O => rx_input_fifo_fifo_N2401
    );
  rx_input_fifo_fifo_N2401_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2401_FFX_RST
    );
  memcontroller_Mmux_addrn_inst_mux_f5_4111 : X_MUX2
    port map (
      IA => memcontroller_N82389,
      IB => memcontroller_N82391,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_4_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_4111_G : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => addr2ext(4),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr4ext(4),
      O => memcontroller_N82391
    );
  memcontroller_Mmux_addrn_inst_mux_f5_4111_F : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => addr3ext(4),
      ADR1 => addr1ext(4),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82389
    );
  memcontroller_addrn_4_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_4_F5MUX,
      O => memcontroller_addrn(4)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_1711 : X_MUX2
    port map (
      IA => memcontroller_N82374,
      IB => memcontroller_N82376,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_1_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_1711_G : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => addr4ext(1),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr2ext(1),
      O => memcontroller_N82376
    );
  memcontroller_Mmux_addrn_inst_mux_f5_1711_F : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr1ext(1),
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr3ext(1),
      O => memcontroller_N82374
    );
  memcontroller_addrn_1_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_1_F5MUX,
      O => memcontroller_addrn(1)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_5111 : X_MUX2
    port map (
      IA => memcontroller_N82394,
      IB => memcontroller_N82396,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_5_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_5111_G : X_LUT4
    generic map(
      INIT => X"B8B8"
    )
    port map (
      ADR0 => addr4ext(5),
      ADR1 => memcontroller_clknum(1),
      ADR2 => addr2ext(5),
      ADR3 => VCC,
      O => memcontroller_N82396
    );
  memcontroller_Mmux_addrn_inst_mux_f5_5111_F : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(5),
      ADR2 => memcontroller_clknum(1),
      ADR3 => addr1ext(5),
      O => memcontroller_N82394
    );
  memcontroller_addrn_5_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_5_F5MUX,
      O => memcontroller_addrn(5)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_6111 : X_MUX2
    port map (
      IA => memcontroller_N82399,
      IB => memcontroller_N82401,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_6_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_6111_G : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => addr4ext(6),
      ADR1 => memcontroller_clknum(1),
      ADR2 => VCC,
      ADR3 => addr2ext(6),
      O => memcontroller_N82401
    );
  memcontroller_Mmux_addrn_inst_mux_f5_6111_F : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => addr3ext(6),
      ADR1 => memcontroller_clknum(1),
      ADR2 => VCC,
      ADR3 => addr1ext(6),
      O => memcontroller_N82399
    );
  memcontroller_addrn_6_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_6_F5MUX,
      O => memcontroller_addrn(6)
    );
  rx_input_fifo_fifo_BU196 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2483,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2502_FFY_RST,
      O => rx_input_fifo_fifo_N2503
    );
  rx_input_fifo_fifo_N2502_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2502_FFY_RST
    );
  memcontroller_Mmux_addrn_inst_mux_f5_7111 : X_MUX2
    port map (
      IA => memcontroller_N82404,
      IB => memcontroller_N82406,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_7_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_7111_G : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => addr2ext(7),
      ADR1 => addr4ext(7),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82406
    );
  memcontroller_Mmux_addrn_inst_mux_f5_7111_F : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => addr3ext(7),
      ADR1 => VCC,
      ADR2 => addr1ext(7),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82404
    );
  memcontroller_addrn_7_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_7_F5MUX,
      O => memcontroller_addrn(7)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_8111 : X_MUX2
    port map (
      IA => memcontroller_N82409,
      IB => memcontroller_N82411,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_8_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_8111_G : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => addr4ext(8),
      ADR1 => addr2ext(8),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82411
    );
  memcontroller_Mmux_addrn_inst_mux_f5_8111_F : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => addr3ext(8),
      ADR1 => addr1ext(8),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82409
    );
  memcontroller_addrn_8_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_8_F5MUX,
      O => memcontroller_addrn(8)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_9111 : X_MUX2
    port map (
      IA => memcontroller_N82414,
      IB => memcontroller_N82416,
      SEL => memcontroller_clknum(0),
      O => memcontroller_addrn_9_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_9111_G : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => addr2ext(9),
      ADR1 => VCC,
      ADR2 => addr4ext(9),
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_N82416
    );
  memcontroller_Mmux_addrn_inst_mux_f5_9111_F : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => addr3ext(9),
      ADR1 => addr1ext(9),
      ADR2 => memcontroller_clknum(1),
      ADR3 => VCC,
      O => memcontroller_N82414
    );
  memcontroller_addrn_9_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_9_F5MUX,
      O => memcontroller_addrn(9)
    );
  addr2ext_0_LOGIC_ZERO_296 : X_ZERO
    port map (
      O => addr2ext_0_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_0_297 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_6,
      IB => addr2ext_0_LOGIC_ZERO,
      SEL => tx_output_addr_Madd_n0000_inst_lut2_0,
      O => tx_output_addr_Madd_n0000_inst_cy_0
    );
  tx_output_addr_Madd_n0000_inst_lut2_01 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_6,
      ADR1 => addr2ext(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_output_addr_Madd_n0000_inst_lut2_0
    );
  addr2ext_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_50,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(1),
      O => addr2ext_0_GROM
    );
  addr2ext_0_COUTUSED : X_BUF
    port map (
      I => addr2ext_0_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_1
    );
  tx_output_addr_Madd_n0000_inst_cy_1_298 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_50,
      IB => tx_output_addr_Madd_n0000_inst_cy_0,
      SEL => addr2ext_0_GROM,
      O => addr2ext_0_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_1 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_0,
      I1 => addr2ext_0_GROM,
      O => tx_output_addr_n0000(1)
    );
  addr2ext_2_LOGIC_ZERO_299 : X_ZERO
    port map (
      O => addr2ext_2_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_2_300 : X_MUX2
    port map (
      IA => addr2ext_2_LOGIC_ZERO,
      IB => addr2ext_2_CYINIT,
      SEL => addr2ext_2_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_2
    );
  tx_output_addr_Madd_n0000_inst_sum_2 : X_XOR2
    port map (
      I0 => addr2ext_2_CYINIT,
      I1 => addr2ext_2_FROM,
      O => tx_output_addr_n0000(2)
    );
  addr2ext_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(2),
      O => addr2ext_2_FROM
    );
  addr2ext_2_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr2ext_2_GROM
    );
  addr2ext_2_COUTUSED : X_BUF
    port map (
      I => addr2ext_2_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_3
    );
  tx_output_addr_Madd_n0000_inst_cy_3_301 : X_MUX2
    port map (
      IA => addr2ext_2_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_2,
      SEL => addr2ext_2_GROM,
      O => addr2ext_2_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_3 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_2,
      I1 => addr2ext_2_GROM,
      O => tx_output_addr_n0000(3)
    );
  addr2ext_2_CYINIT_302 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_1,
      O => addr2ext_2_CYINIT
    );
  addr2ext_4_LOGIC_ZERO_303 : X_ZERO
    port map (
      O => addr2ext_4_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_4_304 : X_MUX2
    port map (
      IA => addr2ext_4_LOGIC_ZERO,
      IB => addr2ext_4_CYINIT,
      SEL => addr2ext_4_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_4
    );
  tx_output_addr_Madd_n0000_inst_sum_4 : X_XOR2
    port map (
      I0 => addr2ext_4_CYINIT,
      I1 => addr2ext_4_FROM,
      O => tx_output_addr_n0000(4)
    );
  addr2ext_4_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => addr2ext(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr2ext_4_FROM
    );
  addr2ext_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr2ext(5),
      ADR3 => VCC,
      O => addr2ext_4_GROM
    );
  addr2ext_4_COUTUSED : X_BUF
    port map (
      I => addr2ext_4_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_5
    );
  tx_output_addr_Madd_n0000_inst_cy_5_305 : X_MUX2
    port map (
      IA => addr2ext_4_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_4,
      SEL => addr2ext_4_GROM,
      O => addr2ext_4_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_5 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_4,
      I1 => addr2ext_4_GROM,
      O => tx_output_addr_n0000(5)
    );
  addr2ext_4_CYINIT_306 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_3,
      O => addr2ext_4_CYINIT
    );
  addr2ext_6_LOGIC_ZERO_307 : X_ZERO
    port map (
      O => addr2ext_6_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_6_308 : X_MUX2
    port map (
      IA => addr2ext_6_LOGIC_ZERO,
      IB => addr2ext_6_CYINIT,
      SEL => addr2ext_6_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_6
    );
  tx_output_addr_Madd_n0000_inst_sum_6 : X_XOR2
    port map (
      I0 => addr2ext_6_CYINIT,
      I1 => addr2ext_6_FROM,
      O => tx_output_addr_n0000(6)
    );
  addr2ext_6_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr2ext(6),
      ADR3 => VCC,
      O => addr2ext_6_FROM
    );
  addr2ext_6_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(7),
      O => addr2ext_6_GROM
    );
  addr2ext_6_COUTUSED : X_BUF
    port map (
      I => addr2ext_6_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_7
    );
  tx_output_addr_Madd_n0000_inst_cy_7_309 : X_MUX2
    port map (
      IA => addr2ext_6_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_6,
      SEL => addr2ext_6_GROM,
      O => addr2ext_6_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_7 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_6,
      I1 => addr2ext_6_GROM,
      O => tx_output_addr_n0000(7)
    );
  addr2ext_6_CYINIT_310 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_5,
      O => addr2ext_6_CYINIT
    );
  addr2ext_8_LOGIC_ZERO_311 : X_ZERO
    port map (
      O => addr2ext_8_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_8_312 : X_MUX2
    port map (
      IA => addr2ext_8_LOGIC_ZERO,
      IB => addr2ext_8_CYINIT,
      SEL => addr2ext_8_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_8
    );
  tx_output_addr_Madd_n0000_inst_sum_8 : X_XOR2
    port map (
      I0 => addr2ext_8_CYINIT,
      I1 => addr2ext_8_FROM,
      O => tx_output_addr_n0000(8)
    );
  addr2ext_8_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr2ext_8_FROM
    );
  addr2ext_8_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(9),
      O => addr2ext_8_GROM
    );
  addr2ext_8_COUTUSED : X_BUF
    port map (
      I => addr2ext_8_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_9
    );
  tx_output_addr_Madd_n0000_inst_cy_9_313 : X_MUX2
    port map (
      IA => addr2ext_8_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_8,
      SEL => addr2ext_8_GROM,
      O => addr2ext_8_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_9 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_8,
      I1 => addr2ext_8_GROM,
      O => tx_output_addr_n0000(9)
    );
  addr2ext_8_CYINIT_314 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_7,
      O => addr2ext_8_CYINIT
    );
  addr2ext_10_LOGIC_ZERO_315 : X_ZERO
    port map (
      O => addr2ext_10_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_10_316 : X_MUX2
    port map (
      IA => addr2ext_10_LOGIC_ZERO,
      IB => addr2ext_10_CYINIT,
      SEL => addr2ext_10_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_10
    );
  tx_output_addr_Madd_n0000_inst_sum_10 : X_XOR2
    port map (
      I0 => addr2ext_10_CYINIT,
      I1 => addr2ext_10_FROM,
      O => tx_output_addr_n0000(10)
    );
  addr2ext_10_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr2ext_10_FROM
    );
  addr2ext_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(11),
      O => addr2ext_10_GROM
    );
  addr2ext_10_COUTUSED : X_BUF
    port map (
      I => addr2ext_10_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_11
    );
  tx_output_addr_Madd_n0000_inst_cy_11_317 : X_MUX2
    port map (
      IA => addr2ext_10_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_10,
      SEL => addr2ext_10_GROM,
      O => addr2ext_10_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_11 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_10,
      I1 => addr2ext_10_GROM,
      O => tx_output_addr_n0000(11)
    );
  addr2ext_10_CYINIT_318 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_9,
      O => addr2ext_10_CYINIT
    );
  addr2ext_12_LOGIC_ZERO_319 : X_ZERO
    port map (
      O => addr2ext_12_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_12_320 : X_MUX2
    port map (
      IA => addr2ext_12_LOGIC_ZERO,
      IB => addr2ext_12_CYINIT,
      SEL => addr2ext_12_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_12
    );
  tx_output_addr_Madd_n0000_inst_sum_12 : X_XOR2
    port map (
      I0 => addr2ext_12_CYINIT,
      I1 => addr2ext_12_FROM,
      O => tx_output_addr_n0000(12)
    );
  addr2ext_12_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr2ext(12),
      ADR3 => VCC,
      O => addr2ext_12_FROM
    );
  addr2ext_12_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr2ext_12_GROM
    );
  addr2ext_12_COUTUSED : X_BUF
    port map (
      I => addr2ext_12_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_13
    );
  tx_output_addr_Madd_n0000_inst_cy_13_321 : X_MUX2
    port map (
      IA => addr2ext_12_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_12,
      SEL => addr2ext_12_GROM,
      O => addr2ext_12_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_13 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_12,
      I1 => addr2ext_12_GROM,
      O => tx_output_addr_n0000(13)
    );
  addr2ext_12_CYINIT_322 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_11,
      O => addr2ext_12_CYINIT
    );
  addr2ext_14_LOGIC_ZERO_323 : X_ZERO
    port map (
      O => addr2ext_14_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_14_324 : X_MUX2
    port map (
      IA => addr2ext_14_LOGIC_ZERO,
      IB => addr2ext_14_CYINIT,
      SEL => addr2ext_14_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_14
    );
  tx_output_addr_Madd_n0000_inst_sum_14 : X_XOR2
    port map (
      I0 => addr2ext_14_CYINIT,
      I1 => addr2ext_14_FROM,
      O => tx_output_addr_n0000(14)
    );
  addr2ext_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr2ext_14_FROM
    );
  addr2ext_15_rt_325 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(15),
      O => addr2ext_15_rt
    );
  tx_output_addr_Madd_n0000_inst_sum_15 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_14,
      I1 => addr2ext_15_rt,
      O => tx_output_addr_n0000(15)
    );
  addr2ext_14_CYINIT_326 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_13,
      O => addr2ext_14_CYINIT
    );
  rx_input_memio_bcnt_86_LOGIC_ZERO_327 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_86_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_270_328 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1,
      IB => rx_input_memio_bcnt_86_LOGIC_ZERO,
      SEL => rx_input_memio_cs_FFd16_rt,
      O => rx_input_memio_bcnt_inst_cy_270
    );
  rx_input_memio_cs_FFd16_rt_329 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_cs_FFd16_rt
    );
  rx_input_memio_bcnt_inst_lut3_721 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_0,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcnt_86,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_72
    );
  rx_input_memio_bcnt_86_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_86_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_271
    );
  rx_input_memio_bcnt_inst_cy_271_330 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_0,
      IB => rx_input_memio_bcnt_inst_cy_270,
      SEL => rx_input_memio_bcnt_inst_lut3_72,
      O => rx_input_memio_bcnt_86_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_235_331 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_270,
      I1 => rx_input_memio_bcnt_inst_lut3_72,
      O => rx_input_memio_bcnt_inst_sum_235
    );
  rx_input_memio_bcnt_87_LOGIC_ZERO_332 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_87_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_272_333 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_87_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_87_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_73,
      O => rx_input_memio_bcnt_inst_cy_272
    );
  rx_input_memio_bcnt_inst_sum_236_334 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_87_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_73,
      O => rx_input_memio_bcnt_inst_sum_236
    );
  rx_input_memio_bcnt_inst_lut3_731 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcnt_87,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_73
    );
  rx_input_memio_bcnt_inst_lut3_741 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_88,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_74
    );
  rx_input_memio_bcnt_87_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_87_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_273
    );
  rx_input_memio_bcnt_inst_cy_273_335 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_87_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_272,
      SEL => rx_input_memio_bcnt_inst_lut3_74,
      O => rx_input_memio_bcnt_87_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_237_336 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_272,
      I1 => rx_input_memio_bcnt_inst_lut3_74,
      O => rx_input_memio_bcnt_inst_sum_237
    );
  rx_input_memio_bcnt_87_CYINIT_337 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_271,
      O => rx_input_memio_bcnt_87_CYINIT
    );
  rx_input_memio_bcnt_89_LOGIC_ZERO_338 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_89_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_274_339 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_89_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_89_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_75,
      O => rx_input_memio_bcnt_inst_cy_274
    );
  rx_input_memio_bcnt_inst_sum_238_340 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_89_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_75,
      O => rx_input_memio_bcnt_inst_sum_238
    );
  rx_input_memio_bcnt_inst_lut3_751 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => rx_input_memio_bcnt_89,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_75
    );
  rx_input_memio_bcnt_inst_lut3_761 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => rx_input_memio_bcnt_90,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_76
    );
  rx_input_memio_bcnt_89_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_89_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_275
    );
  rx_input_memio_bcnt_inst_cy_275_341 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_89_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_274,
      SEL => rx_input_memio_bcnt_inst_lut3_76,
      O => rx_input_memio_bcnt_89_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_239_342 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_274,
      I1 => rx_input_memio_bcnt_inst_lut3_76,
      O => rx_input_memio_bcnt_inst_sum_239
    );
  rx_input_memio_bcnt_89_CYINIT_343 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_273,
      O => rx_input_memio_bcnt_89_CYINIT
    );
  rx_input_memio_bcnt_91_LOGIC_ZERO_344 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_91_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_276_345 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_91_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_91_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_77,
      O => rx_input_memio_bcnt_inst_cy_276
    );
  rx_input_memio_bcnt_inst_sum_240_346 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_91_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_77,
      O => rx_input_memio_bcnt_inst_sum_240
    );
  rx_input_memio_bcnt_inst_lut3_771 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcnt_91,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_77
    );
  rx_input_memio_bcnt_inst_lut3_781 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_92,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_78
    );
  rx_input_memio_bcnt_91_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_91_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_277
    );
  rx_input_memio_bcnt_inst_cy_277_347 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_91_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_276,
      SEL => rx_input_memio_bcnt_inst_lut3_78,
      O => rx_input_memio_bcnt_91_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_241_348 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_276,
      I1 => rx_input_memio_bcnt_inst_lut3_78,
      O => rx_input_memio_bcnt_inst_sum_241
    );
  rx_input_memio_bcnt_91_CYINIT_349 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_275,
      O => rx_input_memio_bcnt_91_CYINIT
    );
  rx_input_memio_bcnt_93_LOGIC_ZERO_350 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_93_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_278_351 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_93_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_93_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_79,
      O => rx_input_memio_bcnt_inst_cy_278
    );
  rx_input_memio_bcnt_inst_sum_242_352 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_93_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_79,
      O => rx_input_memio_bcnt_inst_sum_242
    );
  rx_input_memio_bcnt_inst_lut3_791 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcnt_93,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_79
    );
  rx_input_memio_bcnt_inst_lut3_801 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcnt_94,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_80
    );
  rx_input_memio_bcnt_93_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_93_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_279
    );
  rx_input_memio_bcnt_inst_cy_279_353 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_93_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_278,
      SEL => rx_input_memio_bcnt_inst_lut3_80,
      O => rx_input_memio_bcnt_93_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_243_354 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_278,
      I1 => rx_input_memio_bcnt_inst_lut3_80,
      O => rx_input_memio_bcnt_inst_sum_243
    );
  rx_input_memio_bcnt_93_CYINIT_355 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_277,
      O => rx_input_memio_bcnt_93_CYINIT
    );
  rx_input_memio_bcnt_95_LOGIC_ZERO_356 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_95_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_280_357 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_95_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_95_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_81,
      O => rx_input_memio_bcnt_inst_cy_280
    );
  rx_input_memio_bcnt_inst_sum_244_358 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_95_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_81,
      O => rx_input_memio_bcnt_inst_sum_244
    );
  rx_input_memio_bcnt_inst_lut3_811 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => rx_input_memio_bcnt_95,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_81
    );
  rx_input_memio_bcnt_inst_lut3_821 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => rx_input_memio_bcnt_96,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_82
    );
  rx_input_memio_bcnt_95_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_95_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_281
    );
  rx_input_memio_bcnt_inst_cy_281_359 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_95_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_280,
      SEL => rx_input_memio_bcnt_inst_lut3_82,
      O => rx_input_memio_bcnt_95_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_245_360 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_280,
      I1 => rx_input_memio_bcnt_inst_lut3_82,
      O => rx_input_memio_bcnt_inst_sum_245
    );
  rx_input_memio_bcnt_95_CYINIT_361 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_279,
      O => rx_input_memio_bcnt_95_CYINIT
    );
  rx_input_memio_bcnt_97_LOGIC_ZERO_362 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_97_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_282_363 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_97_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_97_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_83,
      O => rx_input_memio_bcnt_inst_cy_282
    );
  rx_input_memio_bcnt_inst_sum_246_364 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_97_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_83,
      O => rx_input_memio_bcnt_inst_sum_246
    );
  rx_input_memio_bcnt_inst_lut3_831 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcnt_97,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_83
    );
  rx_input_memio_bcnt_inst_lut3_841 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcnt_98,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_84
    );
  rx_input_memio_bcnt_97_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_97_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_283
    );
  rx_input_memio_bcnt_inst_cy_283_365 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_97_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_282,
      SEL => rx_input_memio_bcnt_inst_lut3_84,
      O => rx_input_memio_bcnt_97_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_247_366 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_282,
      I1 => rx_input_memio_bcnt_inst_lut3_84,
      O => rx_input_memio_bcnt_inst_sum_247
    );
  rx_input_memio_bcnt_97_CYINIT_367 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_281,
      O => rx_input_memio_bcnt_97_CYINIT
    );
  rx_input_memio_bcnt_99_LOGIC_ZERO_368 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_99_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_284_369 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_99_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_99_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_85,
      O => rx_input_memio_bcnt_inst_cy_284
    );
  rx_input_memio_bcnt_inst_sum_248_370 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_99_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_85,
      O => rx_input_memio_bcnt_inst_sum_248
    );
  rx_input_memio_bcnt_inst_lut3_851 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcnt_99,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_85
    );
  rx_input_memio_bcnt_inst_lut3_861 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_100,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_86
    );
  rx_input_memio_bcnt_99_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_99_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_285
    );
  rx_input_memio_bcnt_inst_cy_285_371 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_99_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_284,
      SEL => rx_input_memio_bcnt_inst_lut3_86,
      O => rx_input_memio_bcnt_99_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_249_372 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_284,
      I1 => rx_input_memio_bcnt_inst_lut3_86,
      O => rx_input_memio_bcnt_inst_sum_249
    );
  rx_input_memio_bcnt_99_CYINIT_373 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_283,
      O => rx_input_memio_bcnt_99_CYINIT
    );
  rx_input_memio_bcnt_inst_sum_250_374 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_101_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_87,
      O => rx_input_memio_bcnt_inst_sum_250
    );
  rx_input_memio_bcnt_inst_lut3_871 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_101,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_87
    );
  rx_input_memio_cs_Out916_SW0_2_375 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd1,
      ADR2 => rx_input_memio_cs_FFd15,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_101_GROM
    );
  rx_input_memio_bcnt_101_YUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_101_GROM,
      O => rx_input_memio_cs_Out916_SW0_2
    );
  rx_input_memio_bcnt_101_CYINIT_376 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_285,
      O => rx_input_memio_bcnt_101_CYINIT
    );
  rx_output_Madd_n0060_inst_cy_49_LOGIC_ZERO_377 : X_ZERO
    port map (
      O => rx_output_Madd_n0060_inst_cy_49_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_48_378 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_19,
      IB => rx_output_Madd_n0060_inst_cy_49_LOGIC_ZERO,
      SEL => rx_output_Madd_n0060_inst_lut2_48,
      O => rx_output_Madd_n0060_inst_cy_48
    );
  rx_output_Madd_n0060_inst_lut2_4811 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_19,
      ADR1 => rx_output_len(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_Madd_n0060_inst_lut2_48
    );
  rx_output_Madd_n0060_inst_lut2_491 : X_LUT4
    generic map(
      INIT => X"EEEE"
    )
    port map (
      ADR0 => rx_output_len(1),
      ADR1 => rx_output_len(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_Madd_n0060_inst_lut2_49
    );
  rx_output_Madd_n0060_inst_cy_49_COUTUSED : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_49_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_49
    );
  rx_output_Madd_n0060_inst_cy_49_379 : X_MUX2
    port map (
      IA => rx_output_len(1),
      IB => rx_output_Madd_n0060_inst_cy_48,
      SEL => rx_output_Madd_n0060_inst_lut2_49,
      O => rx_output_Madd_n0060_inst_cy_49_CYMUXG
    );
  rx_output_n0060_2_LOGIC_ZERO_380 : X_ZERO
    port map (
      O => rx_output_n0060_2_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_50_381 : X_MUX2
    port map (
      IA => rx_output_n0060_2_LOGIC_ZERO,
      IB => rx_output_n0060_2_CYINIT,
      SEL => rx_output_n0060_2_FROM,
      O => rx_output_Madd_n0060_inst_cy_50
    );
  rx_output_Madd_n0060_inst_sum_50 : X_XOR2
    port map (
      I0 => rx_output_n0060_2_CYINIT,
      I1 => rx_output_n0060_2_FROM,
      O => rx_output_n0060_2_XORF
    );
  rx_output_n0060_2_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_2_FROM
    );
  rx_output_n0060_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(3),
      ADR3 => VCC,
      O => rx_output_n0060_2_GROM
    );
  rx_output_n0060_2_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_2_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_51
    );
  rx_output_n0060_2_XUSED : X_BUF
    port map (
      I => rx_output_n0060_2_XORF,
      O => rx_output_n0060(2)
    );
  rx_output_n0060_2_YUSED : X_BUF
    port map (
      I => rx_output_n0060_2_XORG,
      O => rx_output_n0060(3)
    );
  rx_output_Madd_n0060_inst_cy_51_382 : X_MUX2
    port map (
      IA => rx_output_n0060_2_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_50,
      SEL => rx_output_n0060_2_GROM,
      O => rx_output_n0060_2_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_51 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_50,
      I1 => rx_output_n0060_2_GROM,
      O => rx_output_n0060_2_XORG
    );
  rx_output_n0060_2_CYINIT_383 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_49,
      O => rx_output_n0060_2_CYINIT
    );
  rx_output_n0060_4_LOGIC_ZERO_384 : X_ZERO
    port map (
      O => rx_output_n0060_4_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_52_385 : X_MUX2
    port map (
      IA => rx_output_n0060_4_LOGIC_ZERO,
      IB => rx_output_n0060_4_CYINIT,
      SEL => rx_output_n0060_4_FROM,
      O => rx_output_Madd_n0060_inst_cy_52
    );
  rx_output_Madd_n0060_inst_sum_52 : X_XOR2
    port map (
      I0 => rx_output_n0060_4_CYINIT,
      I1 => rx_output_n0060_4_FROM,
      O => rx_output_n0060_4_XORF
    );
  rx_output_n0060_4_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(4),
      O => rx_output_n0060_4_FROM
    );
  rx_output_n0060_4_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_4_GROM
    );
  rx_output_n0060_4_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_4_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_53
    );
  rx_output_n0060_4_XUSED : X_BUF
    port map (
      I => rx_output_n0060_4_XORF,
      O => rx_output_n0060(4)
    );
  rx_output_n0060_4_YUSED : X_BUF
    port map (
      I => rx_output_n0060_4_XORG,
      O => rx_output_n0060(5)
    );
  rx_output_Madd_n0060_inst_cy_53_386 : X_MUX2
    port map (
      IA => rx_output_n0060_4_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_52,
      SEL => rx_output_n0060_4_GROM,
      O => rx_output_n0060_4_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_53 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_52,
      I1 => rx_output_n0060_4_GROM,
      O => rx_output_n0060_4_XORG
    );
  rx_output_n0060_4_CYINIT_387 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_51,
      O => rx_output_n0060_4_CYINIT
    );
  rx_output_n0060_6_LOGIC_ZERO_388 : X_ZERO
    port map (
      O => rx_output_n0060_6_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_54_389 : X_MUX2
    port map (
      IA => rx_output_n0060_6_LOGIC_ZERO,
      IB => rx_output_n0060_6_CYINIT,
      SEL => rx_output_n0060_6_FROM,
      O => rx_output_Madd_n0060_inst_cy_54
    );
  rx_output_Madd_n0060_inst_sum_54 : X_XOR2
    port map (
      I0 => rx_output_n0060_6_CYINIT,
      I1 => rx_output_n0060_6_FROM,
      O => rx_output_n0060_6_XORF
    );
  rx_output_n0060_6_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(6),
      O => rx_output_n0060_6_FROM
    );
  rx_output_n0060_6_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_6_GROM
    );
  rx_output_n0060_6_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_6_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_55
    );
  rx_output_n0060_6_XUSED : X_BUF
    port map (
      I => rx_output_n0060_6_XORF,
      O => rx_output_n0060(6)
    );
  rx_output_n0060_6_YUSED : X_BUF
    port map (
      I => rx_output_n0060_6_XORG,
      O => rx_output_n0060(7)
    );
  rx_output_Madd_n0060_inst_cy_55_390 : X_MUX2
    port map (
      IA => rx_output_n0060_6_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_54,
      SEL => rx_output_n0060_6_GROM,
      O => rx_output_n0060_6_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_55 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_54,
      I1 => rx_output_n0060_6_GROM,
      O => rx_output_n0060_6_XORG
    );
  rx_output_n0060_6_CYINIT_391 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_53,
      O => rx_output_n0060_6_CYINIT
    );
  rx_output_n0060_8_LOGIC_ZERO_392 : X_ZERO
    port map (
      O => rx_output_n0060_8_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_56_393 : X_MUX2
    port map (
      IA => rx_output_n0060_8_LOGIC_ZERO,
      IB => rx_output_n0060_8_CYINIT,
      SEL => rx_output_n0060_8_FROM,
      O => rx_output_Madd_n0060_inst_cy_56
    );
  rx_output_Madd_n0060_inst_sum_56 : X_XOR2
    port map (
      I0 => rx_output_n0060_8_CYINIT,
      I1 => rx_output_n0060_8_FROM,
      O => rx_output_n0060_8_XORF
    );
  rx_output_n0060_8_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_8_FROM
    );
  rx_output_n0060_8_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_8_GROM
    );
  rx_output_n0060_8_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_8_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_57
    );
  rx_output_n0060_8_XUSED : X_BUF
    port map (
      I => rx_output_n0060_8_XORF,
      O => rx_output_n0060(8)
    );
  rx_output_n0060_8_YUSED : X_BUF
    port map (
      I => rx_output_n0060_8_XORG,
      O => rx_output_n0060(9)
    );
  rx_output_Madd_n0060_inst_cy_57_394 : X_MUX2
    port map (
      IA => rx_output_n0060_8_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_56,
      SEL => rx_output_n0060_8_GROM,
      O => rx_output_n0060_8_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_57 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_56,
      I1 => rx_output_n0060_8_GROM,
      O => rx_output_n0060_8_XORG
    );
  rx_output_n0060_8_CYINIT_395 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_55,
      O => rx_output_n0060_8_CYINIT
    );
  rx_output_n0060_10_LOGIC_ZERO_396 : X_ZERO
    port map (
      O => rx_output_n0060_10_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_58_397 : X_MUX2
    port map (
      IA => rx_output_n0060_10_LOGIC_ZERO,
      IB => rx_output_n0060_10_CYINIT,
      SEL => rx_output_n0060_10_FROM,
      O => rx_output_Madd_n0060_inst_cy_58
    );
  rx_output_Madd_n0060_inst_sum_58 : X_XOR2
    port map (
      I0 => rx_output_n0060_10_CYINIT,
      I1 => rx_output_n0060_10_FROM,
      O => rx_output_n0060_10_XORF
    );
  rx_output_n0060_10_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(10),
      O => rx_output_n0060_10_FROM
    );
  rx_output_n0060_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(11),
      O => rx_output_n0060_10_GROM
    );
  rx_output_n0060_10_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_10_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_59
    );
  rx_output_n0060_10_XUSED : X_BUF
    port map (
      I => rx_output_n0060_10_XORF,
      O => rx_output_n0060(10)
    );
  rx_output_n0060_10_YUSED : X_BUF
    port map (
      I => rx_output_n0060_10_XORG,
      O => rx_output_n0060(11)
    );
  rx_output_Madd_n0060_inst_cy_59_398 : X_MUX2
    port map (
      IA => rx_output_n0060_10_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_58,
      SEL => rx_output_n0060_10_GROM,
      O => rx_output_n0060_10_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_59 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_58,
      I1 => rx_output_n0060_10_GROM,
      O => rx_output_n0060_10_XORG
    );
  rx_output_n0060_10_CYINIT_399 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_57,
      O => rx_output_n0060_10_CYINIT
    );
  rx_output_n0060_12_LOGIC_ZERO_400 : X_ZERO
    port map (
      O => rx_output_n0060_12_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_60_401 : X_MUX2
    port map (
      IA => rx_output_n0060_12_LOGIC_ZERO,
      IB => rx_output_n0060_12_CYINIT,
      SEL => rx_output_n0060_12_FROM,
      O => rx_output_Madd_n0060_inst_cy_60
    );
  rx_output_Madd_n0060_inst_sum_60 : X_XOR2
    port map (
      I0 => rx_output_n0060_12_CYINIT,
      I1 => rx_output_n0060_12_FROM,
      O => rx_output_n0060_12_XORF
    );
  rx_output_n0060_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_12_FROM
    );
  rx_output_n0060_12_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_12_GROM
    );
  rx_output_n0060_12_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_12_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_61
    );
  rx_output_n0060_12_XUSED : X_BUF
    port map (
      I => rx_output_n0060_12_XORF,
      O => rx_output_n0060(12)
    );
  rx_output_n0060_12_YUSED : X_BUF
    port map (
      I => rx_output_n0060_12_XORG,
      O => rx_output_n0060(13)
    );
  rx_output_Madd_n0060_inst_cy_61_402 : X_MUX2
    port map (
      IA => rx_output_n0060_12_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_60,
      SEL => rx_output_n0060_12_GROM,
      O => rx_output_n0060_12_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_61 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_60,
      I1 => rx_output_n0060_12_GROM,
      O => rx_output_n0060_12_XORG
    );
  rx_output_n0060_12_CYINIT_403 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_59,
      O => rx_output_n0060_12_CYINIT
    );
  rx_output_n0060_14_LOGIC_ZERO_404 : X_ZERO
    port map (
      O => rx_output_n0060_14_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_62_405 : X_MUX2
    port map (
      IA => rx_output_n0060_14_LOGIC_ZERO,
      IB => rx_output_n0060_14_CYINIT,
      SEL => rx_output_n0060_14_FROM,
      O => rx_output_Madd_n0060_inst_cy_62
    );
  rx_output_Madd_n0060_inst_sum_62 : X_XOR2
    port map (
      I0 => rx_output_n0060_14_CYINIT,
      I1 => rx_output_n0060_14_FROM,
      O => rx_output_n0060_14_XORF
    );
  rx_output_n0060_14_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(14),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_14_FROM
    );
  rx_output_len_15_rt_406 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(15),
      ADR3 => VCC,
      O => rx_output_len_15_rt
    );
  rx_output_n0060_14_XUSED : X_BUF
    port map (
      I => rx_output_n0060_14_XORF,
      O => rx_output_n0060(14)
    );
  rx_output_n0060_14_YUSED : X_BUF
    port map (
      I => rx_output_n0060_14_XORG,
      O => rx_output_n0060(15)
    );
  rx_output_Madd_n0060_inst_sum_63 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_62,
      I1 => rx_output_len_15_rt,
      O => rx_output_n0060_14_XORG
    );
  rx_output_n0060_14_CYINIT_407 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_61,
      O => rx_output_n0060_14_CYINIT
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ONE_408 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ZERO_409 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_177_410 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(8),
      ADR1 => rx_input_memio_addrchk_datal(9),
      ADR2 => rx_input_memio_addrchk_macaddrl(9),
      ADR3 => rx_input_memio_addrchk_macaddrl(8),
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(10),
      ADR1 => rx_input_memio_addrchk_datal(11),
      ADR2 => rx_input_memio_addrchk_macaddrl(11),
      ADR3 => rx_input_memio_addrchk_macaddrl(10),
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_411 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_4_LOGIC_ZERO_412 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_4_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_179_413 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_4_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_4_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(13),
      ADR1 => rx_input_memio_addrchk_datal(12),
      ADR2 => rx_input_memio_addrchk_macaddrl(12),
      ADR3 => rx_input_memio_addrchk_macaddrl(13),
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(15),
      ADR1 => rx_input_memio_addrchk_datal(14),
      ADR2 => rx_input_memio_addrchk_macaddrl(14),
      ADR3 => rx_input_memio_addrchk_macaddrl(15),
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_4_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_4_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(4)
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_4_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_4_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_4_CYINIT_414 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_4_CYINIT
    );
  mac_control_rxcrcerr_cnt_0_LOGIC_ZERO_415 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_0_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_16_416 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_31,
      IB => mac_control_rxcrcerr_cnt_0_LOGIC_ZERO,
      SEL => mac_control_rxcrcerr_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_31,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(0),
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_rxcrcerr_cnt_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_57,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(1),
      O => mac_control_rxcrcerr_cnt_0_GROM
    );
  mac_control_rxcrcerr_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_0_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_17_417 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_57,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_rxcrcerr_cnt_0_GROM,
      O => mac_control_rxcrcerr_cnt_0_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_rxcrcerr_cnt_0_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(1)
    );
  mac_control_rxcrcerr_cnt_2_LOGIC_ZERO_418 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_2_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_18_419 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_2_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_2_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_2_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_2_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(2)
    );
  mac_control_rxcrcerr_cnt_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(2),
      O => mac_control_rxcrcerr_cnt_2_FROM
    );
  mac_control_rxcrcerr_cnt_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(3),
      O => mac_control_rxcrcerr_cnt_2_GROM
    );
  mac_control_rxcrcerr_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_2_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_19_420 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_rxcrcerr_cnt_2_GROM,
      O => mac_control_rxcrcerr_cnt_2_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_rxcrcerr_cnt_2_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(3)
    );
  mac_control_rxcrcerr_cnt_2_CYINIT_421 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_rxcrcerr_cnt_2_CYINIT
    );
  mac_control_rxcrcerr_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(5),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(5)
    );
  mac_control_rxcrcerr_cnt_4_LOGIC_ZERO_422 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_4_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_20_423 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_4_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_4_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_4_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_4_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(4)
    );
  mac_control_rxcrcerr_cnt_4_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(4),
      O => mac_control_rxcrcerr_cnt_4_FROM
    );
  mac_control_rxcrcerr_cnt_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(5),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_4_GROM
    );
  mac_control_rxcrcerr_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_4_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_21_424 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_rxcrcerr_cnt_4_GROM,
      O => mac_control_rxcrcerr_cnt_4_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_rxcrcerr_cnt_4_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(5)
    );
  mac_control_rxcrcerr_cnt_4_CYINIT_425 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_rxcrcerr_cnt_4_CYINIT
    );
  mac_control_rxcrcerr_cnt_6_LOGIC_ZERO_426 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_6_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_22_427 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_6_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_6_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_6_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_6_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(6)
    );
  mac_control_rxcrcerr_cnt_6_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxcrcerr_cnt(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_6_FROM
    );
  mac_control_rxcrcerr_cnt_6_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(7),
      O => mac_control_rxcrcerr_cnt_6_GROM
    );
  mac_control_rxcrcerr_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_6_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_23_428 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_rxcrcerr_cnt_6_GROM,
      O => mac_control_rxcrcerr_cnt_6_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_rxcrcerr_cnt_6_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(7)
    );
  mac_control_rxcrcerr_cnt_6_CYINIT_429 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_rxcrcerr_cnt_6_CYINIT
    );
  mac_control_rxcrcerr_cnt_8_LOGIC_ZERO_430 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_8_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_24_431 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_8_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_8_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_8_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_8_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(8)
    );
  mac_control_rxcrcerr_cnt_8_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(8),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_8_FROM
    );
  mac_control_rxcrcerr_cnt_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(9),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_8_GROM
    );
  mac_control_rxcrcerr_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_8_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_25_432 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_rxcrcerr_cnt_8_GROM,
      O => mac_control_rxcrcerr_cnt_8_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_rxcrcerr_cnt_8_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(9)
    );
  mac_control_rxcrcerr_cnt_8_CYINIT_433 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_rxcrcerr_cnt_8_CYINIT
    );
  mac_control_rxcrcerr_cnt_10_LOGIC_ZERO_434 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_10_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_26_435 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_10_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_10_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_10_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_10_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(10)
    );
  mac_control_rxcrcerr_cnt_10_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxcrcerr_cnt(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_10_FROM
    );
  mac_control_rxcrcerr_cnt_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(11),
      O => mac_control_rxcrcerr_cnt_10_GROM
    );
  mac_control_rxcrcerr_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_10_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_27_436 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_rxcrcerr_cnt_10_GROM,
      O => mac_control_rxcrcerr_cnt_10_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_rxcrcerr_cnt_10_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(11)
    );
  mac_control_rxcrcerr_cnt_10_CYINIT_437 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_rxcrcerr_cnt_10_CYINIT
    );
  rx_input_fifo_fifo_BU77 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2809,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N17_FFX_RST,
      O => rx_input_fifo_fifo_N17
    );
  rx_input_fifo_fifo_N17_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N17_FFX_RST
    );
  mac_control_rxcrcerr_cnt_12_LOGIC_ZERO_438 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_12_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_28_439 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_12_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_12_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_12_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_12_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(12)
    );
  mac_control_rxcrcerr_cnt_12_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(12),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_12_FROM
    );
  mac_control_rxcrcerr_cnt_12_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(13),
      O => mac_control_rxcrcerr_cnt_12_GROM
    );
  mac_control_rxcrcerr_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_12_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_29_440 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_rxcrcerr_cnt_12_GROM,
      O => mac_control_rxcrcerr_cnt_12_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_rxcrcerr_cnt_12_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(13)
    );
  mac_control_rxcrcerr_cnt_12_CYINIT_441 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_rxcrcerr_cnt_12_CYINIT
    );
  mac_control_rxcrcerr_cnt_14_LOGIC_ZERO_442 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_14_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_30_443 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_14_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_14_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_14_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_14_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(14)
    );
  mac_control_rxcrcerr_cnt_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxcrcerr_cnt(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_14_FROM
    );
  mac_control_rxcrcerr_cnt_14_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(15),
      O => mac_control_rxcrcerr_cnt_14_GROM
    );
  mac_control_rxcrcerr_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_14_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_31_444 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_rxcrcerr_cnt_14_GROM,
      O => mac_control_rxcrcerr_cnt_14_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_rxcrcerr_cnt_14_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(15)
    );
  mac_control_rxcrcerr_cnt_14_CYINIT_445 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_rxcrcerr_cnt_14_CYINIT
    );
  mac_control_rxcrcerr_cnt_16_LOGIC_ZERO_446 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_16_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_32_447 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_16_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_16_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_16_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_16_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(16)
    );
  mac_control_rxcrcerr_cnt_16_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(16),
      O => mac_control_rxcrcerr_cnt_16_FROM
    );
  mac_control_rxcrcerr_cnt_16_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(17),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_16_GROM
    );
  mac_control_rxcrcerr_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_16_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_33_448 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_rxcrcerr_cnt_16_GROM,
      O => mac_control_rxcrcerr_cnt_16_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_rxcrcerr_cnt_16_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(17)
    );
  mac_control_rxcrcerr_cnt_16_CYINIT_449 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_rxcrcerr_cnt_16_CYINIT
    );
  mac_control_rxcrcerr_cnt_18_LOGIC_ZERO_450 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_18_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_34_451 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_18_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_18_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_18_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_18_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(18)
    );
  mac_control_rxcrcerr_cnt_18_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxcrcerr_cnt(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_18_FROM
    );
  mac_control_rxcrcerr_cnt_18_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(19),
      O => mac_control_rxcrcerr_cnt_18_GROM
    );
  mac_control_rxcrcerr_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_18_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_35_452 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_rxcrcerr_cnt_18_GROM,
      O => mac_control_rxcrcerr_cnt_18_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_rxcrcerr_cnt_18_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(19)
    );
  mac_control_rxcrcerr_cnt_18_CYINIT_453 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_rxcrcerr_cnt_18_CYINIT
    );
  mac_control_rxcrcerr_cnt_20_LOGIC_ZERO_454 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_20_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_36_455 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_20_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_20_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_20_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_20_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(20)
    );
  mac_control_rxcrcerr_cnt_20_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(20),
      O => mac_control_rxcrcerr_cnt_20_FROM
    );
  mac_control_rxcrcerr_cnt_20_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxcrcerr_cnt(21),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_20_GROM
    );
  mac_control_rxcrcerr_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_20_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_37_456 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_rxcrcerr_cnt_20_GROM,
      O => mac_control_rxcrcerr_cnt_20_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_rxcrcerr_cnt_20_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(21)
    );
  mac_control_rxcrcerr_cnt_20_CYINIT_457 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_rxcrcerr_cnt_20_CYINIT
    );
  mac_control_rxcrcerr_cnt_22_LOGIC_ZERO_458 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_22_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_38_459 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_22_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_22_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_22_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_22_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(22)
    );
  mac_control_rxcrcerr_cnt_22_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxcrcerr_cnt(22),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_22_FROM
    );
  mac_control_rxcrcerr_cnt_22_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(23),
      O => mac_control_rxcrcerr_cnt_22_GROM
    );
  mac_control_rxcrcerr_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_22_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_39_460 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_rxcrcerr_cnt_22_GROM,
      O => mac_control_rxcrcerr_cnt_22_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_rxcrcerr_cnt_22_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(23)
    );
  mac_control_rxcrcerr_cnt_22_CYINIT_461 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_rxcrcerr_cnt_22_CYINIT
    );
  mac_control_rxcrcerr_cnt_24_LOGIC_ZERO_462 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_24_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_40_463 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_24_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_24_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_24_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_24_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(24)
    );
  mac_control_rxcrcerr_cnt_24_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(24),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_24_FROM
    );
  mac_control_rxcrcerr_cnt_24_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(25),
      O => mac_control_rxcrcerr_cnt_24_GROM
    );
  mac_control_rxcrcerr_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_24_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_41_464 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_rxcrcerr_cnt_24_GROM,
      O => mac_control_rxcrcerr_cnt_24_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_rxcrcerr_cnt_24_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(25)
    );
  mac_control_rxcrcerr_cnt_24_CYINIT_465 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_rxcrcerr_cnt_24_CYINIT
    );
  mac_control_rxcrcerr_cnt_26_LOGIC_ZERO_466 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_26_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_42_467 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_26_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_26_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_26_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_26_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(26)
    );
  mac_control_rxcrcerr_cnt_26_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(26),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_26_FROM
    );
  mac_control_rxcrcerr_cnt_26_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(27),
      O => mac_control_rxcrcerr_cnt_26_GROM
    );
  mac_control_rxcrcerr_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_26_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_43_468 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_rxcrcerr_cnt_26_GROM,
      O => mac_control_rxcrcerr_cnt_26_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_rxcrcerr_cnt_26_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(27)
    );
  mac_control_rxcrcerr_cnt_26_CYINIT_469 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_rxcrcerr_cnt_26_CYINIT
    );
  mac_control_rxcrcerr_cnt_28_LOGIC_ZERO_470 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_28_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_44_471 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_28_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_28_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_28_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_28_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(28)
    );
  mac_control_rxcrcerr_cnt_28_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(28),
      O => mac_control_rxcrcerr_cnt_28_FROM
    );
  mac_control_rxcrcerr_cnt_28_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(29),
      O => mac_control_rxcrcerr_cnt_28_GROM
    );
  mac_control_rxcrcerr_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_28_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_45_472 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_rxcrcerr_cnt_28_GROM,
      O => mac_control_rxcrcerr_cnt_28_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_rxcrcerr_cnt_28_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(29)
    );
  mac_control_rxcrcerr_cnt_28_CYINIT_473 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_rxcrcerr_cnt_28_CYINIT
    );
  mac_control_rxcrcerr_cnt_30_LOGIC_ZERO_474 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_30_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_46_475 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_30_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_30_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_30_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_30_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_30_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(30)
    );
  mac_control_rxcrcerr_cnt_30_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(30),
      O => mac_control_rxcrcerr_cnt_30_FROM
    );
  mac_control_rxcrcerr_cnt_31_rt_476 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(31),
      O => mac_control_rxcrcerr_cnt_31_rt
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_rxcrcerr_cnt_31_rt,
      O => mac_control_rxcrcerr_cnt_n0000(31)
    );
  mac_control_rxcrcerr_cnt_30_CYINIT_477 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_rxcrcerr_cnt_30_CYINIT
    );
  rx_input_memio_bp_0_LOGIC_ONE_478 : X_ONE
    port map (
      O => rx_input_memio_bp_0_LOGIC_ONE
    );
  rx_input_memio_Msub_n0043_inst_cy_221_479 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_42,
      IB => rx_input_memio_bp_0_CYINIT,
      SEL => rx_input_memio_bp_0_FROM,
      O => rx_input_memio_Msub_n0043_inst_cy_221
    );
  rx_input_memio_Msub_n0043_inst_sum_187 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_0_CYINIT,
      I1 => rx_input_memio_bp_0_FROM,
      O => rx_input_memio_n0043(0)
    );
  rx_input_memio_bp_0_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_42,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_macnt_70,
      O => rx_input_memio_bp_0_FROM
    );
  rx_input_memio_Msub_n0043_inst_lut2_1341 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_71,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_134
    );
  rx_input_memio_bp_0_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_0_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_222
    );
  rx_input_memio_Msub_n0043_inst_cy_222_480 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_71,
      IB => rx_input_memio_Msub_n0043_inst_cy_221,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_134,
      O => rx_input_memio_bp_0_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_188 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_221,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_134,
      O => rx_input_memio_n0043(1)
    );
  rx_input_memio_bp_0_CYINIT_481 : X_BUF
    port map (
      I => rx_input_memio_bp_0_LOGIC_ONE,
      O => rx_input_memio_bp_0_CYINIT
    );
  rx_input_memio_bp_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_2_FFY_RST
    );
  rx_input_memio_bp_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(3),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_2_FFY_RST,
      O => rx_input_memio_bp(3)
    );
  rx_input_memio_Msub_n0043_inst_cy_223_482 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_72,
      IB => rx_input_memio_bp_2_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_135,
      O => rx_input_memio_Msub_n0043_inst_cy_223
    );
  rx_input_memio_Msub_n0043_inst_sum_189 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_2_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_135,
      O => rx_input_memio_n0043(2)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1351 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_72,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_135
    );
  rx_input_memio_Msub_n0043_inst_lut2_1361 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_73,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_136
    );
  rx_input_memio_bp_2_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_2_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_224
    );
  rx_input_memio_Msub_n0043_inst_cy_224_483 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_73,
      IB => rx_input_memio_Msub_n0043_inst_cy_223,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_136,
      O => rx_input_memio_bp_2_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_190 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_223,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_136,
      O => rx_input_memio_n0043(3)
    );
  rx_input_memio_bp_2_CYINIT_484 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_222,
      O => rx_input_memio_bp_2_CYINIT
    );
  rx_input_fifo_fifo_BU136 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3360,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2404_FFY_RST,
      O => rx_input_fifo_fifo_N2403
    );
  rx_input_fifo_fifo_N2404_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2404_FFY_RST
    );
  rx_input_memio_bp_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_4_FFY_RST
    );
  rx_input_memio_bp_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(5),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_4_FFY_RST,
      O => rx_input_memio_bp(5)
    );
  rx_input_memio_Msub_n0043_inst_cy_225_485 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_74,
      IB => rx_input_memio_bp_4_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_137,
      O => rx_input_memio_Msub_n0043_inst_cy_225
    );
  rx_input_memio_Msub_n0043_inst_sum_191 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_4_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_137,
      O => rx_input_memio_n0043(4)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1371 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_74,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_137
    );
  rx_input_memio_Msub_n0043_inst_lut2_1381 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_75,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_138
    );
  rx_input_memio_bp_4_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_4_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_226
    );
  rx_input_memio_Msub_n0043_inst_cy_226_486 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_75,
      IB => rx_input_memio_Msub_n0043_inst_cy_225,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_138,
      O => rx_input_memio_bp_4_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_192 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_225,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_138,
      O => rx_input_memio_n0043(5)
    );
  rx_input_memio_bp_4_CYINIT_487 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_224,
      O => rx_input_memio_bp_4_CYINIT
    );
  rx_input_memio_bp_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_6_FFY_RST
    );
  rx_input_memio_bp_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(7),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_6_FFY_RST,
      O => rx_input_memio_bp(7)
    );
  rx_input_memio_Msub_n0043_inst_cy_227_488 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_76,
      IB => rx_input_memio_bp_6_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_139,
      O => rx_input_memio_Msub_n0043_inst_cy_227
    );
  rx_input_memio_Msub_n0043_inst_sum_193 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_6_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_139,
      O => rx_input_memio_n0043(6)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1391 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_76,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_139
    );
  rx_input_memio_Msub_n0043_inst_lut2_1401 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_77,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_140
    );
  rx_input_memio_bp_6_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_6_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_228
    );
  rx_input_memio_Msub_n0043_inst_cy_228_489 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_77,
      IB => rx_input_memio_Msub_n0043_inst_cy_227,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_140,
      O => rx_input_memio_bp_6_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_194 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_227,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_140,
      O => rx_input_memio_n0043(7)
    );
  rx_input_memio_bp_6_CYINIT_490 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_226,
      O => rx_input_memio_bp_6_CYINIT
    );
  rx_input_memio_bp_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_8_FFY_RST
    );
  rx_input_memio_bp_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(9),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_8_FFY_RST,
      O => rx_input_memio_bp(9)
    );
  rx_input_memio_Msub_n0043_inst_cy_229_491 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_78,
      IB => rx_input_memio_bp_8_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_141,
      O => rx_input_memio_Msub_n0043_inst_cy_229
    );
  rx_input_memio_Msub_n0043_inst_sum_195 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_8_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_141,
      O => rx_input_memio_n0043(8)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1411 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_78,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_141
    );
  rx_input_memio_Msub_n0043_inst_lut2_1421 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_79,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_142
    );
  rx_input_memio_bp_8_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_8_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_230
    );
  rx_input_memio_Msub_n0043_inst_cy_230_492 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_79,
      IB => rx_input_memio_Msub_n0043_inst_cy_229,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_142,
      O => rx_input_memio_bp_8_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_196 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_229,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_142,
      O => rx_input_memio_n0043(9)
    );
  rx_input_memio_bp_8_CYINIT_493 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_228,
      O => rx_input_memio_bp_8_CYINIT
    );
  rx_input_memio_bp_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_10_FFY_RST
    );
  rx_input_memio_bp_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(11),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_10_FFY_RST,
      O => rx_input_memio_bp(11)
    );
  rx_input_memio_Msub_n0043_inst_cy_231_494 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_80,
      IB => rx_input_memio_bp_10_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_143,
      O => rx_input_memio_Msub_n0043_inst_cy_231
    );
  rx_input_memio_Msub_n0043_inst_sum_197 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_10_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_143,
      O => rx_input_memio_n0043(10)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1431 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_80,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_143
    );
  rx_input_memio_Msub_n0043_inst_lut2_1441 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_81,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_144
    );
  rx_input_memio_bp_10_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_10_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_232
    );
  rx_input_memio_Msub_n0043_inst_cy_232_495 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_81,
      IB => rx_input_memio_Msub_n0043_inst_cy_231,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_144,
      O => rx_input_memio_bp_10_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_198 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_231,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_144,
      O => rx_input_memio_n0043(11)
    );
  rx_input_memio_bp_10_CYINIT_496 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_230,
      O => rx_input_memio_bp_10_CYINIT
    );
  rx_input_memio_Msub_n0043_inst_cy_233_497 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_82,
      IB => rx_input_memio_bp_12_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_145,
      O => rx_input_memio_Msub_n0043_inst_cy_233
    );
  rx_input_memio_Msub_n0043_inst_sum_199 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_12_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_145,
      O => rx_input_memio_n0043(12)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1451 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_82,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_145
    );
  rx_input_memio_Msub_n0043_inst_lut2_1461 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_83,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_146
    );
  rx_input_memio_bp_12_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_12_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_234
    );
  rx_input_memio_Msub_n0043_inst_cy_234_498 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_83,
      IB => rx_input_memio_Msub_n0043_inst_cy_233,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_146,
      O => rx_input_memio_bp_12_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_200 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_233,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_146,
      O => rx_input_memio_n0043(13)
    );
  rx_input_memio_bp_12_CYINIT_499 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_232,
      O => rx_input_memio_bp_12_CYINIT
    );
  rx_input_memio_Msub_n0043_inst_cy_235_500 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_84,
      IB => rx_input_memio_bp_14_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_147,
      O => rx_input_memio_Msub_n0043_inst_cy_235
    );
  rx_input_memio_Msub_n0043_inst_sum_201 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_14_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_147,
      O => rx_input_memio_n0043(14)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1471 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_84,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_147
    );
  rx_input_memio_Msub_n0043_inst_lut2_1481 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_85,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_148
    );
  rx_input_memio_Msub_n0043_inst_sum_202 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_235,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_148,
      O => rx_input_memio_n0043(15)
    );
  rx_input_memio_bp_14_CYINIT_501 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_234,
      O => rx_input_memio_bp_14_CYINIT
    );
  mac_control_rxoferr_cnt_0_LOGIC_ZERO_502 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_0_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_16_503 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_33,
      IB => mac_control_rxoferr_cnt_0_LOGIC_ZERO,
      SEL => mac_control_rxoferr_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_33,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(0),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_rxoferr_cnt_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_16,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(1),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_0_GROM
    );
  mac_control_rxoferr_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_0_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_17_504 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_16,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_rxoferr_cnt_0_GROM,
      O => mac_control_rxoferr_cnt_0_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_rxoferr_cnt_0_GROM,
      O => mac_control_rxoferr_cnt_n0000(1)
    );
  mac_control_rxoferr_cnt_2_LOGIC_ZERO_505 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_2_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_18_506 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_2_CYINIT,
      SEL => mac_control_rxoferr_cnt_2_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_2_CYINIT,
      I1 => mac_control_rxoferr_cnt_2_FROM,
      O => mac_control_rxoferr_cnt_n0000(2)
    );
  mac_control_rxoferr_cnt_2_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxoferr_cnt(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_2_FROM
    );
  mac_control_rxoferr_cnt_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(3),
      O => mac_control_rxoferr_cnt_2_GROM
    );
  mac_control_rxoferr_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_2_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_19_507 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_rxoferr_cnt_2_GROM,
      O => mac_control_rxoferr_cnt_2_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_rxoferr_cnt_2_GROM,
      O => mac_control_rxoferr_cnt_n0000(3)
    );
  mac_control_rxoferr_cnt_2_CYINIT_508 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_rxoferr_cnt_2_CYINIT
    );
  mac_control_rxoferr_cnt_4_LOGIC_ZERO_509 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_4_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_20_510 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_4_CYINIT,
      SEL => mac_control_rxoferr_cnt_4_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_4_CYINIT,
      I1 => mac_control_rxoferr_cnt_4_FROM,
      O => mac_control_rxoferr_cnt_n0000(4)
    );
  mac_control_rxoferr_cnt_4_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(4),
      O => mac_control_rxoferr_cnt_4_FROM
    );
  mac_control_rxoferr_cnt_4_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(5),
      O => mac_control_rxoferr_cnt_4_GROM
    );
  mac_control_rxoferr_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_4_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_21_511 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_rxoferr_cnt_4_GROM,
      O => mac_control_rxoferr_cnt_4_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_rxoferr_cnt_4_GROM,
      O => mac_control_rxoferr_cnt_n0000(5)
    );
  mac_control_rxoferr_cnt_4_CYINIT_512 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_rxoferr_cnt_4_CYINIT
    );
  rx_input_fifo_fifo_BU71 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2808,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N19_FFY_RST,
      O => rx_input_fifo_fifo_N18
    );
  rx_input_fifo_fifo_N19_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N19_FFY_RST
    );
  mac_control_rxoferr_cnt_6_LOGIC_ZERO_513 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_6_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_22_514 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_6_CYINIT,
      SEL => mac_control_rxoferr_cnt_6_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_6_CYINIT,
      I1 => mac_control_rxoferr_cnt_6_FROM,
      O => mac_control_rxoferr_cnt_n0000(6)
    );
  mac_control_rxoferr_cnt_6_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxoferr_cnt(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_6_FROM
    );
  mac_control_rxoferr_cnt_6_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxoferr_cnt(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_6_GROM
    );
  mac_control_rxoferr_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_6_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_23_515 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_rxoferr_cnt_6_GROM,
      O => mac_control_rxoferr_cnt_6_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_rxoferr_cnt_6_GROM,
      O => mac_control_rxoferr_cnt_n0000(7)
    );
  mac_control_rxoferr_cnt_6_CYINIT_516 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_rxoferr_cnt_6_CYINIT
    );
  mac_control_rxoferr_cnt_8_LOGIC_ZERO_517 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_8_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_24_518 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_8_CYINIT,
      SEL => mac_control_rxoferr_cnt_8_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_8_CYINIT,
      I1 => mac_control_rxoferr_cnt_8_FROM,
      O => mac_control_rxoferr_cnt_n0000(8)
    );
  mac_control_rxoferr_cnt_8_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(8),
      O => mac_control_rxoferr_cnt_8_FROM
    );
  mac_control_rxoferr_cnt_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(9),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_8_GROM
    );
  mac_control_rxoferr_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_8_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_25_519 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_rxoferr_cnt_8_GROM,
      O => mac_control_rxoferr_cnt_8_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_rxoferr_cnt_8_GROM,
      O => mac_control_rxoferr_cnt_n0000(9)
    );
  mac_control_rxoferr_cnt_8_CYINIT_520 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_rxoferr_cnt_8_CYINIT
    );
  mac_control_rxoferr_cnt_10_LOGIC_ZERO_521 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_10_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_26_522 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_10_CYINIT,
      SEL => mac_control_rxoferr_cnt_10_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_10_CYINIT,
      I1 => mac_control_rxoferr_cnt_10_FROM,
      O => mac_control_rxoferr_cnt_n0000(10)
    );
  mac_control_rxoferr_cnt_10_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(10),
      O => mac_control_rxoferr_cnt_10_FROM
    );
  mac_control_rxoferr_cnt_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(11),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_10_GROM
    );
  mac_control_rxoferr_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_10_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_27_523 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_rxoferr_cnt_10_GROM,
      O => mac_control_rxoferr_cnt_10_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_rxoferr_cnt_10_GROM,
      O => mac_control_rxoferr_cnt_n0000(11)
    );
  mac_control_rxoferr_cnt_10_CYINIT_524 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_rxoferr_cnt_10_CYINIT
    );
  mac_control_rxoferr_cnt_12_LOGIC_ZERO_525 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_12_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_28_526 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_12_CYINIT,
      SEL => mac_control_rxoferr_cnt_12_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_12_CYINIT,
      I1 => mac_control_rxoferr_cnt_12_FROM,
      O => mac_control_rxoferr_cnt_n0000(12)
    );
  mac_control_rxoferr_cnt_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxoferr_cnt(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_12_FROM
    );
  mac_control_rxoferr_cnt_12_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxoferr_cnt(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_12_GROM
    );
  mac_control_rxoferr_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_12_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_29_527 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_rxoferr_cnt_12_GROM,
      O => mac_control_rxoferr_cnt_12_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_rxoferr_cnt_12_GROM,
      O => mac_control_rxoferr_cnt_n0000(13)
    );
  mac_control_rxoferr_cnt_12_CYINIT_528 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_rxoferr_cnt_12_CYINIT
    );
  mac_control_rxoferr_cnt_14_LOGIC_ZERO_529 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_14_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_30_530 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_14_CYINIT,
      SEL => mac_control_rxoferr_cnt_14_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_14_CYINIT,
      I1 => mac_control_rxoferr_cnt_14_FROM,
      O => mac_control_rxoferr_cnt_n0000(14)
    );
  mac_control_rxoferr_cnt_14_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(14),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_14_FROM
    );
  mac_control_rxoferr_cnt_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(15),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_14_GROM
    );
  mac_control_rxoferr_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_14_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_31_531 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_rxoferr_cnt_14_GROM,
      O => mac_control_rxoferr_cnt_14_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_rxoferr_cnt_14_GROM,
      O => mac_control_rxoferr_cnt_n0000(15)
    );
  mac_control_rxoferr_cnt_14_CYINIT_532 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_rxoferr_cnt_14_CYINIT
    );
  mac_control_rxoferr_cnt_16_LOGIC_ZERO_533 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_16_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_32_534 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_16_CYINIT,
      SEL => mac_control_rxoferr_cnt_16_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_16_CYINIT,
      I1 => mac_control_rxoferr_cnt_16_FROM,
      O => mac_control_rxoferr_cnt_n0000(16)
    );
  mac_control_rxoferr_cnt_16_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(16),
      O => mac_control_rxoferr_cnt_16_FROM
    );
  mac_control_rxoferr_cnt_16_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(17),
      O => mac_control_rxoferr_cnt_16_GROM
    );
  mac_control_rxoferr_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_16_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_33_535 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_rxoferr_cnt_16_GROM,
      O => mac_control_rxoferr_cnt_16_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_rxoferr_cnt_16_GROM,
      O => mac_control_rxoferr_cnt_n0000(17)
    );
  mac_control_rxoferr_cnt_16_CYINIT_536 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_rxoferr_cnt_16_CYINIT
    );
  mac_control_rxoferr_cnt_18_LOGIC_ZERO_537 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_18_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_34_538 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_18_CYINIT,
      SEL => mac_control_rxoferr_cnt_18_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_18_CYINIT,
      I1 => mac_control_rxoferr_cnt_18_FROM,
      O => mac_control_rxoferr_cnt_n0000(18)
    );
  mac_control_rxoferr_cnt_18_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(18),
      O => mac_control_rxoferr_cnt_18_FROM
    );
  mac_control_rxoferr_cnt_18_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(19),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_18_GROM
    );
  mac_control_rxoferr_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_18_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_35_539 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_rxoferr_cnt_18_GROM,
      O => mac_control_rxoferr_cnt_18_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_rxoferr_cnt_18_GROM,
      O => mac_control_rxoferr_cnt_n0000(19)
    );
  mac_control_rxoferr_cnt_18_CYINIT_540 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_rxoferr_cnt_18_CYINIT
    );
  mac_control_rxoferr_cnt_20_LOGIC_ZERO_541 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_20_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_36_542 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_20_CYINIT,
      SEL => mac_control_rxoferr_cnt_20_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_20_CYINIT,
      I1 => mac_control_rxoferr_cnt_20_FROM,
      O => mac_control_rxoferr_cnt_n0000(20)
    );
  mac_control_rxoferr_cnt_20_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(20),
      O => mac_control_rxoferr_cnt_20_FROM
    );
  mac_control_rxoferr_cnt_20_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(21),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_20_GROM
    );
  mac_control_rxoferr_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_20_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_37_543 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_rxoferr_cnt_20_GROM,
      O => mac_control_rxoferr_cnt_20_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_rxoferr_cnt_20_GROM,
      O => mac_control_rxoferr_cnt_n0000(21)
    );
  mac_control_rxoferr_cnt_20_CYINIT_544 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_rxoferr_cnt_20_CYINIT
    );
  mac_control_rxoferr_cnt_22_LOGIC_ZERO_545 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_22_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_38_546 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_22_CYINIT,
      SEL => mac_control_rxoferr_cnt_22_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_22_CYINIT,
      I1 => mac_control_rxoferr_cnt_22_FROM,
      O => mac_control_rxoferr_cnt_n0000(22)
    );
  mac_control_rxoferr_cnt_22_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(22),
      O => mac_control_rxoferr_cnt_22_FROM
    );
  mac_control_rxoferr_cnt_22_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(23),
      O => mac_control_rxoferr_cnt_22_GROM
    );
  mac_control_rxoferr_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_22_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_39_547 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_rxoferr_cnt_22_GROM,
      O => mac_control_rxoferr_cnt_22_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_rxoferr_cnt_22_GROM,
      O => mac_control_rxoferr_cnt_n0000(23)
    );
  mac_control_rxoferr_cnt_22_CYINIT_548 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_rxoferr_cnt_22_CYINIT
    );
  mac_control_rxoferr_cnt_24_LOGIC_ZERO_549 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_24_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_40_550 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_24_CYINIT,
      SEL => mac_control_rxoferr_cnt_24_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_24_CYINIT,
      I1 => mac_control_rxoferr_cnt_24_FROM,
      O => mac_control_rxoferr_cnt_n0000(24)
    );
  mac_control_rxoferr_cnt_24_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(24),
      O => mac_control_rxoferr_cnt_24_FROM
    );
  mac_control_rxoferr_cnt_24_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(25),
      O => mac_control_rxoferr_cnt_24_GROM
    );
  mac_control_rxoferr_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_24_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_41_551 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_rxoferr_cnt_24_GROM,
      O => mac_control_rxoferr_cnt_24_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_rxoferr_cnt_24_GROM,
      O => mac_control_rxoferr_cnt_n0000(25)
    );
  mac_control_rxoferr_cnt_24_CYINIT_552 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_rxoferr_cnt_24_CYINIT
    );
  rx_input_fifo_fifo_BU199 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2482,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2502_FFX_RST,
      O => rx_input_fifo_fifo_N2502
    );
  rx_input_fifo_fifo_N2502_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2502_FFX_RST
    );
  mac_control_rxoferr_cnt_26_LOGIC_ZERO_553 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_26_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_42_554 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_26_CYINIT,
      SEL => mac_control_rxoferr_cnt_26_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_26_CYINIT,
      I1 => mac_control_rxoferr_cnt_26_FROM,
      O => mac_control_rxoferr_cnt_n0000(26)
    );
  mac_control_rxoferr_cnt_26_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(26),
      O => mac_control_rxoferr_cnt_26_FROM
    );
  mac_control_rxoferr_cnt_26_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(27),
      O => mac_control_rxoferr_cnt_26_GROM
    );
  mac_control_rxoferr_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_26_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_43_555 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_rxoferr_cnt_26_GROM,
      O => mac_control_rxoferr_cnt_26_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_rxoferr_cnt_26_GROM,
      O => mac_control_rxoferr_cnt_n0000(27)
    );
  mac_control_rxoferr_cnt_26_CYINIT_556 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_rxoferr_cnt_26_CYINIT
    );
  mac_control_rxoferr_cnt_28_LOGIC_ZERO_557 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_28_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_44_558 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_28_CYINIT,
      SEL => mac_control_rxoferr_cnt_28_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_28_CYINIT,
      I1 => mac_control_rxoferr_cnt_28_FROM,
      O => mac_control_rxoferr_cnt_n0000(28)
    );
  mac_control_rxoferr_cnt_28_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(28),
      O => mac_control_rxoferr_cnt_28_FROM
    );
  mac_control_rxoferr_cnt_28_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(29),
      O => mac_control_rxoferr_cnt_28_GROM
    );
  mac_control_rxoferr_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_28_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_45_559 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_rxoferr_cnt_28_GROM,
      O => mac_control_rxoferr_cnt_28_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_rxoferr_cnt_28_GROM,
      O => mac_control_rxoferr_cnt_n0000(29)
    );
  mac_control_rxoferr_cnt_28_CYINIT_560 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_rxoferr_cnt_28_CYINIT
    );
  mac_control_rxoferr_cnt_30_LOGIC_ZERO_561 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_30_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_46_562 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_30_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_30_CYINIT,
      SEL => mac_control_rxoferr_cnt_30_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_30_CYINIT,
      I1 => mac_control_rxoferr_cnt_30_FROM,
      O => mac_control_rxoferr_cnt_n0000(30)
    );
  mac_control_rxoferr_cnt_30_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(30),
      O => mac_control_rxoferr_cnt_30_FROM
    );
  mac_control_rxoferr_cnt_31_rt_563 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(31),
      O => mac_control_rxoferr_cnt_31_rt
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_rxoferr_cnt_31_rt,
      O => mac_control_rxoferr_cnt_n0000(31)
    );
  mac_control_rxoferr_cnt_30_CYINIT_564 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_rxoferr_cnt_30_CYINIT
    );
  mac_control_ledrx_cnt_154_LOGIC_ONE_565 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_154_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_340_566 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_21,
      IB => mac_control_ledrx_cnt_154_LOGIC_ONE,
      SEL => mac_control_ledrx_rst_rt,
      O => mac_control_ledrx_cnt_inst_cy_340
    );
  mac_control_ledrx_rst_rt_567 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_21,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_rst,
      ADR3 => VCC,
      O => mac_control_ledrx_rst_rt
    );
  mac_control_ledrx_cnt_inst_lut3_2361 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_28,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_cnt_154,
      ADR3 => mac_control_ledrx_rst,
      O => mac_control_ledrx_cnt_inst_lut3_236
    );
  mac_control_ledrx_cnt_154_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_154_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_341
    );
  mac_control_ledrx_cnt_inst_cy_341_568 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_28,
      IB => mac_control_ledrx_cnt_inst_cy_340,
      SEL => mac_control_ledrx_cnt_inst_lut3_236,
      O => mac_control_ledrx_cnt_154_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_301_569 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_340,
      I1 => mac_control_ledrx_cnt_inst_lut3_236,
      O => mac_control_ledrx_cnt_inst_sum_301
    );
  mac_control_ledrx_cnt_155_LOGIC_ONE_570 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_155_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_342_571 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_155_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_155_CYINIT,
      SEL => mac_control_ledrx_cnt_inst_lut3_237,
      O => mac_control_ledrx_cnt_inst_cy_342
    );
  mac_control_ledrx_cnt_inst_sum_302_572 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_155_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_237,
      O => mac_control_ledrx_cnt_inst_sum_302
    );
  mac_control_ledrx_cnt_inst_lut3_2371 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_ledrx_rst,
      ADR1 => mac_control_ledrx_cnt_155,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledrx_cnt_inst_lut3_237
    );
  mac_control_ledrx_cnt_inst_lut3_2381 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_rst,
      ADR3 => mac_control_ledrx_cnt_156,
      O => mac_control_ledrx_cnt_inst_lut3_238
    );
  mac_control_ledrx_cnt_155_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_155_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_343
    );
  mac_control_ledrx_cnt_inst_cy_343_573 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_155_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_inst_cy_342,
      SEL => mac_control_ledrx_cnt_inst_lut3_238,
      O => mac_control_ledrx_cnt_155_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_303_574 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_342,
      I1 => mac_control_ledrx_cnt_inst_lut3_238,
      O => mac_control_ledrx_cnt_inst_sum_303
    );
  mac_control_ledrx_cnt_155_CYINIT_575 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_341,
      O => mac_control_ledrx_cnt_155_CYINIT
    );
  mac_control_ledrx_cnt_157_LOGIC_ONE_576 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_157_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_344_577 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_157_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_157_CYINIT,
      SEL => mac_control_ledrx_cnt_inst_lut3_239,
      O => mac_control_ledrx_cnt_inst_cy_344
    );
  mac_control_ledrx_cnt_inst_sum_304_578 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_157_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_239,
      O => mac_control_ledrx_cnt_inst_sum_304
    );
  mac_control_ledrx_cnt_inst_lut3_2391 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_cnt_157,
      ADR3 => mac_control_ledrx_rst,
      O => mac_control_ledrx_cnt_inst_lut3_239
    );
  mac_control_ledrx_cnt_inst_lut3_2401 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledrx_cnt_158,
      ADR2 => VCC,
      ADR3 => mac_control_ledrx_rst,
      O => mac_control_ledrx_cnt_inst_lut3_240
    );
  mac_control_ledrx_cnt_157_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_157_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_345
    );
  mac_control_ledrx_cnt_inst_cy_345_579 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_157_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_inst_cy_344,
      SEL => mac_control_ledrx_cnt_inst_lut3_240,
      O => mac_control_ledrx_cnt_157_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_305_580 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_344,
      I1 => mac_control_ledrx_cnt_inst_lut3_240,
      O => mac_control_ledrx_cnt_inst_sum_305
    );
  mac_control_ledrx_cnt_157_CYINIT_581 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_343,
      O => mac_control_ledrx_cnt_157_CYINIT
    );
  mac_control_ledrx_cnt_159_LOGIC_ONE_582 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_159_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_346_583 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_159_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_159_CYINIT,
      SEL => mac_control_ledrx_cnt_inst_lut3_241,
      O => mac_control_ledrx_cnt_inst_cy_346
    );
  mac_control_ledrx_cnt_inst_sum_306_584 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_159_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_241,
      O => mac_control_ledrx_cnt_inst_sum_306
    );
  mac_control_ledrx_cnt_inst_lut3_2411 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledrx_rst,
      ADR2 => VCC,
      ADR3 => mac_control_ledrx_cnt_159,
      O => mac_control_ledrx_cnt_inst_lut3_241
    );
  mac_control_ledrx_cnt_inst_lut3_2421 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_160,
      ADR1 => mac_control_ledrx_rst,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledrx_cnt_inst_lut3_242
    );
  mac_control_ledrx_cnt_159_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_159_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_347
    );
  mac_control_ledrx_cnt_inst_cy_347_585 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_159_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_inst_cy_346,
      SEL => mac_control_ledrx_cnt_inst_lut3_242,
      O => mac_control_ledrx_cnt_159_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_307_586 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_346,
      I1 => mac_control_ledrx_cnt_inst_lut3_242,
      O => mac_control_ledrx_cnt_inst_sum_307
    );
  mac_control_ledrx_cnt_159_CYINIT_587 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_345,
      O => mac_control_ledrx_cnt_159_CYINIT
    );
  mac_control_ledrx_cnt_161_LOGIC_ONE_588 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_161_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_348_589 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_161_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_161_CYINIT,
      SEL => mac_control_ledrx_cnt_inst_lut3_243,
      O => mac_control_ledrx_cnt_inst_cy_348
    );
  mac_control_ledrx_cnt_inst_sum_308_590 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_161_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_243,
      O => mac_control_ledrx_cnt_inst_sum_308
    );
  mac_control_ledrx_cnt_inst_lut3_2431 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledrx_rst,
      ADR2 => VCC,
      ADR3 => mac_control_ledrx_cnt_161,
      O => mac_control_ledrx_cnt_inst_lut3_243
    );
  mac_control_ledrx_cnt_inst_lut3_2441 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_162,
      ADR1 => mac_control_ledrx_rst,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledrx_cnt_inst_lut3_244
    );
  mac_control_ledrx_cnt_161_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_161_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_349
    );
  mac_control_ledrx_cnt_inst_cy_349_591 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_161_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_inst_cy_348,
      SEL => mac_control_ledrx_cnt_inst_lut3_244,
      O => mac_control_ledrx_cnt_161_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_309_592 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_348,
      I1 => mac_control_ledrx_cnt_inst_lut3_244,
      O => mac_control_ledrx_cnt_inst_sum_309
    );
  mac_control_ledrx_cnt_161_CYINIT_593 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_347,
      O => mac_control_ledrx_cnt_161_CYINIT
    );
  mac_control_ledrx_cnt_163_LOGIC_ONE_594 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_163_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_350_595 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_163_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_163_CYINIT,
      SEL => mac_control_ledrx_cnt_inst_lut3_245,
      O => mac_control_ledrx_cnt_inst_cy_350
    );
  mac_control_ledrx_cnt_inst_sum_310_596 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_163_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_245,
      O => mac_control_ledrx_cnt_inst_sum_310
    );
  mac_control_ledrx_cnt_inst_lut3_2451 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_cnt_163,
      ADR3 => mac_control_ledrx_rst,
      O => mac_control_ledrx_cnt_inst_lut3_245
    );
  mac_control_ledrx_cnt_inst_lut3_2461 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_rst,
      ADR3 => mac_control_ledrx_cnt_164,
      O => mac_control_ledrx_cnt_inst_lut3_246
    );
  mac_control_ledrx_cnt_163_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_163_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_351
    );
  mac_control_ledrx_cnt_inst_cy_351_597 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_163_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_inst_cy_350,
      SEL => mac_control_ledrx_cnt_inst_lut3_246,
      O => mac_control_ledrx_cnt_163_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_311_598 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_350,
      I1 => mac_control_ledrx_cnt_inst_lut3_246,
      O => mac_control_ledrx_cnt_inst_sum_311
    );
  mac_control_ledrx_cnt_163_CYINIT_599 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_349,
      O => mac_control_ledrx_cnt_163_CYINIT
    );
  mac_control_ledrx_cnt_inst_sum_312_600 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_165_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_247,
      O => mac_control_ledrx_cnt_inst_sum_312
    );
  mac_control_ledrx_cnt_inst_lut3_2471 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_165,
      ADR1 => mac_control_ledrx_rst,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledrx_cnt_inst_lut3_247
    );
  mac_control_ledrx_cnt_165_CYINIT_601 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_351,
      O => mac_control_ledrx_cnt_165_CYINIT
    );
  tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ONE_602 : X_ONE
    port map (
      O => tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ONE
    );
  tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ZERO_603 : X_ZERO
    port map (
      O => tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ZERO
    );
  tx_output_Mcompar_n0035_inst_cy_194_604 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ONE,
      SEL => tx_output_bcntl_1_rt,
      O => tx_output_Mcompar_n0035_inst_cy_194
    );
  tx_output_bcntl_1_rt_605 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_bcntl(1),
      ADR3 => VCC,
      O => tx_output_bcntl_1_rt
    );
  tx_output_BEL_0 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_bcntl(1),
      O => tx_output_SIG_25
    );
  tx_output_Mcompar_n0035_inst_cy_195_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_195_CYMUXG,
      O => tx_output_Mcompar_n0035_inst_cy_195
    );
  tx_output_Mcompar_n0035_inst_cy_195_606 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0035_inst_cy_194,
      SEL => tx_output_SIG_25,
      O => tx_output_Mcompar_n0035_inst_cy_195_CYMUXG
    );
  tx_output_Mcompar_n0035_inst_cy_197_LOGIC_ONE_607 : X_ONE
    port map (
      O => tx_output_Mcompar_n0035_inst_cy_197_LOGIC_ONE
    );
  tx_output_Mcompar_n0035_inst_cy_196_608 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_197_LOGIC_ONE,
      IB => tx_output_Mcompar_n0035_inst_cy_197_CYINIT,
      SEL => tx_output_Mcompar_n0035_inst_lut1_6,
      O => tx_output_Mcompar_n0035_inst_cy_196
    );
  tx_output_Mcompar_n0035_inst_lut1_61 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_bcntl(2),
      ADR3 => VCC,
      O => tx_output_Mcompar_n0035_inst_lut1_6
    );
  tx_output_Mcompar_n0035_inst_lut1_71 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_bcntl(2),
      ADR3 => VCC,
      O => tx_output_Mcompar_n0035_inst_lut1_7
    );
  tx_output_Mcompar_n0035_inst_cy_197_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_197_CYMUXG,
      O => tx_output_Mcompar_n0035_inst_cy_197
    );
  tx_output_Mcompar_n0035_inst_cy_197_609 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_197_LOGIC_ONE,
      IB => tx_output_Mcompar_n0035_inst_cy_196,
      SEL => tx_output_Mcompar_n0035_inst_lut1_7,
      O => tx_output_Mcompar_n0035_inst_cy_197_CYMUXG
    );
  tx_output_Mcompar_n0035_inst_cy_197_CYINIT_610 : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_195,
      O => tx_output_Mcompar_n0035_inst_cy_197_CYINIT
    );
  tx_output_Mcompar_n0035_inst_cy_199_LOGIC_ZERO_611 : X_ZERO
    port map (
      O => tx_output_Mcompar_n0035_inst_cy_199_LOGIC_ZERO
    );
  tx_output_Mcompar_n0035_inst_cy_198_612 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_199_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0035_inst_cy_199_CYINIT,
      SEL => tx_output_bcntl_3_rt,
      O => tx_output_Mcompar_n0035_inst_cy_198
    );
  tx_output_bcntl_3_rt_613 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_bcntl(3),
      ADR3 => VCC,
      O => tx_output_bcntl_3_rt
    );
  tx_output_BEL_1 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_bcntl(3),
      ADR3 => VCC,
      O => tx_output_SIG_26
    );
  tx_output_Mcompar_n0035_inst_cy_199_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_199_CYMUXG,
      O => tx_output_Mcompar_n0035_inst_cy_199
    );
  tx_output_Mcompar_n0035_inst_cy_199_614 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_199_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0035_inst_cy_198,
      SEL => tx_output_SIG_26,
      O => tx_output_Mcompar_n0035_inst_cy_199_CYMUXG
    );
  tx_output_Mcompar_n0035_inst_cy_199_CYINIT_615 : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_197,
      O => tx_output_Mcompar_n0035_inst_cy_199_CYINIT
    );
  tx_output_Mcompar_n0035_inst_cy_201_LOGIC_ONE_616 : X_ONE
    port map (
      O => tx_output_Mcompar_n0035_inst_cy_201_LOGIC_ONE
    );
  tx_output_Mcompar_n0035_inst_cy_200_617 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_201_LOGIC_ONE,
      IB => tx_output_Mcompar_n0035_inst_cy_201_CYINIT,
      SEL => tx_output_Mcompar_n0035_inst_lut4_16,
      O => tx_output_Mcompar_n0035_inst_cy_200
    );
  tx_output_Mcompar_n0035_inst_lut4_161 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcntl(6),
      ADR1 => tx_output_bcntl(5),
      ADR2 => tx_output_bcntl(4),
      ADR3 => tx_output_bcntl(7),
      O => tx_output_Mcompar_n0035_inst_lut4_16
    );
  tx_output_Mcompar_n0035_inst_lut4_171 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcntl(6),
      ADR1 => tx_output_bcntl(5),
      ADR2 => tx_output_bcntl(4),
      ADR3 => tx_output_bcntl(7),
      O => tx_output_Mcompar_n0035_inst_lut4_17
    );
  tx_output_Mcompar_n0035_inst_cy_201_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_201_CYMUXG,
      O => tx_output_Mcompar_n0035_inst_cy_201
    );
  tx_output_Mcompar_n0035_inst_cy_201_618 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_201_LOGIC_ONE,
      IB => tx_output_Mcompar_n0035_inst_cy_200,
      SEL => tx_output_Mcompar_n0035_inst_lut4_17,
      O => tx_output_Mcompar_n0035_inst_cy_201_CYMUXG
    );
  tx_output_Mcompar_n0035_inst_cy_201_CYINIT_619 : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_199,
      O => tx_output_Mcompar_n0035_inst_cy_201_CYINIT
    );
  rx_input_fifo_fifo_BU129 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3320,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2404_FFX_RST,
      O => rx_input_fifo_fifo_N2404
    );
  rx_input_fifo_fifo_N2404_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2404_FFX_RST
    );
  tx_output_n0035_LOGIC_ONE_620 : X_ONE
    port map (
      O => tx_output_n0035_LOGIC_ONE
    );
  tx_output_Mcompar_n0035_inst_cy_202_621 : X_MUX2
    port map (
      IA => tx_output_n0035_LOGIC_ONE,
      IB => tx_output_n0035_CYINIT,
      SEL => tx_output_Mcompar_n0035_inst_lut4_18,
      O => tx_output_Mcompar_n0035_inst_cy_202
    );
  tx_output_Mcompar_n0035_inst_lut4_181 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcntl(9),
      ADR1 => tx_output_bcntl(11),
      ADR2 => tx_output_bcntl(10),
      ADR3 => tx_output_bcntl(8),
      O => tx_output_Mcompar_n0035_inst_lut4_18
    );
  tx_output_Mcompar_n0035_inst_lut4_191 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcntl(15),
      ADR1 => tx_output_bcntl(12),
      ADR2 => tx_output_bcntl(14),
      ADR3 => tx_output_bcntl(13),
      O => tx_output_Mcompar_n0035_inst_lut4_19
    );
  tx_output_n0035_COUTUSED : X_BUF
    port map (
      I => tx_output_n0035_CYMUXG,
      O => tx_output_n0035
    );
  tx_output_Mcompar_n0035_inst_cy_203 : X_MUX2
    port map (
      IA => tx_output_n0035_LOGIC_ONE,
      IB => tx_output_Mcompar_n0035_inst_cy_202,
      SEL => tx_output_Mcompar_n0035_inst_lut4_19,
      O => tx_output_n0035_CYMUXG
    );
  tx_output_n0035_CYINIT_622 : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_201,
      O => tx_output_n0035_CYINIT
    );
  mac_control_rxphyerr_cnt_0_LOGIC_ZERO_623 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_0_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_16_624 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_33,
      IB => mac_control_rxphyerr_cnt_0_LOGIC_ZERO,
      SEL => mac_control_rxphyerr_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_33,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(0),
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_rxphyerr_cnt_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_16,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(1),
      O => mac_control_rxphyerr_cnt_0_GROM
    );
  mac_control_rxphyerr_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_0_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_17_625 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_16,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_rxphyerr_cnt_0_GROM,
      O => mac_control_rxphyerr_cnt_0_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_rxphyerr_cnt_0_GROM,
      O => mac_control_rxphyerr_cnt_n0000(1)
    );
  rx_input_fifo_fifo_BU193 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2484,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2504_FFY_RST,
      O => rx_input_fifo_fifo_N2504
    );
  rx_input_fifo_fifo_N2504_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2504_FFY_RST
    );
  mac_control_rxphyerr_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(3),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(3)
    );
  mac_control_rxphyerr_cnt_2_LOGIC_ZERO_626 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_2_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_18_627 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_2_CYINIT,
      SEL => mac_control_rxphyerr_cnt_2_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_2_CYINIT,
      I1 => mac_control_rxphyerr_cnt_2_FROM,
      O => mac_control_rxphyerr_cnt_n0000(2)
    );
  mac_control_rxphyerr_cnt_2_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(2),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_2_FROM
    );
  mac_control_rxphyerr_cnt_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(3),
      O => mac_control_rxphyerr_cnt_2_GROM
    );
  mac_control_rxphyerr_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_2_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_19_628 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_rxphyerr_cnt_2_GROM,
      O => mac_control_rxphyerr_cnt_2_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_rxphyerr_cnt_2_GROM,
      O => mac_control_rxphyerr_cnt_n0000(3)
    );
  mac_control_rxphyerr_cnt_2_CYINIT_629 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_rxphyerr_cnt_2_CYINIT
    );
  mac_control_rxphyerr_cnt_4_LOGIC_ZERO_630 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_4_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_20_631 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_4_CYINIT,
      SEL => mac_control_rxphyerr_cnt_4_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_4_CYINIT,
      I1 => mac_control_rxphyerr_cnt_4_FROM,
      O => mac_control_rxphyerr_cnt_n0000(4)
    );
  mac_control_rxphyerr_cnt_4_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(4),
      O => mac_control_rxphyerr_cnt_4_FROM
    );
  mac_control_rxphyerr_cnt_4_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(5),
      O => mac_control_rxphyerr_cnt_4_GROM
    );
  mac_control_rxphyerr_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_4_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_21_632 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_rxphyerr_cnt_4_GROM,
      O => mac_control_rxphyerr_cnt_4_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_rxphyerr_cnt_4_GROM,
      O => mac_control_rxphyerr_cnt_n0000(5)
    );
  mac_control_rxphyerr_cnt_4_CYINIT_633 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_rxphyerr_cnt_4_CYINIT
    );
  mac_control_rxphyerr_cnt_6_LOGIC_ZERO_634 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_6_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_22_635 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_6_CYINIT,
      SEL => mac_control_rxphyerr_cnt_6_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_6_CYINIT,
      I1 => mac_control_rxphyerr_cnt_6_FROM,
      O => mac_control_rxphyerr_cnt_n0000(6)
    );
  mac_control_rxphyerr_cnt_6_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(6),
      O => mac_control_rxphyerr_cnt_6_FROM
    );
  mac_control_rxphyerr_cnt_6_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(7),
      O => mac_control_rxphyerr_cnt_6_GROM
    );
  mac_control_rxphyerr_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_6_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_23_636 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_rxphyerr_cnt_6_GROM,
      O => mac_control_rxphyerr_cnt_6_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_rxphyerr_cnt_6_GROM,
      O => mac_control_rxphyerr_cnt_n0000(7)
    );
  mac_control_rxphyerr_cnt_6_CYINIT_637 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_rxphyerr_cnt_6_CYINIT
    );
  mac_control_rxphyerr_cnt_8_LOGIC_ZERO_638 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_8_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_24_639 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_8_CYINIT,
      SEL => mac_control_rxphyerr_cnt_8_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_8_CYINIT,
      I1 => mac_control_rxphyerr_cnt_8_FROM,
      O => mac_control_rxphyerr_cnt_n0000(8)
    );
  mac_control_rxphyerr_cnt_8_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(8),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_8_FROM
    );
  mac_control_rxphyerr_cnt_8_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_8_GROM
    );
  mac_control_rxphyerr_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_8_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_25_640 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_rxphyerr_cnt_8_GROM,
      O => mac_control_rxphyerr_cnt_8_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_rxphyerr_cnt_8_GROM,
      O => mac_control_rxphyerr_cnt_n0000(9)
    );
  mac_control_rxphyerr_cnt_8_CYINIT_641 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_rxphyerr_cnt_8_CYINIT
    );
  mac_control_rxphyerr_cnt_10_LOGIC_ZERO_642 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_10_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_26_643 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_10_CYINIT,
      SEL => mac_control_rxphyerr_cnt_10_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_10_CYINIT,
      I1 => mac_control_rxphyerr_cnt_10_FROM,
      O => mac_control_rxphyerr_cnt_n0000(10)
    );
  mac_control_rxphyerr_cnt_10_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(10),
      O => mac_control_rxphyerr_cnt_10_FROM
    );
  mac_control_rxphyerr_cnt_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(11),
      O => mac_control_rxphyerr_cnt_10_GROM
    );
  mac_control_rxphyerr_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_10_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_27_644 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_rxphyerr_cnt_10_GROM,
      O => mac_control_rxphyerr_cnt_10_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_rxphyerr_cnt_10_GROM,
      O => mac_control_rxphyerr_cnt_n0000(11)
    );
  mac_control_rxphyerr_cnt_10_CYINIT_645 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_rxphyerr_cnt_10_CYINIT
    );
  mac_control_rxphyerr_cnt_12_LOGIC_ZERO_646 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_12_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_28_647 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_12_CYINIT,
      SEL => mac_control_rxphyerr_cnt_12_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_12_CYINIT,
      I1 => mac_control_rxphyerr_cnt_12_FROM,
      O => mac_control_rxphyerr_cnt_n0000(12)
    );
  mac_control_rxphyerr_cnt_12_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(12),
      O => mac_control_rxphyerr_cnt_12_FROM
    );
  mac_control_rxphyerr_cnt_12_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_12_GROM
    );
  mac_control_rxphyerr_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_12_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_29_648 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_rxphyerr_cnt_12_GROM,
      O => mac_control_rxphyerr_cnt_12_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_rxphyerr_cnt_12_GROM,
      O => mac_control_rxphyerr_cnt_n0000(13)
    );
  mac_control_rxphyerr_cnt_12_CYINIT_649 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_rxphyerr_cnt_12_CYINIT
    );
  mac_control_rxphyerr_cnt_14_LOGIC_ZERO_650 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_14_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_30_651 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_14_CYINIT,
      SEL => mac_control_rxphyerr_cnt_14_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_14_CYINIT,
      I1 => mac_control_rxphyerr_cnt_14_FROM,
      O => mac_control_rxphyerr_cnt_n0000(14)
    );
  mac_control_rxphyerr_cnt_14_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(14),
      O => mac_control_rxphyerr_cnt_14_FROM
    );
  mac_control_rxphyerr_cnt_14_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(15),
      O => mac_control_rxphyerr_cnt_14_GROM
    );
  mac_control_rxphyerr_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_14_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_31_652 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_rxphyerr_cnt_14_GROM,
      O => mac_control_rxphyerr_cnt_14_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_rxphyerr_cnt_14_GROM,
      O => mac_control_rxphyerr_cnt_n0000(15)
    );
  mac_control_rxphyerr_cnt_14_CYINIT_653 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_rxphyerr_cnt_14_CYINIT
    );
  memcontroller_dnout_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_30_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_30_OFF_RST,
      O => memcontroller_dnout(30)
    );
  MD_30_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_30_OFF_RST
    );
  memcontroller_ts_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_30_TFF_RST,
      O => memcontroller_ts(30)
    );
  MD_30_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_30_TFF_RST
    );
  memcontroller_qn_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(23),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_23_IFF_RST,
      O => memcontroller_qn(23)
    );
  MD_23_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_23_IFF_RST
    );
  memcontroller_dnout_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_23_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_23_OFF_RST,
      O => memcontroller_dnout(23)
    );
  MD_23_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_23_OFF_RST
    );
  memcontroller_ts_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_23_TFF_RST,
      O => memcontroller_ts(23)
    );
  MD_23_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_23_TFF_RST
    );
  memcontroller_qn_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_15_IFF_RST,
      O => memcontroller_qn(15)
    );
  MD_15_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_15_IFF_RST
    );
  memcontroller_qn_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(31),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_31_IFF_RST,
      O => memcontroller_qn(31)
    );
  MD_31_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_31_IFF_RST
    );
  memcontroller_dnout_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_15_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_15_OFF_RST,
      O => memcontroller_dnout(15)
    );
  MD_15_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_15_OFF_RST
    );
  memcontroller_ts_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_15_TFF_RST,
      O => memcontroller_ts(15)
    );
  MD_15_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_15_TFF_RST
    );
  tx_input_dinl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_3_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_3_IFF_RST,
      O => tx_input_dinl(3)
    );
  DIN_3_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_3_IFF_RST
    );
  tx_input_dinl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_4_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_4_IFF_RST,
      O => tx_input_dinl(4)
    );
  DIN_4_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_4_IFF_RST
    );
  tx_input_dinl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_5_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_5_IFF_RST,
      O => tx_input_dinl(5)
    );
  DIN_5_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_5_IFF_RST
    );
  tx_input_dinl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_6_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_6_IFF_RST,
      O => tx_input_dinl(6)
    );
  DIN_6_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_6_IFF_RST
    );
  tx_input_dinl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_7_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_7_IFF_RST,
      O => tx_input_dinl(7)
    );
  DIN_7_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_7_IFF_RST
    );
  tx_input_dinl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_8_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_8_IFF_RST,
      O => tx_input_dinl(8)
    );
  DIN_8_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_8_IFF_RST
    );
  tx_input_dinl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_9_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_9_IFF_RST,
      O => tx_input_dinl(9)
    );
  DIN_9_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_9_IFF_RST
    );
  rx_input_GMII_rx_erl_654 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RX_ER_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RX_ER_IFF_RST,
      O => rx_input_GMII_rx_erl
    );
  RX_ER_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RX_ER_IFF_RST
    );
  rx_input_GMII_rx_dvl_655 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RX_DV_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RX_DV_IFF_RST,
      O => rx_input_GMII_rx_dvl
    );
  RX_DV_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RX_DV_IFF_RST
    );
  memcontroller_addr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_10_OD,
      CE => MA_10_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_10_OFF_RST,
      O => memcontroller_ADDREXT(10)
    );
  MA_10_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_10_OFF_RST
    );
  memcontroller_dnout_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_26_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_26_OFF_RST,
      O => memcontroller_dnout(26)
    );
  MD_26_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_26_OFF_RST
    );
  memcontroller_ts_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_26_TFF_RST,
      O => memcontroller_ts(26)
    );
  MD_26_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_26_TFF_RST
    );
  memcontroller_qn_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(19),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_19_IFF_RST,
      O => memcontroller_qn(19)
    );
  MD_19_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_19_IFF_RST
    );
  memcontroller_dnout_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_19_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_19_OFF_RST,
      O => memcontroller_dnout(19)
    );
  MD_19_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_19_OFF_RST
    );
  memcontroller_ts_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_19_TFF_RST,
      O => memcontroller_ts(19)
    );
  MD_19_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_19_TFF_RST
    );
  memcontroller_qn_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(27),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_27_IFF_RST,
      O => memcontroller_qn(27)
    );
  MD_27_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_27_IFF_RST
    );
  memcontroller_qn_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(28),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_28_IFF_RST,
      O => memcontroller_qn(28)
    );
  MD_28_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_28_IFF_RST
    );
  memcontroller_dnout_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_27_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_27_OFF_RST,
      O => memcontroller_dnout(27)
    );
  MD_27_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_27_OFF_RST
    );
  memcontroller_ts_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_27_TFF_RST,
      O => memcontroller_ts(27)
    );
  MD_27_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_27_TFF_RST
    );
  mac_control_rxphyerr_cnt_16_LOGIC_ZERO_656 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_16_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_32_657 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_16_CYINIT,
      SEL => mac_control_rxphyerr_cnt_16_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_16_CYINIT,
      I1 => mac_control_rxphyerr_cnt_16_FROM,
      O => mac_control_rxphyerr_cnt_n0000(16)
    );
  mac_control_rxphyerr_cnt_16_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(16),
      O => mac_control_rxphyerr_cnt_16_FROM
    );
  mac_control_rxphyerr_cnt_16_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(17),
      O => mac_control_rxphyerr_cnt_16_GROM
    );
  mac_control_rxphyerr_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_16_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_33_658 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_rxphyerr_cnt_16_GROM,
      O => mac_control_rxphyerr_cnt_16_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_rxphyerr_cnt_16_GROM,
      O => mac_control_rxphyerr_cnt_n0000(17)
    );
  mac_control_rxphyerr_cnt_16_CYINIT_659 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_rxphyerr_cnt_16_CYINIT
    );
  mac_control_rxphyerr_cnt_18_LOGIC_ZERO_660 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_18_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_34_661 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_18_CYINIT,
      SEL => mac_control_rxphyerr_cnt_18_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_18_CYINIT,
      I1 => mac_control_rxphyerr_cnt_18_FROM,
      O => mac_control_rxphyerr_cnt_n0000(18)
    );
  mac_control_rxphyerr_cnt_18_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(18),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_18_FROM
    );
  mac_control_rxphyerr_cnt_18_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(19),
      O => mac_control_rxphyerr_cnt_18_GROM
    );
  mac_control_rxphyerr_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_18_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_35_662 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_rxphyerr_cnt_18_GROM,
      O => mac_control_rxphyerr_cnt_18_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_rxphyerr_cnt_18_GROM,
      O => mac_control_rxphyerr_cnt_n0000(19)
    );
  mac_control_rxphyerr_cnt_18_CYINIT_663 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_rxphyerr_cnt_18_CYINIT
    );
  mac_control_rxphyerr_cnt_20_LOGIC_ZERO_664 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_20_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_36_665 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_20_CYINIT,
      SEL => mac_control_rxphyerr_cnt_20_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_20_CYINIT,
      I1 => mac_control_rxphyerr_cnt_20_FROM,
      O => mac_control_rxphyerr_cnt_n0000(20)
    );
  mac_control_rxphyerr_cnt_20_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(20),
      O => mac_control_rxphyerr_cnt_20_FROM
    );
  mac_control_rxphyerr_cnt_20_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(21),
      O => mac_control_rxphyerr_cnt_20_GROM
    );
  mac_control_rxphyerr_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_20_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_37_666 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_rxphyerr_cnt_20_GROM,
      O => mac_control_rxphyerr_cnt_20_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_rxphyerr_cnt_20_GROM,
      O => mac_control_rxphyerr_cnt_n0000(21)
    );
  mac_control_rxphyerr_cnt_20_CYINIT_667 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_rxphyerr_cnt_20_CYINIT
    );
  mac_control_rxphyerr_cnt_22_LOGIC_ZERO_668 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_22_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_38_669 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_22_CYINIT,
      SEL => mac_control_rxphyerr_cnt_22_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_22_CYINIT,
      I1 => mac_control_rxphyerr_cnt_22_FROM,
      O => mac_control_rxphyerr_cnt_n0000(22)
    );
  mac_control_rxphyerr_cnt_22_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(22),
      O => mac_control_rxphyerr_cnt_22_FROM
    );
  mac_control_rxphyerr_cnt_22_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(23),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_22_GROM
    );
  mac_control_rxphyerr_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_22_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_39_670 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_rxphyerr_cnt_22_GROM,
      O => mac_control_rxphyerr_cnt_22_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_rxphyerr_cnt_22_GROM,
      O => mac_control_rxphyerr_cnt_n0000(23)
    );
  mac_control_rxphyerr_cnt_22_CYINIT_671 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_rxphyerr_cnt_22_CYINIT
    );
  mac_control_rxphyerr_cnt_24_LOGIC_ZERO_672 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_24_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_40_673 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_24_CYINIT,
      SEL => mac_control_rxphyerr_cnt_24_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_24_CYINIT,
      I1 => mac_control_rxphyerr_cnt_24_FROM,
      O => mac_control_rxphyerr_cnt_n0000(24)
    );
  mac_control_rxphyerr_cnt_24_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(24),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_24_FROM
    );
  mac_control_rxphyerr_cnt_24_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(25),
      O => mac_control_rxphyerr_cnt_24_GROM
    );
  mac_control_rxphyerr_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_24_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_41_674 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_rxphyerr_cnt_24_GROM,
      O => mac_control_rxphyerr_cnt_24_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_rxphyerr_cnt_24_GROM,
      O => mac_control_rxphyerr_cnt_n0000(25)
    );
  mac_control_rxphyerr_cnt_24_CYINIT_675 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_rxphyerr_cnt_24_CYINIT
    );
  mac_control_rxphyerr_cnt_26_LOGIC_ZERO_676 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_26_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_42_677 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_26_CYINIT,
      SEL => mac_control_rxphyerr_cnt_26_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_26_CYINIT,
      I1 => mac_control_rxphyerr_cnt_26_FROM,
      O => mac_control_rxphyerr_cnt_n0000(26)
    );
  mac_control_rxphyerr_cnt_26_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(26),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_26_FROM
    );
  mac_control_rxphyerr_cnt_26_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(27),
      O => mac_control_rxphyerr_cnt_26_GROM
    );
  mac_control_rxphyerr_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_26_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_43_678 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_rxphyerr_cnt_26_GROM,
      O => mac_control_rxphyerr_cnt_26_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_rxphyerr_cnt_26_GROM,
      O => mac_control_rxphyerr_cnt_n0000(27)
    );
  mac_control_rxphyerr_cnt_26_CYINIT_679 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_rxphyerr_cnt_26_CYINIT
    );
  mac_control_rxphyerr_cnt_28_LOGIC_ZERO_680 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_28_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_44_681 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_28_CYINIT,
      SEL => mac_control_rxphyerr_cnt_28_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_28_CYINIT,
      I1 => mac_control_rxphyerr_cnt_28_FROM,
      O => mac_control_rxphyerr_cnt_n0000(28)
    );
  mac_control_rxphyerr_cnt_28_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(28),
      O => mac_control_rxphyerr_cnt_28_FROM
    );
  mac_control_rxphyerr_cnt_28_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(29),
      O => mac_control_rxphyerr_cnt_28_GROM
    );
  mac_control_rxphyerr_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_28_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_45_682 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_rxphyerr_cnt_28_GROM,
      O => mac_control_rxphyerr_cnt_28_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_rxphyerr_cnt_28_GROM,
      O => mac_control_rxphyerr_cnt_n0000(29)
    );
  mac_control_rxphyerr_cnt_28_CYINIT_683 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_rxphyerr_cnt_28_CYINIT
    );
  mac_control_rxphyerr_cnt_30_LOGIC_ZERO_684 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_30_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_46_685 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_30_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_30_CYINIT,
      SEL => mac_control_rxphyerr_cnt_30_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_30_CYINIT,
      I1 => mac_control_rxphyerr_cnt_30_FROM,
      O => mac_control_rxphyerr_cnt_n0000(30)
    );
  mac_control_rxphyerr_cnt_30_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(30),
      O => mac_control_rxphyerr_cnt_30_FROM
    );
  mac_control_rxphyerr_cnt_31_rt_686 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(31),
      O => mac_control_rxphyerr_cnt_31_rt
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_rxphyerr_cnt_31_rt,
      O => mac_control_rxphyerr_cnt_n0000(31)
    );
  mac_control_rxphyerr_cnt_30_CYINIT_687 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_rxphyerr_cnt_30_CYINIT
    );
  mac_control_rxfifowerr_cnt_0_LOGIC_ZERO_688 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_0_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_16_689 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_31,
      IB => mac_control_rxfifowerr_cnt_0_LOGIC_ZERO,
      SEL => mac_control_rxfifowerr_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_31,
      ADR1 => mac_control_rxfifowerr_cnt(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_rxfifowerr_cnt_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_17,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(1),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_0_GROM
    );
  mac_control_rxfifowerr_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_0_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_17_690 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_17,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_rxfifowerr_cnt_0_GROM,
      O => mac_control_rxfifowerr_cnt_0_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_rxfifowerr_cnt_0_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(1)
    );
  mac_control_rxfifowerr_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(3),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(3)
    );
  mac_control_rxfifowerr_cnt_2_LOGIC_ZERO_691 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_2_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_18_692 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_2_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_2_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_2_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_2_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(2)
    );
  mac_control_rxfifowerr_cnt_2_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_2_FROM
    );
  mac_control_rxfifowerr_cnt_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(3),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_2_GROM
    );
  mac_control_rxfifowerr_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_2_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_19_693 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_rxfifowerr_cnt_2_GROM,
      O => mac_control_rxfifowerr_cnt_2_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_rxfifowerr_cnt_2_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(3)
    );
  mac_control_rxfifowerr_cnt_2_CYINIT_694 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_rxfifowerr_cnt_2_CYINIT
    );
  mac_control_rxfifowerr_cnt_4_LOGIC_ZERO_695 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_4_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_20_696 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_4_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_4_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_4_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_4_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(4)
    );
  mac_control_rxfifowerr_cnt_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_4_FROM
    );
  mac_control_rxfifowerr_cnt_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(5),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_4_GROM
    );
  mac_control_rxfifowerr_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_4_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_21_697 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_rxfifowerr_cnt_4_GROM,
      O => mac_control_rxfifowerr_cnt_4_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_rxfifowerr_cnt_4_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(5)
    );
  mac_control_rxfifowerr_cnt_4_CYINIT_698 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_rxfifowerr_cnt_4_CYINIT
    );
  mac_control_rxfifowerr_cnt_6_LOGIC_ZERO_699 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_6_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_22_700 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_6_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_6_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_6_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_6_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(6)
    );
  mac_control_rxfifowerr_cnt_6_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(6),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_6_FROM
    );
  mac_control_rxfifowerr_cnt_6_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(7),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_6_GROM
    );
  mac_control_rxfifowerr_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_6_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_23_701 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_rxfifowerr_cnt_6_GROM,
      O => mac_control_rxfifowerr_cnt_6_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_rxfifowerr_cnt_6_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(7)
    );
  mac_control_rxfifowerr_cnt_6_CYINIT_702 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_rxfifowerr_cnt_6_CYINIT
    );
  mac_control_rxfifowerr_cnt_8_LOGIC_ZERO_703 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_8_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_24_704 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_8_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_8_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_8_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_8_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(8)
    );
  mac_control_rxfifowerr_cnt_8_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_8_FROM
    );
  mac_control_rxfifowerr_cnt_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(9),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_8_GROM
    );
  mac_control_rxfifowerr_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_8_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_25_705 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_rxfifowerr_cnt_8_GROM,
      O => mac_control_rxfifowerr_cnt_8_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_rxfifowerr_cnt_8_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(9)
    );
  mac_control_rxfifowerr_cnt_8_CYINIT_706 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_rxfifowerr_cnt_8_CYINIT
    );
  mac_control_rxfifowerr_cnt_10_LOGIC_ZERO_707 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_10_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_26_708 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_10_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_10_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_10_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_10_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(10)
    );
  mac_control_rxfifowerr_cnt_10_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxfifowerr_cnt(10),
      O => mac_control_rxfifowerr_cnt_10_FROM
    );
  mac_control_rxfifowerr_cnt_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(11),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_10_GROM
    );
  mac_control_rxfifowerr_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_10_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_27_709 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_rxfifowerr_cnt_10_GROM,
      O => mac_control_rxfifowerr_cnt_10_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_rxfifowerr_cnt_10_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(11)
    );
  mac_control_rxfifowerr_cnt_10_CYINIT_710 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_rxfifowerr_cnt_10_CYINIT
    );
  mac_control_rxfifowerr_cnt_12_LOGIC_ZERO_711 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_12_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_28_712 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_12_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_12_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_12_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_12_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(12)
    );
  mac_control_rxfifowerr_cnt_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_12_FROM
    );
  mac_control_rxfifowerr_cnt_12_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(13),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_12_GROM
    );
  mac_control_rxfifowerr_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_12_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_29_713 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_rxfifowerr_cnt_12_GROM,
      O => mac_control_rxfifowerr_cnt_12_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_rxfifowerr_cnt_12_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(13)
    );
  mac_control_rxfifowerr_cnt_12_CYINIT_714 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_rxfifowerr_cnt_12_CYINIT
    );
  mac_control_rxfifowerr_cnt_14_LOGIC_ZERO_715 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_14_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_30_716 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_14_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_14_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_14_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_14_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(14)
    );
  mac_control_rxfifowerr_cnt_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_14_FROM
    );
  mac_control_rxfifowerr_cnt_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(15),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_14_GROM
    );
  mac_control_rxfifowerr_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_14_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_31_717 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_rxfifowerr_cnt_14_GROM,
      O => mac_control_rxfifowerr_cnt_14_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_rxfifowerr_cnt_14_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(15)
    );
  mac_control_rxfifowerr_cnt_14_CYINIT_718 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_rxfifowerr_cnt_14_CYINIT
    );
  mac_control_rxfifowerr_cnt_16_LOGIC_ZERO_719 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_16_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_32_720 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_16_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_16_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_16_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_16_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(16)
    );
  mac_control_rxfifowerr_cnt_16_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_16_FROM
    );
  mac_control_rxfifowerr_cnt_16_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(17),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_16_GROM
    );
  mac_control_rxfifowerr_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_16_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_33_721 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_rxfifowerr_cnt_16_GROM,
      O => mac_control_rxfifowerr_cnt_16_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_rxfifowerr_cnt_16_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(17)
    );
  mac_control_rxfifowerr_cnt_16_CYINIT_722 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_rxfifowerr_cnt_16_CYINIT
    );
  mac_control_rxfifowerr_cnt_18_LOGIC_ZERO_723 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_18_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_34_724 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_18_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_18_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_18_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_18_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(18)
    );
  mac_control_rxfifowerr_cnt_18_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_18_FROM
    );
  mac_control_rxfifowerr_cnt_18_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(19),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_18_GROM
    );
  mac_control_rxfifowerr_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_18_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_35_725 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_rxfifowerr_cnt_18_GROM,
      O => mac_control_rxfifowerr_cnt_18_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_rxfifowerr_cnt_18_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(19)
    );
  mac_control_rxfifowerr_cnt_18_CYINIT_726 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_rxfifowerr_cnt_18_CYINIT
    );
  mac_control_rxfifowerr_cnt_20_LOGIC_ZERO_727 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_20_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_36_728 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_20_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_20_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_20_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_20_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(20)
    );
  mac_control_rxfifowerr_cnt_20_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(20),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_20_FROM
    );
  mac_control_rxfifowerr_cnt_20_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(21),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_20_GROM
    );
  mac_control_rxfifowerr_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_20_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_37_729 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_rxfifowerr_cnt_20_GROM,
      O => mac_control_rxfifowerr_cnt_20_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_rxfifowerr_cnt_20_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(21)
    );
  mac_control_rxfifowerr_cnt_20_CYINIT_730 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_rxfifowerr_cnt_20_CYINIT
    );
  mac_control_rxfifowerr_cnt_22_LOGIC_ZERO_731 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_22_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_38_732 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_22_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_22_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_22_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_22_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(22)
    );
  mac_control_rxfifowerr_cnt_22_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(22),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_22_FROM
    );
  mac_control_rxfifowerr_cnt_22_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(23),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_22_GROM
    );
  mac_control_rxfifowerr_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_22_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_39_733 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_rxfifowerr_cnt_22_GROM,
      O => mac_control_rxfifowerr_cnt_22_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_rxfifowerr_cnt_22_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(23)
    );
  mac_control_rxfifowerr_cnt_22_CYINIT_734 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_rxfifowerr_cnt_22_CYINIT
    );
  mac_control_rxfifowerr_cnt_24_LOGIC_ZERO_735 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_24_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_40_736 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_24_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_24_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_24_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_24_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(24)
    );
  mac_control_rxfifowerr_cnt_24_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(24),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_24_FROM
    );
  mac_control_rxfifowerr_cnt_24_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(25),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_24_GROM
    );
  mac_control_rxfifowerr_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_24_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_41_737 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_rxfifowerr_cnt_24_GROM,
      O => mac_control_rxfifowerr_cnt_24_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_rxfifowerr_cnt_24_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(25)
    );
  mac_control_rxfifowerr_cnt_24_CYINIT_738 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_rxfifowerr_cnt_24_CYINIT
    );
  rx_input_fifo_fifo_BU65 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2807,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N19_FFX_RST,
      O => rx_input_fifo_fifo_N19
    );
  rx_input_fifo_fifo_N19_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N19_FFX_RST
    );
  mac_control_rxfifowerr_cnt_26_LOGIC_ZERO_739 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_26_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_42_740 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_26_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_26_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_26_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_26_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(26)
    );
  mac_control_rxfifowerr_cnt_26_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(26),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_26_FROM
    );
  mac_control_rxfifowerr_cnt_26_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(27),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_26_GROM
    );
  mac_control_rxfifowerr_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_26_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_43_741 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_rxfifowerr_cnt_26_GROM,
      O => mac_control_rxfifowerr_cnt_26_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_rxfifowerr_cnt_26_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(27)
    );
  mac_control_rxfifowerr_cnt_26_CYINIT_742 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_rxfifowerr_cnt_26_CYINIT
    );
  mac_control_rxfifowerr_cnt_28_LOGIC_ZERO_743 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_28_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_44_744 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_28_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_28_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_28_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_28_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(28)
    );
  mac_control_rxfifowerr_cnt_28_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(28),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_28_FROM
    );
  mac_control_rxfifowerr_cnt_28_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(29),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_28_GROM
    );
  mac_control_rxfifowerr_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_28_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_45_745 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_rxfifowerr_cnt_28_GROM,
      O => mac_control_rxfifowerr_cnt_28_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_rxfifowerr_cnt_28_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(29)
    );
  mac_control_rxfifowerr_cnt_28_CYINIT_746 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_rxfifowerr_cnt_28_CYINIT
    );
  mac_control_rxfifowerr_cnt_30_LOGIC_ZERO_747 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_30_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_46_748 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_30_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_30_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_30_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_30_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_30_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(30)
    );
  mac_control_rxfifowerr_cnt_30_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(30),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_30_FROM
    );
  mac_control_rxfifowerr_cnt_31_rt_749 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(31),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_31_rt
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_rxfifowerr_cnt_31_rt,
      O => mac_control_rxfifowerr_cnt_n0000(31)
    );
  mac_control_rxfifowerr_cnt_30_CYINIT_750 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_rxfifowerr_cnt_30_CYINIT
    );
  mac_control_txfifowerr_cnt_0_LOGIC_ZERO_751 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_0_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_16_752 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_1,
      IB => mac_control_txfifowerr_cnt_0_LOGIC_ZERO,
      SEL => mac_control_txfifowerr_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_1,
      ADR1 => mac_control_txfifowerr_cnt(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_txfifowerr_cnt_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_56,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(1),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_0_GROM
    );
  mac_control_txfifowerr_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_0_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_17_753 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_56,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_txfifowerr_cnt_0_GROM,
      O => mac_control_txfifowerr_cnt_0_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_txfifowerr_cnt_0_GROM,
      O => mac_control_txfifowerr_cnt_n0000(1)
    );
  mac_control_txfifowerr_cnt_2_LOGIC_ZERO_754 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_2_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_18_755 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_2_CYINIT,
      SEL => mac_control_txfifowerr_cnt_2_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_2_CYINIT,
      I1 => mac_control_txfifowerr_cnt_2_FROM,
      O => mac_control_txfifowerr_cnt_n0000(2)
    );
  mac_control_txfifowerr_cnt_2_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_2_FROM
    );
  mac_control_txfifowerr_cnt_2_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_2_GROM
    );
  mac_control_txfifowerr_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_2_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_19_756 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_txfifowerr_cnt_2_GROM,
      O => mac_control_txfifowerr_cnt_2_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_txfifowerr_cnt_2_GROM,
      O => mac_control_txfifowerr_cnt_n0000(3)
    );
  mac_control_txfifowerr_cnt_2_CYINIT_757 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_txfifowerr_cnt_2_CYINIT
    );
  mac_control_txfifowerr_cnt_4_LOGIC_ZERO_758 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_4_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_20_759 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_4_CYINIT,
      SEL => mac_control_txfifowerr_cnt_4_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_4_CYINIT,
      I1 => mac_control_txfifowerr_cnt_4_FROM,
      O => mac_control_txfifowerr_cnt_n0000(4)
    );
  mac_control_txfifowerr_cnt_4_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_4_FROM
    );
  mac_control_txfifowerr_cnt_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(5),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_4_GROM
    );
  mac_control_txfifowerr_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_4_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_21_760 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_txfifowerr_cnt_4_GROM,
      O => mac_control_txfifowerr_cnt_4_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_txfifowerr_cnt_4_GROM,
      O => mac_control_txfifowerr_cnt_n0000(5)
    );
  mac_control_txfifowerr_cnt_4_CYINIT_761 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_txfifowerr_cnt_4_CYINIT
    );
  mac_control_txfifowerr_cnt_6_LOGIC_ZERO_762 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_6_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_22_763 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_6_CYINIT,
      SEL => mac_control_txfifowerr_cnt_6_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_6_CYINIT,
      I1 => mac_control_txfifowerr_cnt_6_FROM,
      O => mac_control_txfifowerr_cnt_n0000(6)
    );
  mac_control_txfifowerr_cnt_6_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txfifowerr_cnt(6),
      O => mac_control_txfifowerr_cnt_6_FROM
    );
  mac_control_txfifowerr_cnt_6_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(7),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_6_GROM
    );
  mac_control_txfifowerr_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_6_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_23_764 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_txfifowerr_cnt_6_GROM,
      O => mac_control_txfifowerr_cnt_6_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_txfifowerr_cnt_6_GROM,
      O => mac_control_txfifowerr_cnt_n0000(7)
    );
  mac_control_txfifowerr_cnt_6_CYINIT_765 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_txfifowerr_cnt_6_CYINIT
    );
  mac_control_txfifowerr_cnt_8_LOGIC_ZERO_766 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_8_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_24_767 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_8_CYINIT,
      SEL => mac_control_txfifowerr_cnt_8_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_8_CYINIT,
      I1 => mac_control_txfifowerr_cnt_8_FROM,
      O => mac_control_txfifowerr_cnt_n0000(8)
    );
  mac_control_txfifowerr_cnt_8_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_8_FROM
    );
  mac_control_txfifowerr_cnt_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(9),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_8_GROM
    );
  mac_control_txfifowerr_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_8_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_25_768 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_txfifowerr_cnt_8_GROM,
      O => mac_control_txfifowerr_cnt_8_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_txfifowerr_cnt_8_GROM,
      O => mac_control_txfifowerr_cnt_n0000(9)
    );
  mac_control_txfifowerr_cnt_8_CYINIT_769 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_txfifowerr_cnt_8_CYINIT
    );
  mac_control_txfifowerr_cnt_10_LOGIC_ZERO_770 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_10_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_26_771 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_10_CYINIT,
      SEL => mac_control_txfifowerr_cnt_10_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_10_CYINIT,
      I1 => mac_control_txfifowerr_cnt_10_FROM,
      O => mac_control_txfifowerr_cnt_n0000(10)
    );
  mac_control_txfifowerr_cnt_10_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(10),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_10_FROM
    );
  mac_control_txfifowerr_cnt_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(11),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_10_GROM
    );
  mac_control_txfifowerr_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_10_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_27_772 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_txfifowerr_cnt_10_GROM,
      O => mac_control_txfifowerr_cnt_10_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_txfifowerr_cnt_10_GROM,
      O => mac_control_txfifowerr_cnt_n0000(11)
    );
  mac_control_txfifowerr_cnt_10_CYINIT_773 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_txfifowerr_cnt_10_CYINIT
    );
  mac_control_txfifowerr_cnt_12_LOGIC_ZERO_774 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_12_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_28_775 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_12_CYINIT,
      SEL => mac_control_txfifowerr_cnt_12_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_12_CYINIT,
      I1 => mac_control_txfifowerr_cnt_12_FROM,
      O => mac_control_txfifowerr_cnt_n0000(12)
    );
  mac_control_txfifowerr_cnt_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_12_FROM
    );
  mac_control_txfifowerr_cnt_12_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_12_GROM
    );
  mac_control_txfifowerr_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_12_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_29_776 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_txfifowerr_cnt_12_GROM,
      O => mac_control_txfifowerr_cnt_12_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_txfifowerr_cnt_12_GROM,
      O => mac_control_txfifowerr_cnt_n0000(13)
    );
  mac_control_txfifowerr_cnt_12_CYINIT_777 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_txfifowerr_cnt_12_CYINIT
    );
  mac_control_txfifowerr_cnt_14_LOGIC_ZERO_778 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_14_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_30_779 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_14_CYINIT,
      SEL => mac_control_txfifowerr_cnt_14_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_14_CYINIT,
      I1 => mac_control_txfifowerr_cnt_14_FROM,
      O => mac_control_txfifowerr_cnt_n0000(14)
    );
  mac_control_txfifowerr_cnt_14_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(14),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_14_FROM
    );
  mac_control_txfifowerr_cnt_14_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(15),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_14_GROM
    );
  mac_control_txfifowerr_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_14_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_31_780 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_txfifowerr_cnt_14_GROM,
      O => mac_control_txfifowerr_cnt_14_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_txfifowerr_cnt_14_GROM,
      O => mac_control_txfifowerr_cnt_n0000(15)
    );
  mac_control_txfifowerr_cnt_14_CYINIT_781 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_txfifowerr_cnt_14_CYINIT
    );
  mac_control_txfifowerr_cnt_16_LOGIC_ZERO_782 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_16_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_32_783 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_16_CYINIT,
      SEL => mac_control_txfifowerr_cnt_16_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_16_CYINIT,
      I1 => mac_control_txfifowerr_cnt_16_FROM,
      O => mac_control_txfifowerr_cnt_n0000(16)
    );
  mac_control_txfifowerr_cnt_16_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_16_FROM
    );
  mac_control_txfifowerr_cnt_16_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(17),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_16_GROM
    );
  mac_control_txfifowerr_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_16_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_33_784 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_txfifowerr_cnt_16_GROM,
      O => mac_control_txfifowerr_cnt_16_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_txfifowerr_cnt_16_GROM,
      O => mac_control_txfifowerr_cnt_n0000(17)
    );
  mac_control_txfifowerr_cnt_16_CYINIT_785 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_txfifowerr_cnt_16_CYINIT
    );
  rx_input_fifo_fifo_BU122 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3280,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2406_FFY_RST,
      O => rx_input_fifo_fifo_N2405
    );
  rx_input_fifo_fifo_N2406_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2406_FFY_RST
    );
  mac_control_txfifowerr_cnt_18_LOGIC_ZERO_786 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_18_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_34_787 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_18_CYINIT,
      SEL => mac_control_txfifowerr_cnt_18_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_18_CYINIT,
      I1 => mac_control_txfifowerr_cnt_18_FROM,
      O => mac_control_txfifowerr_cnt_n0000(18)
    );
  mac_control_txfifowerr_cnt_18_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_18_FROM
    );
  mac_control_txfifowerr_cnt_18_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(19),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_18_GROM
    );
  mac_control_txfifowerr_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_18_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_35_788 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_txfifowerr_cnt_18_GROM,
      O => mac_control_txfifowerr_cnt_18_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_txfifowerr_cnt_18_GROM,
      O => mac_control_txfifowerr_cnt_n0000(19)
    );
  mac_control_txfifowerr_cnt_18_CYINIT_789 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_txfifowerr_cnt_18_CYINIT
    );
  mac_control_txfifowerr_cnt_20_LOGIC_ZERO_790 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_20_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_36_791 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_20_CYINIT,
      SEL => mac_control_txfifowerr_cnt_20_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_20_CYINIT,
      I1 => mac_control_txfifowerr_cnt_20_FROM,
      O => mac_control_txfifowerr_cnt_n0000(20)
    );
  mac_control_txfifowerr_cnt_20_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(20),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_20_FROM
    );
  mac_control_txfifowerr_cnt_20_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(21),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_20_GROM
    );
  mac_control_txfifowerr_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_20_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_37_792 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_txfifowerr_cnt_20_GROM,
      O => mac_control_txfifowerr_cnt_20_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_txfifowerr_cnt_20_GROM,
      O => mac_control_txfifowerr_cnt_n0000(21)
    );
  mac_control_txfifowerr_cnt_20_CYINIT_793 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_txfifowerr_cnt_20_CYINIT
    );
  mac_control_txfifowerr_cnt_22_LOGIC_ZERO_794 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_22_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_38_795 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_22_CYINIT,
      SEL => mac_control_txfifowerr_cnt_22_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_22_CYINIT,
      I1 => mac_control_txfifowerr_cnt_22_FROM,
      O => mac_control_txfifowerr_cnt_n0000(22)
    );
  mac_control_txfifowerr_cnt_22_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(22),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_22_FROM
    );
  mac_control_txfifowerr_cnt_22_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txfifowerr_cnt(23),
      O => mac_control_txfifowerr_cnt_22_GROM
    );
  mac_control_txfifowerr_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_22_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_39_796 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_txfifowerr_cnt_22_GROM,
      O => mac_control_txfifowerr_cnt_22_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_txfifowerr_cnt_22_GROM,
      O => mac_control_txfifowerr_cnt_n0000(23)
    );
  mac_control_txfifowerr_cnt_22_CYINIT_797 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_txfifowerr_cnt_22_CYINIT
    );
  mac_control_txfifowerr_cnt_24_LOGIC_ZERO_798 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_24_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_40_799 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_24_CYINIT,
      SEL => mac_control_txfifowerr_cnt_24_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_24_CYINIT,
      I1 => mac_control_txfifowerr_cnt_24_FROM,
      O => mac_control_txfifowerr_cnt_n0000(24)
    );
  mac_control_txfifowerr_cnt_24_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(24),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_24_FROM
    );
  mac_control_txfifowerr_cnt_24_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(25),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_24_GROM
    );
  mac_control_txfifowerr_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_24_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_41_800 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_txfifowerr_cnt_24_GROM,
      O => mac_control_txfifowerr_cnt_24_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_txfifowerr_cnt_24_GROM,
      O => mac_control_txfifowerr_cnt_n0000(25)
    );
  mac_control_txfifowerr_cnt_24_CYINIT_801 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_txfifowerr_cnt_24_CYINIT
    );
  mac_control_txfifowerr_cnt_26_LOGIC_ZERO_802 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_26_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_42_803 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_26_CYINIT,
      SEL => mac_control_txfifowerr_cnt_26_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_26_CYINIT,
      I1 => mac_control_txfifowerr_cnt_26_FROM,
      O => mac_control_txfifowerr_cnt_n0000(26)
    );
  mac_control_txfifowerr_cnt_26_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(26),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_26_FROM
    );
  mac_control_txfifowerr_cnt_26_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(27),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_26_GROM
    );
  mac_control_txfifowerr_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_26_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_43_804 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_txfifowerr_cnt_26_GROM,
      O => mac_control_txfifowerr_cnt_26_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_txfifowerr_cnt_26_GROM,
      O => mac_control_txfifowerr_cnt_n0000(27)
    );
  mac_control_txfifowerr_cnt_26_CYINIT_805 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_txfifowerr_cnt_26_CYINIT
    );
  mac_control_txfifowerr_cnt_28_LOGIC_ZERO_806 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_28_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_44_807 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_28_CYINIT,
      SEL => mac_control_txfifowerr_cnt_28_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_28_CYINIT,
      I1 => mac_control_txfifowerr_cnt_28_FROM,
      O => mac_control_txfifowerr_cnt_n0000(28)
    );
  mac_control_txfifowerr_cnt_28_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(28),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_28_FROM
    );
  mac_control_txfifowerr_cnt_28_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(29),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_28_GROM
    );
  mac_control_txfifowerr_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_28_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_45_808 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_txfifowerr_cnt_28_GROM,
      O => mac_control_txfifowerr_cnt_28_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_txfifowerr_cnt_28_GROM,
      O => mac_control_txfifowerr_cnt_n0000(29)
    );
  mac_control_txfifowerr_cnt_28_CYINIT_809 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_txfifowerr_cnt_28_CYINIT
    );
  mac_control_txfifowerr_cnt_30_LOGIC_ZERO_810 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_30_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_46_811 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_30_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_30_CYINIT,
      SEL => mac_control_txfifowerr_cnt_30_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_30_CYINIT,
      I1 => mac_control_txfifowerr_cnt_30_FROM,
      O => mac_control_txfifowerr_cnt_n0000(30)
    );
  mac_control_txfifowerr_cnt_30_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(30),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_30_FROM
    );
  mac_control_txfifowerr_cnt_31_rt_812 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(31),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_31_rt
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_txfifowerr_cnt_31_rt,
      O => mac_control_txfifowerr_cnt_n0000(31)
    );
  mac_control_txfifowerr_cnt_30_CYINIT_813 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_txfifowerr_cnt_30_CYINIT
    );
  rx_input_fifo_fifo_BU59 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2806,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N21_FFY_RST,
      O => rx_input_fifo_fifo_N20
    );
  rx_input_fifo_fifo_N21_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N21_FFY_RST
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ONE_814 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ZERO_815 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_177_816 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(25),
      ADR1 => rx_input_memio_addrchk_datal(24),
      ADR2 => rx_input_memio_addrchk_macaddrl(25),
      ADR3 => rx_input_memio_addrchk_macaddrl(24),
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(27),
      ADR1 => rx_input_memio_addrchk_datal(26),
      ADR2 => rx_input_memio_addrchk_macaddrl(27),
      ADR3 => rx_input_memio_addrchk_macaddrl(26),
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_817 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_2_LOGIC_ZERO_818 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_2_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_179_819 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_2_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_2_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(28),
      ADR1 => rx_input_memio_addrchk_datal(29),
      ADR2 => rx_input_memio_addrchk_macaddrl(29),
      ADR3 => rx_input_memio_addrchk_macaddrl(28),
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(30),
      ADR1 => rx_input_memio_addrchk_datal(31),
      ADR2 => rx_input_memio_addrchk_macaddrl(31),
      ADR3 => rx_input_memio_addrchk_macaddrl(30),
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_2_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_2_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(2)
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_2_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_2_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_2_CYINIT_820 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_2_CYINIT
    );
  rx_output_bp_0_LOGIC_ONE_821 : X_ONE
    port map (
      O => rx_output_bp_0_LOGIC_ONE
    );
  rx_output_Madd_lbp_inst_cy_86_822 : X_MUX2
    port map (
      IA => rx_output_lenr(2),
      IB => rx_output_bp_0_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_79,
      O => rx_output_Madd_lbp_inst_cy_86
    );
  rx_output_Madd_lbp_inst_sum_79 : X_XOR2
    port map (
      I0 => rx_output_bp_0_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_79,
      O => rx_output_lbp(0)
    );
  rx_output_Madd_lbp_inst_lut2_791 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_lenr(2),
      ADR1 => VCC,
      ADR2 => rx_output_bp(0),
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_79
    );
  rx_output_Madd_lbp_inst_lut2_801 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(1),
      O => rx_output_Madd_lbp_inst_lut2_80
    );
  rx_output_bp_0_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_0_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_87
    );
  rx_output_Madd_lbp_inst_cy_87_823 : X_MUX2
    port map (
      IA => rx_output_lenr(3),
      IB => rx_output_Madd_lbp_inst_cy_86,
      SEL => rx_output_Madd_lbp_inst_lut2_80,
      O => rx_output_bp_0_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_80 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_86,
      I1 => rx_output_Madd_lbp_inst_lut2_80,
      O => rx_output_lbp(1)
    );
  rx_output_bp_0_CYINIT_824 : X_BUF
    port map (
      I => rx_output_bp_0_LOGIC_ONE,
      O => rx_output_bp_0_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_88_825 : X_MUX2
    port map (
      IA => rx_output_lenr(4),
      IB => rx_output_bp_2_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_81,
      O => rx_output_Madd_lbp_inst_cy_88
    );
  rx_output_Madd_lbp_inst_sum_81 : X_XOR2
    port map (
      I0 => rx_output_bp_2_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_81,
      O => rx_output_lbp(2)
    );
  rx_output_Madd_lbp_inst_lut2_811 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_lenr(4),
      ADR1 => VCC,
      ADR2 => rx_output_bp(2),
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_81
    );
  rx_output_Madd_lbp_inst_lut2_821 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(3),
      O => rx_output_Madd_lbp_inst_lut2_82
    );
  rx_output_bp_2_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_2_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_89
    );
  rx_output_Madd_lbp_inst_cy_89_826 : X_MUX2
    port map (
      IA => rx_output_lenr(5),
      IB => rx_output_Madd_lbp_inst_cy_88,
      SEL => rx_output_Madd_lbp_inst_lut2_82,
      O => rx_output_bp_2_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_82 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_88,
      I1 => rx_output_Madd_lbp_inst_lut2_82,
      O => rx_output_lbp(3)
    );
  rx_output_bp_2_CYINIT_827 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_87,
      O => rx_output_bp_2_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_90_828 : X_MUX2
    port map (
      IA => rx_output_lenr(6),
      IB => rx_output_bp_4_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_83,
      O => rx_output_Madd_lbp_inst_cy_90
    );
  rx_output_Madd_lbp_inst_sum_83 : X_XOR2
    port map (
      I0 => rx_output_bp_4_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_83,
      O => rx_output_lbp(4)
    );
  rx_output_Madd_lbp_inst_lut2_831 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_lenr(6),
      ADR1 => VCC,
      ADR2 => rx_output_bp(4),
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_83
    );
  rx_output_Madd_lbp_inst_lut2_841 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(7),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(5),
      O => rx_output_Madd_lbp_inst_lut2_84
    );
  rx_output_bp_4_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_4_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_91
    );
  rx_output_Madd_lbp_inst_cy_91_829 : X_MUX2
    port map (
      IA => rx_output_lenr(7),
      IB => rx_output_Madd_lbp_inst_cy_90,
      SEL => rx_output_Madd_lbp_inst_lut2_84,
      O => rx_output_bp_4_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_84 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_90,
      I1 => rx_output_Madd_lbp_inst_lut2_84,
      O => rx_output_lbp(5)
    );
  rx_output_bp_4_CYINIT_830 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_89,
      O => rx_output_bp_4_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_92_831 : X_MUX2
    port map (
      IA => rx_output_lenr(8),
      IB => rx_output_bp_6_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_85,
      O => rx_output_Madd_lbp_inst_cy_92
    );
  rx_output_Madd_lbp_inst_sum_85 : X_XOR2
    port map (
      I0 => rx_output_bp_6_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_85,
      O => rx_output_lbp(6)
    );
  rx_output_Madd_lbp_inst_lut2_851 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_lenr(8),
      ADR1 => VCC,
      ADR2 => rx_output_bp(6),
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_85
    );
  rx_output_Madd_lbp_inst_lut2_861 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(7),
      O => rx_output_Madd_lbp_inst_lut2_86
    );
  rx_output_bp_6_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_6_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_93
    );
  rx_output_Madd_lbp_inst_cy_93_832 : X_MUX2
    port map (
      IA => rx_output_lenr(9),
      IB => rx_output_Madd_lbp_inst_cy_92,
      SEL => rx_output_Madd_lbp_inst_lut2_86,
      O => rx_output_bp_6_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_86 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_92,
      I1 => rx_output_Madd_lbp_inst_lut2_86,
      O => rx_output_lbp(7)
    );
  rx_output_bp_6_CYINIT_833 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_91,
      O => rx_output_bp_6_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_94_834 : X_MUX2
    port map (
      IA => rx_output_lenr(10),
      IB => rx_output_bp_8_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_87,
      O => rx_output_Madd_lbp_inst_cy_94
    );
  rx_output_Madd_lbp_inst_sum_87 : X_XOR2
    port map (
      I0 => rx_output_bp_8_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_87,
      O => rx_output_lbp(8)
    );
  rx_output_Madd_lbp_inst_lut2_871 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_lenr(10),
      ADR1 => rx_output_bp(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_87
    );
  rx_output_Madd_lbp_inst_lut2_881 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_lenr(11),
      ADR1 => rx_output_bp(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_88
    );
  rx_output_bp_8_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_8_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_95
    );
  rx_output_Madd_lbp_inst_cy_95_835 : X_MUX2
    port map (
      IA => rx_output_lenr(11),
      IB => rx_output_Madd_lbp_inst_cy_94,
      SEL => rx_output_Madd_lbp_inst_lut2_88,
      O => rx_output_bp_8_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_88 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_94,
      I1 => rx_output_Madd_lbp_inst_lut2_88,
      O => rx_output_lbp(9)
    );
  rx_output_bp_8_CYINIT_836 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_93,
      O => rx_output_bp_8_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_96_837 : X_MUX2
    port map (
      IA => rx_output_lenr(12),
      IB => rx_output_bp_10_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_89,
      O => rx_output_Madd_lbp_inst_cy_96
    );
  rx_output_Madd_lbp_inst_sum_89 : X_XOR2
    port map (
      I0 => rx_output_bp_10_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_89,
      O => rx_output_lbp(10)
    );
  rx_output_Madd_lbp_inst_lut2_891 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_lenr(12),
      ADR1 => VCC,
      ADR2 => rx_output_bp(10),
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_89
    );
  rx_output_Madd_lbp_inst_lut2_901 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(11),
      O => rx_output_Madd_lbp_inst_lut2_90
    );
  rx_output_bp_10_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_10_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_97
    );
  rx_output_Madd_lbp_inst_cy_97_838 : X_MUX2
    port map (
      IA => rx_output_lenr(13),
      IB => rx_output_Madd_lbp_inst_cy_96,
      SEL => rx_output_Madd_lbp_inst_lut2_90,
      O => rx_output_bp_10_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_90 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_96,
      I1 => rx_output_Madd_lbp_inst_lut2_90,
      O => rx_output_lbp(11)
    );
  rx_output_bp_10_CYINIT_839 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_95,
      O => rx_output_bp_10_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_98_840 : X_MUX2
    port map (
      IA => rx_output_lenr(14),
      IB => rx_output_bp_12_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_91,
      O => rx_output_Madd_lbp_inst_cy_98
    );
  rx_output_Madd_lbp_inst_sum_91 : X_XOR2
    port map (
      I0 => rx_output_bp_12_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_91,
      O => rx_output_lbp(12)
    );
  rx_output_Madd_lbp_inst_lut2_911 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_lenr(14),
      ADR1 => rx_output_bp(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_91
    );
  rx_output_Madd_lbp_inst_lut2_921 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(15),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(13),
      O => rx_output_Madd_lbp_inst_lut2_92
    );
  rx_output_bp_12_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_12_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_99
    );
  rx_output_Madd_lbp_inst_cy_99_841 : X_MUX2
    port map (
      IA => rx_output_lenr(15),
      IB => rx_output_Madd_lbp_inst_cy_98,
      SEL => rx_output_Madd_lbp_inst_lut2_92,
      O => rx_output_bp_12_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_92 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_98,
      I1 => rx_output_Madd_lbp_inst_lut2_92,
      O => rx_output_lbp(13)
    );
  rx_output_bp_12_CYINIT_842 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_97,
      O => rx_output_bp_12_CYINIT
    );
  rx_output_bp_14_LOGIC_ZERO_843 : X_ZERO
    port map (
      O => rx_output_bp_14_LOGIC_ZERO
    );
  rx_output_Madd_lbp_inst_cy_100_844 : X_MUX2
    port map (
      IA => rx_output_bp_14_LOGIC_ZERO,
      IB => rx_output_bp_14_CYINIT,
      SEL => rx_output_bp_14_FROM,
      O => rx_output_Madd_lbp_inst_cy_100
    );
  rx_output_Madd_lbp_inst_sum_93 : X_XOR2
    port map (
      I0 => rx_output_bp_14_CYINIT,
      I1 => rx_output_bp_14_FROM,
      O => rx_output_lbp(14)
    );
  rx_output_bp_14_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_bp(14),
      ADR3 => VCC,
      O => rx_output_bp_14_FROM
    );
  rx_output_bp_15_rt_845 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(15),
      O => rx_output_bp_15_rt
    );
  rx_output_Madd_lbp_inst_sum_94 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_100,
      I1 => rx_output_bp_15_rt,
      O => rx_output_lbp(15)
    );
  rx_output_bp_14_CYINIT_846 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_99,
      O => rx_output_bp_14_CYINIT
    );
  tx_output_bcnt_38_LOGIC_ONE_847 : X_ONE
    port map (
      O => tx_output_bcnt_38_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_204_848 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_46,
      IB => tx_output_bcnt_38_LOGIC_ONE,
      SEL => tx_output_cs_FFd12_rt,
      O => tx_output_bcnt_inst_cy_204
    );
  tx_output_cs_FFd12_rt_849 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_46,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_output_cs_FFd12_rt
    );
  tx_output_bcnt_inst_lut3_401 : X_LUT4
    generic map(
      INIT => X"0F33"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_8,
      ADR1 => tx_output_bcnt_38,
      ADR2 => q2(0),
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_40
    );
  tx_output_bcnt_38_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_38_CYMUXG,
      O => tx_output_bcnt_inst_cy_205
    );
  tx_output_bcnt_inst_cy_205_850 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_8,
      IB => tx_output_bcnt_inst_cy_204,
      SEL => tx_output_bcnt_inst_lut3_40,
      O => tx_output_bcnt_38_CYMUXG
    );
  tx_output_bcnt_inst_sum_171_851 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_204,
      I1 => tx_output_bcnt_inst_lut3_40,
      O => tx_output_bcnt_inst_sum_171
    );
  tx_output_bcnt_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_39_FFY_RST
    );
  tx_output_bcnt_40_852 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_173,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_39_FFY_RST,
      O => tx_output_bcnt_40
    );
  tx_output_bcnt_39_LOGIC_ONE_853 : X_ONE
    port map (
      O => tx_output_bcnt_39_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_206_854 : X_MUX2
    port map (
      IA => tx_output_bcnt_39_LOGIC_ONE,
      IB => tx_output_bcnt_39_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_41,
      O => tx_output_bcnt_inst_cy_206
    );
  tx_output_bcnt_inst_sum_172_855 : X_XOR2
    port map (
      I0 => tx_output_bcnt_39_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_41,
      O => tx_output_bcnt_inst_sum_172
    );
  tx_output_bcnt_inst_lut3_411 : X_LUT4
    generic map(
      INIT => X"3355"
    )
    port map (
      ADR0 => tx_output_bcnt_39,
      ADR1 => q2(1),
      ADR2 => VCC,
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_41
    );
  tx_output_bcnt_inst_lut3_421 : X_LUT4
    generic map(
      INIT => X"3355"
    )
    port map (
      ADR0 => tx_output_bcnt_40,
      ADR1 => q2(2),
      ADR2 => VCC,
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_42
    );
  tx_output_bcnt_39_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_39_CYMUXG,
      O => tx_output_bcnt_inst_cy_207
    );
  tx_output_bcnt_inst_cy_207_856 : X_MUX2
    port map (
      IA => tx_output_bcnt_39_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_206,
      SEL => tx_output_bcnt_inst_lut3_42,
      O => tx_output_bcnt_39_CYMUXG
    );
  tx_output_bcnt_inst_sum_173_857 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_206,
      I1 => tx_output_bcnt_inst_lut3_42,
      O => tx_output_bcnt_inst_sum_173
    );
  tx_output_bcnt_39_CYINIT_858 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_205,
      O => tx_output_bcnt_39_CYINIT
    );
  tx_output_bcnt_41_LOGIC_ONE_859 : X_ONE
    port map (
      O => tx_output_bcnt_41_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_208_860 : X_MUX2
    port map (
      IA => tx_output_bcnt_41_LOGIC_ONE,
      IB => tx_output_bcnt_41_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_43,
      O => tx_output_bcnt_inst_cy_208
    );
  tx_output_bcnt_inst_sum_174_861 : X_XOR2
    port map (
      I0 => tx_output_bcnt_41_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_43,
      O => tx_output_bcnt_inst_sum_174
    );
  tx_output_bcnt_inst_lut3_431 : X_LUT4
    generic map(
      INIT => X"0F33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_bcnt_41,
      ADR2 => q2(3),
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_43
    );
  tx_output_bcnt_inst_lut3_441 : X_LUT4
    generic map(
      INIT => X"03CF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_bcnt_42,
      ADR3 => q2(4),
      O => tx_output_bcnt_inst_lut3_44
    );
  tx_output_bcnt_41_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_41_CYMUXG,
      O => tx_output_bcnt_inst_cy_209
    );
  tx_output_bcnt_inst_cy_209_862 : X_MUX2
    port map (
      IA => tx_output_bcnt_41_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_208,
      SEL => tx_output_bcnt_inst_lut3_44,
      O => tx_output_bcnt_41_CYMUXG
    );
  tx_output_bcnt_inst_sum_175_863 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_208,
      I1 => tx_output_bcnt_inst_lut3_44,
      O => tx_output_bcnt_inst_sum_175
    );
  tx_output_bcnt_41_CYINIT_864 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_207,
      O => tx_output_bcnt_41_CYINIT
    );
  tx_output_bcnt_43_LOGIC_ONE_865 : X_ONE
    port map (
      O => tx_output_bcnt_43_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_210_866 : X_MUX2
    port map (
      IA => tx_output_bcnt_43_LOGIC_ONE,
      IB => tx_output_bcnt_43_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_45,
      O => tx_output_bcnt_inst_cy_210
    );
  tx_output_bcnt_inst_sum_176_867 : X_XOR2
    port map (
      I0 => tx_output_bcnt_43_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_45,
      O => tx_output_bcnt_inst_sum_176
    );
  tx_output_bcnt_inst_lut3_451 : X_LUT4
    generic map(
      INIT => X"4477"
    )
    port map (
      ADR0 => q2(5),
      ADR1 => tx_output_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_output_bcnt_43,
      O => tx_output_bcnt_inst_lut3_45
    );
  tx_output_bcnt_inst_lut3_461 : X_LUT4
    generic map(
      INIT => X"05F5"
    )
    port map (
      ADR0 => tx_output_bcnt_44,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd12,
      ADR3 => q2(6),
      O => tx_output_bcnt_inst_lut3_46
    );
  tx_output_bcnt_43_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_43_CYMUXG,
      O => tx_output_bcnt_inst_cy_211
    );
  tx_output_bcnt_inst_cy_211_868 : X_MUX2
    port map (
      IA => tx_output_bcnt_43_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_210,
      SEL => tx_output_bcnt_inst_lut3_46,
      O => tx_output_bcnt_43_CYMUXG
    );
  tx_output_bcnt_inst_sum_177_869 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_210,
      I1 => tx_output_bcnt_inst_lut3_46,
      O => tx_output_bcnt_inst_sum_177
    );
  tx_output_bcnt_43_CYINIT_870 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_209,
      O => tx_output_bcnt_43_CYINIT
    );
  tx_output_bcnt_45_LOGIC_ONE_871 : X_ONE
    port map (
      O => tx_output_bcnt_45_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_212_872 : X_MUX2
    port map (
      IA => tx_output_bcnt_45_LOGIC_ONE,
      IB => tx_output_bcnt_45_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_47,
      O => tx_output_bcnt_inst_cy_212
    );
  tx_output_bcnt_inst_sum_178_873 : X_XOR2
    port map (
      I0 => tx_output_bcnt_45_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_47,
      O => tx_output_bcnt_inst_sum_178
    );
  tx_output_bcnt_inst_lut3_471 : X_LUT4
    generic map(
      INIT => X"4477"
    )
    port map (
      ADR0 => q2(7),
      ADR1 => tx_output_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_output_bcnt_45,
      O => tx_output_bcnt_inst_lut3_47
    );
  tx_output_bcnt_inst_lut3_481 : X_LUT4
    generic map(
      INIT => X"0C3F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => q2(8),
      ADR3 => tx_output_bcnt_46,
      O => tx_output_bcnt_inst_lut3_48
    );
  tx_output_bcnt_45_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_45_CYMUXG,
      O => tx_output_bcnt_inst_cy_213
    );
  tx_output_bcnt_inst_cy_213_874 : X_MUX2
    port map (
      IA => tx_output_bcnt_45_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_212,
      SEL => tx_output_bcnt_inst_lut3_48,
      O => tx_output_bcnt_45_CYMUXG
    );
  tx_output_bcnt_inst_sum_179_875 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_212,
      I1 => tx_output_bcnt_inst_lut3_48,
      O => tx_output_bcnt_inst_sum_179
    );
  tx_output_bcnt_45_CYINIT_876 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_211,
      O => tx_output_bcnt_45_CYINIT
    );
  tx_output_bcnt_47_LOGIC_ONE_877 : X_ONE
    port map (
      O => tx_output_bcnt_47_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_214_878 : X_MUX2
    port map (
      IA => tx_output_bcnt_47_LOGIC_ONE,
      IB => tx_output_bcnt_47_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_49,
      O => tx_output_bcnt_inst_cy_214
    );
  tx_output_bcnt_inst_sum_180_879 : X_XOR2
    port map (
      I0 => tx_output_bcnt_47_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_49,
      O => tx_output_bcnt_inst_sum_180
    );
  tx_output_bcnt_inst_lut3_491 : X_LUT4
    generic map(
      INIT => X"03CF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_bcnt_47,
      ADR3 => q2(9),
      O => tx_output_bcnt_inst_lut3_49
    );
  tx_output_bcnt_inst_lut3_501 : X_LUT4
    generic map(
      INIT => X"4747"
    )
    port map (
      ADR0 => q2(10),
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_bcnt_48,
      ADR3 => VCC,
      O => tx_output_bcnt_inst_lut3_50
    );
  tx_output_bcnt_47_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_47_CYMUXG,
      O => tx_output_bcnt_inst_cy_215
    );
  tx_output_bcnt_inst_cy_215_880 : X_MUX2
    port map (
      IA => tx_output_bcnt_47_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_214,
      SEL => tx_output_bcnt_inst_lut3_50,
      O => tx_output_bcnt_47_CYMUXG
    );
  tx_output_bcnt_inst_sum_181_881 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_214,
      I1 => tx_output_bcnt_inst_lut3_50,
      O => tx_output_bcnt_inst_sum_181
    );
  tx_output_bcnt_47_CYINIT_882 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_213,
      O => tx_output_bcnt_47_CYINIT
    );
  tx_output_bcnt_49_LOGIC_ONE_883 : X_ONE
    port map (
      O => tx_output_bcnt_49_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_216_884 : X_MUX2
    port map (
      IA => tx_output_bcnt_49_LOGIC_ONE,
      IB => tx_output_bcnt_49_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_51,
      O => tx_output_bcnt_inst_cy_216
    );
  tx_output_bcnt_inst_sum_182_885 : X_XOR2
    port map (
      I0 => tx_output_bcnt_49_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_51,
      O => tx_output_bcnt_inst_sum_182
    );
  tx_output_bcnt_inst_lut3_511 : X_LUT4
    generic map(
      INIT => X"5353"
    )
    port map (
      ADR0 => q2(11),
      ADR1 => tx_output_bcnt_49,
      ADR2 => tx_output_cs_FFd12,
      ADR3 => VCC,
      O => tx_output_bcnt_inst_lut3_51
    );
  tx_output_bcnt_inst_lut3_521 : X_LUT4
    generic map(
      INIT => X"1D1D"
    )
    port map (
      ADR0 => tx_output_bcnt_50,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => q2(12),
      ADR3 => VCC,
      O => tx_output_bcnt_inst_lut3_52
    );
  tx_output_bcnt_49_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_49_CYMUXG,
      O => tx_output_bcnt_inst_cy_217
    );
  tx_output_bcnt_inst_cy_217_886 : X_MUX2
    port map (
      IA => tx_output_bcnt_49_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_216,
      SEL => tx_output_bcnt_inst_lut3_52,
      O => tx_output_bcnt_49_CYMUXG
    );
  tx_output_bcnt_inst_sum_183_887 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_216,
      I1 => tx_output_bcnt_inst_lut3_52,
      O => tx_output_bcnt_inst_sum_183
    );
  tx_output_bcnt_49_CYINIT_888 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_215,
      O => tx_output_bcnt_49_CYINIT
    );
  tx_output_bcnt_51_LOGIC_ONE_889 : X_ONE
    port map (
      O => tx_output_bcnt_51_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_218_890 : X_MUX2
    port map (
      IA => tx_output_bcnt_51_LOGIC_ONE,
      IB => tx_output_bcnt_51_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_53,
      O => tx_output_bcnt_inst_cy_218
    );
  tx_output_bcnt_inst_sum_184_891 : X_XOR2
    port map (
      I0 => tx_output_bcnt_51_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_53,
      O => tx_output_bcnt_inst_sum_184
    );
  tx_output_bcnt_inst_lut3_531 : X_LUT4
    generic map(
      INIT => X"550F"
    )
    port map (
      ADR0 => q2(13),
      ADR1 => VCC,
      ADR2 => tx_output_bcnt_51,
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_53
    );
  tx_output_bcnt_inst_lut3_541 : X_LUT4
    generic map(
      INIT => X"1B1B"
    )
    port map (
      ADR0 => tx_output_cs_FFd12,
      ADR1 => tx_output_bcnt_52,
      ADR2 => q2(14),
      ADR3 => VCC,
      O => tx_output_bcnt_inst_lut3_54
    );
  tx_output_bcnt_51_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_51_CYMUXG,
      O => tx_output_bcnt_inst_cy_219
    );
  tx_output_bcnt_inst_cy_219_892 : X_MUX2
    port map (
      IA => tx_output_bcnt_51_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_218,
      SEL => tx_output_bcnt_inst_lut3_54,
      O => tx_output_bcnt_51_CYMUXG
    );
  tx_output_bcnt_inst_sum_185_893 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_218,
      I1 => tx_output_bcnt_inst_lut3_54,
      O => tx_output_bcnt_inst_sum_185
    );
  tx_output_bcnt_51_CYINIT_894 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_217,
      O => tx_output_bcnt_51_CYINIT
    );
  tx_output_bcnt_inst_sum_186_895 : X_XOR2
    port map (
      I0 => tx_output_bcnt_53_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_55,
      O => tx_output_bcnt_inst_sum_186
    );
  tx_output_bcnt_inst_lut3_551 : X_LUT4
    generic map(
      INIT => X"550F"
    )
    port map (
      ADR0 => q2(15),
      ADR1 => VCC,
      ADR2 => tx_output_bcnt_53,
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_55
    );
  tx_output_bcnt_53_CYINIT_896 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_219,
      O => tx_output_bcnt_53_CYINIT
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ONE_897 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ZERO_898 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_177_899 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(16),
      ADR1 => rx_input_memio_addrchk_macaddrl(17),
      ADR2 => rx_input_memio_addrchk_datal(16),
      ADR3 => rx_input_memio_addrchk_datal(17),
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(19),
      ADR1 => rx_input_memio_addrchk_macaddrl(18),
      ADR2 => rx_input_memio_addrchk_datal(18),
      ADR3 => rx_input_memio_addrchk_datal(19),
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_900 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_CYMUXG
    );
  rx_input_fifo_fifo_BU115 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3240,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N2406_FFX_RST,
      O => rx_input_fifo_fifo_N2406
    );
  rx_input_fifo_fifo_N2406_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2406_FFX_RST
    );
  rx_input_memio_addrchk_lmaceq_3_LOGIC_ZERO_901 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_3_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_179_902 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_3_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_3_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(20),
      ADR1 => rx_input_memio_addrchk_macaddrl(21),
      ADR2 => rx_input_memio_addrchk_datal(21),
      ADR3 => rx_input_memio_addrchk_datal(20),
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(22),
      ADR1 => rx_input_memio_addrchk_macaddrl(23),
      ADR2 => rx_input_memio_addrchk_datal(22),
      ADR3 => rx_input_memio_addrchk_datal(23),
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_3_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_3_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(3)
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_3_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_3_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_3_CYINIT_903 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_3_CYINIT
    );
  rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ONE_904 : X_ONE
    port map (
      O => rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ONE
    );
  rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ZERO_905 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ZERO
    );
  rx_output_Mcompar_n0017_inst_cy_78_906 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ONE,
      SEL => rx_output_Mcompar_n0017_inst_lut4_0,
      O => rx_output_Mcompar_n0017_inst_cy_78
    );
  rx_output_Mcompar_n0017_inst_lut4_01 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_output_bpl(1),
      ADR1 => rx_output_bpl(0),
      ADR2 => rxbp(1),
      ADR3 => rxbp(0),
      O => rx_output_Mcompar_n0017_inst_lut4_0
    );
  rx_output_Mcompar_n0017_inst_lut4_11 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_output_bpl(2),
      ADR1 => rx_output_bpl(3),
      ADR2 => rxbp(2),
      ADR3 => rxbp(3),
      O => rx_output_Mcompar_n0017_inst_lut4_1
    );
  rx_output_Mcompar_n0017_inst_cy_79_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_79_CYMUXG,
      O => rx_output_Mcompar_n0017_inst_cy_79
    );
  rx_output_Mcompar_n0017_inst_cy_79_907 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_78,
      SEL => rx_output_Mcompar_n0017_inst_lut4_1,
      O => rx_output_Mcompar_n0017_inst_cy_79_CYMUXG
    );
  rx_output_Mcompar_n0017_inst_cy_81_LOGIC_ZERO_908 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0017_inst_cy_81_LOGIC_ZERO
    );
  rx_output_Mcompar_n0017_inst_cy_80_909 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_81_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_81_CYINIT,
      SEL => rx_output_Mcompar_n0017_inst_lut4_2,
      O => rx_output_Mcompar_n0017_inst_cy_80
    );
  rx_output_Mcompar_n0017_inst_lut4_21 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rxbp(5),
      ADR1 => rx_output_bpl(5),
      ADR2 => rx_output_bpl(4),
      ADR3 => rxbp(4),
      O => rx_output_Mcompar_n0017_inst_lut4_2
    );
  rx_output_Mcompar_n0017_inst_lut4_31 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rxbp(7),
      ADR1 => rxbp(6),
      ADR2 => rx_output_bpl(7),
      ADR3 => rx_output_bpl(6),
      O => rx_output_Mcompar_n0017_inst_lut4_3
    );
  rx_output_Mcompar_n0017_inst_cy_81_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_81_CYMUXG,
      O => rx_output_Mcompar_n0017_inst_cy_81
    );
  rx_output_Mcompar_n0017_inst_cy_81_910 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_81_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_80,
      SEL => rx_output_Mcompar_n0017_inst_lut4_3,
      O => rx_output_Mcompar_n0017_inst_cy_81_CYMUXG
    );
  rx_output_Mcompar_n0017_inst_cy_81_CYINIT_911 : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_79,
      O => rx_output_Mcompar_n0017_inst_cy_81_CYINIT
    );
  rx_output_Mcompar_n0017_inst_cy_83_LOGIC_ZERO_912 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0017_inst_cy_83_LOGIC_ZERO
    );
  rx_output_Mcompar_n0017_inst_cy_82_913 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_83_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_83_CYINIT,
      SEL => rx_output_Mcompar_n0017_inst_lut4_4,
      O => rx_output_Mcompar_n0017_inst_cy_82
    );
  rx_output_Mcompar_n0017_inst_lut4_41 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_output_bpl(8),
      ADR1 => rx_output_bpl(9),
      ADR2 => rxbp(8),
      ADR3 => rxbp(9),
      O => rx_output_Mcompar_n0017_inst_lut4_4
    );
  rx_output_Mcompar_n0017_inst_lut4_51 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_output_bpl(10),
      ADR1 => rxbp(10),
      ADR2 => rx_output_bpl(11),
      ADR3 => rxbp(11),
      O => rx_output_Mcompar_n0017_inst_lut4_5
    );
  rx_output_Mcompar_n0017_inst_cy_83_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_83_CYMUXG,
      O => rx_output_Mcompar_n0017_inst_cy_83
    );
  rx_output_Mcompar_n0017_inst_cy_83_914 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_83_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_82,
      SEL => rx_output_Mcompar_n0017_inst_lut4_5,
      O => rx_output_Mcompar_n0017_inst_cy_83_CYMUXG
    );
  rx_output_Mcompar_n0017_inst_cy_83_CYINIT_915 : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_81,
      O => rx_output_Mcompar_n0017_inst_cy_83_CYINIT
    );
  rx_output_n0017_LOGIC_ZERO_916 : X_ZERO
    port map (
      O => rx_output_n0017_LOGIC_ZERO
    );
  rx_output_Mcompar_n0017_inst_cy_84_917 : X_MUX2
    port map (
      IA => rx_output_n0017_LOGIC_ZERO,
      IB => rx_output_n0017_CYINIT,
      SEL => rx_output_Mcompar_n0017_inst_lut4_6,
      O => rx_output_Mcompar_n0017_inst_cy_84
    );
  rx_output_Mcompar_n0017_inst_lut4_61 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_output_bpl(13),
      ADR1 => rx_output_bpl(12),
      ADR2 => rxbp(12),
      ADR3 => rxbp(13),
      O => rx_output_Mcompar_n0017_inst_lut4_6
    );
  rx_output_Mcompar_n0017_inst_lut4_71 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rxbp(15),
      ADR1 => rx_output_bpl(14),
      ADR2 => rx_output_bpl(15),
      ADR3 => rxbp(14),
      O => rx_output_Mcompar_n0017_inst_lut4_7
    );
  rx_output_n0017_COUTUSED : X_BUF
    port map (
      I => rx_output_n0017_CYMUXG,
      O => rx_output_n0017
    );
  rx_output_Mcompar_n0017_inst_cy_85 : X_MUX2
    port map (
      IA => rx_output_n0017_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_84,
      SEL => rx_output_Mcompar_n0017_inst_lut4_7,
      O => rx_output_n0017_CYMUXG
    );
  rx_output_n0017_CYINIT_918 : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_83,
      O => rx_output_n0017_CYINIT
    );
  rx_fifocheck_diff_0_LOGIC_ONE_919 : X_ONE
    port map (
      O => rx_fifocheck_diff_0_LOGIC_ONE
    );
  rx_fifocheck_Msub_n0001_inst_cy_161_920 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(0),
      IB => rx_fifocheck_diff_0_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_111,
      O => rx_fifocheck_Msub_n0001_inst_cy_161
    );
  rx_fifocheck_Msub_n0001_inst_sum_143 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_0_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_111,
      O => rx_fifocheck_n0001(0)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1111 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_bpl(0),
      O => rx_fifocheck_Msub_n0001_inst_lut2_111
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1121 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(1),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(1),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_112
    );
  rx_fifocheck_diff_0_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_0_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_162
    );
  rx_fifocheck_Msub_n0001_inst_cy_162_921 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(1),
      IB => rx_fifocheck_Msub_n0001_inst_cy_161,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_112,
      O => rx_fifocheck_diff_0_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_144 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_161,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_112,
      O => rx_fifocheck_n0001(1)
    );
  rx_fifocheck_diff_0_CYINIT_922 : X_BUF
    port map (
      I => rx_fifocheck_diff_0_LOGIC_ONE,
      O => rx_fifocheck_diff_0_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_163_923 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(2),
      IB => rx_fifocheck_diff_2_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_113,
      O => rx_fifocheck_Msub_n0001_inst_cy_163
    );
  rx_fifocheck_Msub_n0001_inst_sum_145 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_2_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_113,
      O => rx_fifocheck_n0001(2)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1131 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(2),
      ADR1 => rx_fifocheck_bpl(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_113
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1141 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_bpl(3),
      O => rx_fifocheck_Msub_n0001_inst_lut2_114
    );
  rx_fifocheck_diff_2_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_2_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_164
    );
  rx_fifocheck_Msub_n0001_inst_cy_164_924 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(3),
      IB => rx_fifocheck_Msub_n0001_inst_cy_163,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_114,
      O => rx_fifocheck_diff_2_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_146 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_163,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_114,
      O => rx_fifocheck_n0001(3)
    );
  rx_fifocheck_diff_2_CYINIT_925 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_162,
      O => rx_fifocheck_diff_2_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_165_926 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(4),
      IB => rx_fifocheck_diff_4_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_115,
      O => rx_fifocheck_Msub_n0001_inst_cy_165
    );
  rx_fifocheck_Msub_n0001_inst_sum_147 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_4_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_115,
      O => rx_fifocheck_n0001(4)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1151 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(4),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(4),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_115
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1161 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_bpl(5),
      O => rx_fifocheck_Msub_n0001_inst_lut2_116
    );
  rx_fifocheck_diff_4_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_4_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_166
    );
  rx_fifocheck_Msub_n0001_inst_cy_166_927 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(5),
      IB => rx_fifocheck_Msub_n0001_inst_cy_165,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_116,
      O => rx_fifocheck_diff_4_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_148 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_165,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_116,
      O => rx_fifocheck_n0001(5)
    );
  rx_fifocheck_diff_4_CYINIT_928 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_164,
      O => rx_fifocheck_diff_4_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_167_929 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(6),
      IB => rx_fifocheck_diff_6_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_117,
      O => rx_fifocheck_Msub_n0001_inst_cy_167
    );
  rx_fifocheck_Msub_n0001_inst_sum_149 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_6_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_117,
      O => rx_fifocheck_n0001(6)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1171 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(6),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(6),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_117
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1181 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(7),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(7),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_118
    );
  rx_fifocheck_diff_6_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_6_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_168
    );
  rx_fifocheck_Msub_n0001_inst_cy_168_930 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(7),
      IB => rx_fifocheck_Msub_n0001_inst_cy_167,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_118,
      O => rx_fifocheck_diff_6_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_150 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_167,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_118,
      O => rx_fifocheck_n0001(7)
    );
  rx_fifocheck_diff_6_CYINIT_931 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_166,
      O => rx_fifocheck_diff_6_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_169_932 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(8),
      IB => rx_fifocheck_diff_8_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_119,
      O => rx_fifocheck_Msub_n0001_inst_cy_169
    );
  rx_fifocheck_Msub_n0001_inst_sum_151 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_8_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_119,
      O => rx_fifocheck_n0001(8)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1191 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(8),
      ADR1 => rx_fifocheck_bpl(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_119
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1201 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_bpl(9),
      O => rx_fifocheck_Msub_n0001_inst_lut2_120
    );
  rx_fifocheck_diff_8_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_8_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_170
    );
  rx_fifocheck_Msub_n0001_inst_cy_170_933 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(9),
      IB => rx_fifocheck_Msub_n0001_inst_cy_169,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_120,
      O => rx_fifocheck_diff_8_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_152 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_169,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_120,
      O => rx_fifocheck_n0001(9)
    );
  rx_fifocheck_diff_8_CYINIT_934 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_168,
      O => rx_fifocheck_diff_8_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_171_935 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(10),
      IB => rx_fifocheck_diff_10_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_121,
      O => rx_fifocheck_Msub_n0001_inst_cy_171
    );
  rx_fifocheck_Msub_n0001_inst_sum_153 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_10_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_121,
      O => rx_fifocheck_n0001(10)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1211 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(10),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_bpl(10),
      O => rx_fifocheck_Msub_n0001_inst_lut2_121
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1221 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(11),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_bpl(11),
      O => rx_fifocheck_Msub_n0001_inst_lut2_122
    );
  rx_fifocheck_diff_10_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_10_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_172
    );
  rx_fifocheck_Msub_n0001_inst_cy_172_936 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(11),
      IB => rx_fifocheck_Msub_n0001_inst_cy_171,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_122,
      O => rx_fifocheck_diff_10_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_154 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_171,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_122,
      O => rx_fifocheck_n0001(11)
    );
  rx_fifocheck_diff_10_CYINIT_937 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_170,
      O => rx_fifocheck_diff_10_CYINIT
    );
  rx_input_fifo_fifo_BU184 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2486,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N2505_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N2506
    );
  rx_input_fifo_fifo_N2505_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N2505_FFY_SET
    );
  rx_fifocheck_Msub_n0001_inst_cy_173_938 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(12),
      IB => rx_fifocheck_diff_12_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_123,
      O => rx_fifocheck_Msub_n0001_inst_cy_173
    );
  rx_fifocheck_Msub_n0001_inst_sum_155 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_12_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_123,
      O => rx_fifocheck_n0001(12)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1231 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(12),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(12),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_123
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1241 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(13),
      ADR1 => rx_fifocheck_bpl(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_124
    );
  rx_fifocheck_diff_12_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_12_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_174
    );
  rx_fifocheck_Msub_n0001_inst_cy_174_939 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(13),
      IB => rx_fifocheck_Msub_n0001_inst_cy_173,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_124,
      O => rx_fifocheck_diff_12_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_156 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_173,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_124,
      O => rx_fifocheck_n0001(13)
    );
  rx_fifocheck_diff_12_CYINIT_940 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_172,
      O => rx_fifocheck_diff_12_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_175_941 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(14),
      IB => rx_fifocheck_diff_14_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_125,
      O => rx_fifocheck_Msub_n0001_inst_cy_175
    );
  rx_fifocheck_Msub_n0001_inst_sum_157 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_14_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_125,
      O => rx_fifocheck_n0001(14)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1251 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(14),
      ADR1 => rx_fifocheck_bpl(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_125
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1261 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(15),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(15),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_126
    );
  rx_fifocheck_Msub_n0001_inst_sum_158 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_175,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_126,
      O => rx_fifocheck_n0001(15)
    );
  rx_fifocheck_diff_14_CYINIT_942 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_174,
      O => rx_fifocheck_diff_14_CYINIT
    );
  tx_fifocheck_diff_0_LOGIC_ONE_943 : X_ONE
    port map (
      O => tx_fifocheck_diff_0_LOGIC_ONE
    );
  tx_fifocheck_Msub_n0001_inst_cy_161_944 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(0),
      IB => tx_fifocheck_diff_0_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_111,
      O => tx_fifocheck_Msub_n0001_inst_cy_161
    );
  tx_fifocheck_Msub_n0001_inst_sum_143 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_0_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_111,
      O => tx_fifocheck_n0001(0)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1111 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(0),
      O => tx_fifocheck_Msub_n0001_inst_lut2_111
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1121 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(1),
      ADR1 => tx_fifocheck_bpl(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_112
    );
  tx_fifocheck_diff_0_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_0_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_162
    );
  tx_fifocheck_Msub_n0001_inst_cy_162_945 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(1),
      IB => tx_fifocheck_Msub_n0001_inst_cy_161,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_112,
      O => tx_fifocheck_diff_0_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_144 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_161,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_112,
      O => tx_fifocheck_n0001(1)
    );
  tx_fifocheck_diff_0_CYINIT_946 : X_BUF
    port map (
      I => tx_fifocheck_diff_0_LOGIC_ONE,
      O => tx_fifocheck_diff_0_CYINIT
    );
  tx_fifocheck_diff_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_2_FFY_RST
    );
  tx_fifocheck_diff_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_2_FFY_RST,
      O => tx_fifocheck_diff(3)
    );
  tx_fifocheck_Msub_n0001_inst_cy_163_947 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(2),
      IB => tx_fifocheck_diff_2_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_113,
      O => tx_fifocheck_Msub_n0001_inst_cy_163
    );
  tx_fifocheck_Msub_n0001_inst_sum_145 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_2_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_113,
      O => tx_fifocheck_n0001(2)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1131 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(2),
      ADR1 => VCC,
      ADR2 => tx_fifocheck_bpl(2),
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_113
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1141 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(3),
      ADR1 => VCC,
      ADR2 => tx_fifocheck_bpl(3),
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_114
    );
  tx_fifocheck_diff_2_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_2_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_164
    );
  tx_fifocheck_Msub_n0001_inst_cy_164_948 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(3),
      IB => tx_fifocheck_Msub_n0001_inst_cy_163,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_114,
      O => tx_fifocheck_diff_2_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_146 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_163,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_114,
      O => tx_fifocheck_n0001(3)
    );
  tx_fifocheck_diff_2_CYINIT_949 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_162,
      O => tx_fifocheck_diff_2_CYINIT
    );
  tx_fifocheck_diff_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_4_FFY_RST
    );
  tx_fifocheck_diff_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_4_FFY_RST,
      O => tx_fifocheck_diff(5)
    );
  tx_fifocheck_Msub_n0001_inst_cy_165_950 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(4),
      IB => tx_fifocheck_diff_4_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_115,
      O => tx_fifocheck_Msub_n0001_inst_cy_165
    );
  tx_fifocheck_Msub_n0001_inst_sum_147 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_4_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_115,
      O => tx_fifocheck_n0001(4)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1151 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(4),
      ADR1 => VCC,
      ADR2 => tx_fifocheck_bpl(4),
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_115
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1161 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(5),
      O => tx_fifocheck_Msub_n0001_inst_lut2_116
    );
  tx_fifocheck_diff_4_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_4_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_166
    );
  tx_fifocheck_Msub_n0001_inst_cy_166_951 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(5),
      IB => tx_fifocheck_Msub_n0001_inst_cy_165,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_116,
      O => tx_fifocheck_diff_4_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_148 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_165,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_116,
      O => tx_fifocheck_n0001(5)
    );
  tx_fifocheck_diff_4_CYINIT_952 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_164,
      O => tx_fifocheck_diff_4_CYINIT
    );
  tx_fifocheck_diff_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_6_FFY_RST
    );
  tx_fifocheck_diff_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_6_FFY_RST,
      O => tx_fifocheck_diff(7)
    );
  tx_fifocheck_Msub_n0001_inst_cy_167_953 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(6),
      IB => tx_fifocheck_diff_6_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_117,
      O => tx_fifocheck_Msub_n0001_inst_cy_167
    );
  tx_fifocheck_Msub_n0001_inst_sum_149 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_6_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_117,
      O => tx_fifocheck_n0001(6)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1171 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(6),
      ADR1 => tx_fifocheck_bpl(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_117
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1181 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(7),
      ADR1 => VCC,
      ADR2 => tx_fifocheck_bpl(7),
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_118
    );
  tx_fifocheck_diff_6_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_6_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_168
    );
  tx_fifocheck_Msub_n0001_inst_cy_168_954 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(7),
      IB => tx_fifocheck_Msub_n0001_inst_cy_167,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_118,
      O => tx_fifocheck_diff_6_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_150 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_167,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_118,
      O => tx_fifocheck_n0001(7)
    );
  tx_fifocheck_diff_6_CYINIT_955 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_166,
      O => tx_fifocheck_diff_6_CYINIT
    );
  tx_fifocheck_diff_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_8_FFY_RST
    );
  tx_fifocheck_diff_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_8_FFY_RST,
      O => tx_fifocheck_diff(9)
    );
  tx_fifocheck_Msub_n0001_inst_cy_169_956 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(8),
      IB => tx_fifocheck_diff_8_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_119,
      O => tx_fifocheck_Msub_n0001_inst_cy_169
    );
  tx_fifocheck_Msub_n0001_inst_sum_151 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_8_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_119,
      O => tx_fifocheck_n0001(8)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1191 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(8),
      O => tx_fifocheck_Msub_n0001_inst_lut2_119
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1201 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(9),
      ADR1 => tx_fifocheck_bpl(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_120
    );
  tx_fifocheck_diff_8_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_8_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_170
    );
  tx_fifocheck_Msub_n0001_inst_cy_170_957 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(9),
      IB => tx_fifocheck_Msub_n0001_inst_cy_169,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_120,
      O => tx_fifocheck_diff_8_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_152 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_169,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_120,
      O => tx_fifocheck_n0001(9)
    );
  tx_fifocheck_diff_8_CYINIT_958 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_168,
      O => tx_fifocheck_diff_8_CYINIT
    );
  tx_fifocheck_diff_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_10_FFY_RST
    );
  tx_fifocheck_diff_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_10_FFY_RST,
      O => tx_fifocheck_diff(11)
    );
  tx_fifocheck_Msub_n0001_inst_cy_171_959 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(10),
      IB => tx_fifocheck_diff_10_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_121,
      O => tx_fifocheck_Msub_n0001_inst_cy_171
    );
  tx_fifocheck_Msub_n0001_inst_sum_153 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_10_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_121,
      O => tx_fifocheck_n0001(10)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1211 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(10),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(10),
      O => tx_fifocheck_Msub_n0001_inst_lut2_121
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1221 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(11),
      ADR1 => tx_fifocheck_bpl(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_122
    );
  tx_fifocheck_diff_10_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_10_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_172
    );
  tx_fifocheck_Msub_n0001_inst_cy_172_960 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(11),
      IB => tx_fifocheck_Msub_n0001_inst_cy_171,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_122,
      O => tx_fifocheck_diff_10_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_154 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_171,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_122,
      O => tx_fifocheck_n0001(11)
    );
  tx_fifocheck_diff_10_CYINIT_961 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_170,
      O => tx_fifocheck_diff_10_CYINIT
    );
  tx_fifocheck_diff_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_12_FFY_RST
    );
  tx_fifocheck_diff_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_12_FFY_RST,
      O => tx_fifocheck_diff(13)
    );
  tx_fifocheck_Msub_n0001_inst_cy_173_962 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(12),
      IB => tx_fifocheck_diff_12_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_123,
      O => tx_fifocheck_Msub_n0001_inst_cy_173
    );
  tx_fifocheck_Msub_n0001_inst_sum_155 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_12_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_123,
      O => tx_fifocheck_n0001(12)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1231 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(12),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(12),
      O => tx_fifocheck_Msub_n0001_inst_lut2_123
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1241 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(13),
      O => tx_fifocheck_Msub_n0001_inst_lut2_124
    );
  tx_fifocheck_diff_12_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_12_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_174
    );
  tx_fifocheck_Msub_n0001_inst_cy_174_963 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(13),
      IB => tx_fifocheck_Msub_n0001_inst_cy_173,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_124,
      O => tx_fifocheck_diff_12_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_156 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_173,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_124,
      O => tx_fifocheck_n0001(13)
    );
  tx_fifocheck_diff_12_CYINIT_964 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_172,
      O => tx_fifocheck_diff_12_CYINIT
    );
  tx_fifocheck_diff_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_14_FFY_RST
    );
  tx_fifocheck_diff_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_14_FFY_RST,
      O => tx_fifocheck_diff(15)
    );
  tx_fifocheck_Msub_n0001_inst_cy_175_965 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(14),
      IB => tx_fifocheck_diff_14_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_125,
      O => tx_fifocheck_Msub_n0001_inst_cy_175
    );
  tx_fifocheck_Msub_n0001_inst_sum_157 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_14_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_125,
      O => tx_fifocheck_n0001(14)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1251 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(14),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(14),
      O => tx_fifocheck_Msub_n0001_inst_lut2_125
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1261 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(15),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(15),
      O => tx_fifocheck_Msub_n0001_inst_lut2_126
    );
  tx_fifocheck_Msub_n0001_inst_sum_158 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_175,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_126,
      O => tx_fifocheck_n0001(15)
    );
  tx_fifocheck_diff_14_CYINIT_966 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_174,
      O => tx_fifocheck_diff_14_CYINIT
    );
  mac_control_ledtx_cnt_142_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_142_FFY_RST
    );
  mac_control_ledtx_cnt_142_967 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_289,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_142_FFY_RST,
      O => mac_control_ledtx_cnt_142
    );
  mac_control_ledtx_cnt_142_LOGIC_ONE_968 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_142_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_327_969 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_8,
      IB => mac_control_ledtx_cnt_142_LOGIC_ONE,
      SEL => mac_control_ledtx_rst_rt,
      O => mac_control_ledtx_cnt_inst_cy_327
    );
  mac_control_ledtx_rst_rt_970 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_8,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_ledtx_rst,
      O => mac_control_ledtx_rst_rt
    );
  mac_control_ledtx_cnt_inst_lut3_2241 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_3,
      ADR1 => mac_control_ledtx_cnt_142,
      ADR2 => mac_control_ledtx_rst,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_224
    );
  mac_control_ledtx_cnt_142_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_142_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_328
    );
  mac_control_ledtx_cnt_inst_cy_328_971 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_3,
      IB => mac_control_ledtx_cnt_inst_cy_327,
      SEL => mac_control_ledtx_cnt_inst_lut3_224,
      O => mac_control_ledtx_cnt_142_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_289_972 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_327,
      I1 => mac_control_ledtx_cnt_inst_lut3_224,
      O => mac_control_ledtx_cnt_inst_sum_289
    );
  mac_control_ledtx_cnt_143_LOGIC_ONE_973 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_143_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_329_974 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_143_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_143_CYINIT,
      SEL => mac_control_ledtx_cnt_inst_lut3_225,
      O => mac_control_ledtx_cnt_inst_cy_329
    );
  mac_control_ledtx_cnt_inst_sum_290_975 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_143_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_225,
      O => mac_control_ledtx_cnt_inst_sum_290
    );
  mac_control_ledtx_cnt_inst_lut3_2251 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_ledtx_rst,
      ADR1 => mac_control_ledtx_cnt_143,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_225
    );
  mac_control_ledtx_cnt_inst_lut3_2261 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledtx_cnt_144,
      ADR3 => mac_control_ledtx_rst,
      O => mac_control_ledtx_cnt_inst_lut3_226
    );
  mac_control_ledtx_cnt_143_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_143_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_330
    );
  mac_control_ledtx_cnt_inst_cy_330_976 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_143_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_inst_cy_329,
      SEL => mac_control_ledtx_cnt_inst_lut3_226,
      O => mac_control_ledtx_cnt_143_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_291_977 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_329,
      I1 => mac_control_ledtx_cnt_inst_lut3_226,
      O => mac_control_ledtx_cnt_inst_sum_291
    );
  mac_control_ledtx_cnt_143_CYINIT_978 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_328,
      O => mac_control_ledtx_cnt_143_CYINIT
    );
  mac_control_ledtx_cnt_145_LOGIC_ONE_979 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_145_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_331_980 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_145_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_145_CYINIT,
      SEL => mac_control_ledtx_cnt_inst_lut3_227,
      O => mac_control_ledtx_cnt_inst_cy_331
    );
  mac_control_ledtx_cnt_inst_sum_292_981 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_145_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_227,
      O => mac_control_ledtx_cnt_inst_sum_292
    );
  mac_control_ledtx_cnt_inst_lut3_2271 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledtx_rst,
      ADR2 => VCC,
      ADR3 => mac_control_ledtx_cnt_145,
      O => mac_control_ledtx_cnt_inst_lut3_227
    );
  mac_control_ledtx_cnt_inst_lut3_2281 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => mac_control_ledtx_rst,
      ADR1 => VCC,
      ADR2 => mac_control_ledtx_cnt_146,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_228
    );
  mac_control_ledtx_cnt_145_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_145_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_332
    );
  mac_control_ledtx_cnt_inst_cy_332_982 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_145_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_inst_cy_331,
      SEL => mac_control_ledtx_cnt_inst_lut3_228,
      O => mac_control_ledtx_cnt_145_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_293_983 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_331,
      I1 => mac_control_ledtx_cnt_inst_lut3_228,
      O => mac_control_ledtx_cnt_inst_sum_293
    );
  mac_control_ledtx_cnt_145_CYINIT_984 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_330,
      O => mac_control_ledtx_cnt_145_CYINIT
    );
  mac_control_ledtx_cnt_147_LOGIC_ONE_985 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_147_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_333_986 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_147_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_147_CYINIT,
      SEL => mac_control_ledtx_cnt_inst_lut3_229,
      O => mac_control_ledtx_cnt_inst_cy_333
    );
  mac_control_ledtx_cnt_inst_sum_294_987 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_147_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_229,
      O => mac_control_ledtx_cnt_inst_sum_294
    );
  mac_control_ledtx_cnt_inst_lut3_2291 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledtx_rst,
      ADR2 => VCC,
      ADR3 => mac_control_ledtx_cnt_147,
      O => mac_control_ledtx_cnt_inst_lut3_229
    );
  mac_control_ledtx_cnt_inst_lut3_2301 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledtx_rst,
      ADR2 => mac_control_ledtx_cnt_148,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_230
    );
  mac_control_ledtx_cnt_147_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_147_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_334
    );
  mac_control_ledtx_cnt_inst_cy_334_988 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_147_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_inst_cy_333,
      SEL => mac_control_ledtx_cnt_inst_lut3_230,
      O => mac_control_ledtx_cnt_147_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_295_989 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_333,
      I1 => mac_control_ledtx_cnt_inst_lut3_230,
      O => mac_control_ledtx_cnt_inst_sum_295
    );
  mac_control_ledtx_cnt_147_CYINIT_990 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_332,
      O => mac_control_ledtx_cnt_147_CYINIT
    );
  mac_control_ledtx_cnt_149_LOGIC_ONE_991 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_149_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_335_992 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_149_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_149_CYINIT,
      SEL => mac_control_ledtx_cnt_inst_lut3_231,
      O => mac_control_ledtx_cnt_inst_cy_335
    );
  mac_control_ledtx_cnt_inst_sum_296_993 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_149_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_231,
      O => mac_control_ledtx_cnt_inst_sum_296
    );
  mac_control_ledtx_cnt_inst_lut3_2311 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_149,
      ADR1 => mac_control_ledtx_rst,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_231
    );
  mac_control_ledtx_cnt_inst_lut3_2321 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledtx_rst,
      ADR3 => mac_control_ledtx_cnt_150,
      O => mac_control_ledtx_cnt_inst_lut3_232
    );
  mac_control_ledtx_cnt_149_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_149_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_336
    );
  mac_control_ledtx_cnt_inst_cy_336_994 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_149_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_inst_cy_335,
      SEL => mac_control_ledtx_cnt_inst_lut3_232,
      O => mac_control_ledtx_cnt_149_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_297_995 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_335,
      I1 => mac_control_ledtx_cnt_inst_lut3_232,
      O => mac_control_ledtx_cnt_inst_sum_297
    );
  mac_control_ledtx_cnt_149_CYINIT_996 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_334,
      O => mac_control_ledtx_cnt_149_CYINIT
    );
  mac_control_ledtx_cnt_151_LOGIC_ONE_997 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_151_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_337_998 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_151_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_151_CYINIT,
      SEL => mac_control_ledtx_cnt_inst_lut3_233,
      O => mac_control_ledtx_cnt_inst_cy_337
    );
  mac_control_ledtx_cnt_inst_sum_298_999 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_151_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_233,
      O => mac_control_ledtx_cnt_inst_sum_298
    );
  mac_control_ledtx_cnt_inst_lut3_2331 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledtx_rst,
      ADR2 => mac_control_ledtx_cnt_151,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_233
    );
  mac_control_ledtx_cnt_inst_lut3_2341 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_152,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_ledtx_rst,
      O => mac_control_ledtx_cnt_inst_lut3_234
    );
  mac_control_ledtx_cnt_151_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_151_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_338
    );
  mac_control_ledtx_cnt_inst_cy_338_1000 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_151_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_inst_cy_337,
      SEL => mac_control_ledtx_cnt_inst_lut3_234,
      O => mac_control_ledtx_cnt_151_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_299_1001 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_337,
      I1 => mac_control_ledtx_cnt_inst_lut3_234,
      O => mac_control_ledtx_cnt_inst_sum_299
    );
  mac_control_ledtx_cnt_151_CYINIT_1002 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_336,
      O => mac_control_ledtx_cnt_151_CYINIT
    );
  mac_control_ledtx_cnt_inst_sum_300_1003 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_153_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_235,
      O => mac_control_ledtx_cnt_inst_sum_300
    );
  mac_control_ledtx_cnt_inst_lut3_2351 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_153,
      ADR1 => mac_control_ledtx_rst,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_235
    );
  mac_control_ledtx_cnt_153_CYINIT_1004 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_338,
      O => mac_control_ledtx_cnt_153_CYINIT
    );
  rx_output_fifo_N17_LOGIC_ZERO_1005 : X_ZERO
    port map (
      O => rx_output_fifo_N17_LOGIC_ZERO
    );
  rx_output_fifo_BU38 : X_MUX2
    port map (
      IA => rx_output_fifo_N17,
      IB => rx_output_fifo_N17_CYINIT,
      SEL => rx_output_fifo_N1912,
      O => rx_output_fifo_N1914
    );
  rx_output_fifo_BU39 : X_XOR2
    port map (
      I0 => rx_output_fifo_N17_CYINIT,
      I1 => rx_output_fifo_N1912,
      O => rx_output_fifo_N1904
    );
  rx_output_fifo_BU37 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_output_fifo_N17,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N1912
    );
  rx_output_fifo_N17_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N16,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N17_GROM
    );
  rx_output_fifo_N17_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N17_CYMUXG,
      O => rx_output_fifo_N1919
    );
  rx_output_fifo_BU44 : X_MUX2
    port map (
      IA => rx_output_fifo_N16,
      IB => rx_output_fifo_N1914,
      SEL => rx_output_fifo_N17_GROM,
      O => rx_output_fifo_N17_CYMUXG
    );
  rx_output_fifo_BU45 : X_XOR2
    port map (
      I0 => rx_output_fifo_N1914,
      I1 => rx_output_fifo_N17_GROM,
      O => rx_output_fifo_N1905
    );
  rx_output_fifo_N17_CYINIT_1006 : X_BUF
    port map (
      I => rx_output_fifo_N17_LOGIC_ZERO,
      O => rx_output_fifo_N17_CYINIT
    );
  rx_output_fifo_BU50 : X_MUX2
    port map (
      IA => rx_output_fifo_N15,
      IB => rx_output_fifo_N15_CYINIT,
      SEL => rx_output_fifo_N15_FROM,
      O => rx_output_fifo_N1924
    );
  rx_output_fifo_BU51 : X_XOR2
    port map (
      I0 => rx_output_fifo_N15_CYINIT,
      I1 => rx_output_fifo_N15_FROM,
      O => rx_output_fifo_N1906
    );
  rx_output_fifo_N15_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N15,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N15_FROM
    );
  rx_output_fifo_N15_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N14,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N15_GROM
    );
  rx_output_fifo_N15_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N15_CYMUXG,
      O => rx_output_fifo_N1929
    );
  rx_output_fifo_BU56 : X_MUX2
    port map (
      IA => rx_output_fifo_N14,
      IB => rx_output_fifo_N1924,
      SEL => rx_output_fifo_N15_GROM,
      O => rx_output_fifo_N15_CYMUXG
    );
  rx_output_fifo_BU57 : X_XOR2
    port map (
      I0 => rx_output_fifo_N1924,
      I1 => rx_output_fifo_N15_GROM,
      O => rx_output_fifo_N1907
    );
  rx_output_fifo_N15_CYINIT_1007 : X_BUF
    port map (
      I => rx_output_fifo_N1919,
      O => rx_output_fifo_N15_CYINIT
    );
  rx_output_fifo_BU62 : X_MUX2
    port map (
      IA => rx_output_fifo_N13,
      IB => rx_output_fifo_N13_CYINIT,
      SEL => rx_output_fifo_N13_FROM,
      O => rx_output_fifo_N1934
    );
  rx_output_fifo_BU63 : X_XOR2
    port map (
      I0 => rx_output_fifo_N13_CYINIT,
      I1 => rx_output_fifo_N13_FROM,
      O => rx_output_fifo_N1908
    );
  rx_output_fifo_N13_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N13,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N13_FROM
    );
  rx_output_fifo_N13_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N12,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N13_GROM
    );
  rx_output_fifo_N13_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N13_CYMUXG,
      O => rx_output_fifo_N1939
    );
  rx_output_fifo_BU68 : X_MUX2
    port map (
      IA => rx_output_fifo_N12,
      IB => rx_output_fifo_N1934,
      SEL => rx_output_fifo_N13_GROM,
      O => rx_output_fifo_N13_CYMUXG
    );
  rx_output_fifo_BU69 : X_XOR2
    port map (
      I0 => rx_output_fifo_N1934,
      I1 => rx_output_fifo_N13_GROM,
      O => rx_output_fifo_N1909
    );
  rx_output_fifo_N13_CYINIT_1008 : X_BUF
    port map (
      I => rx_output_fifo_N1929,
      O => rx_output_fifo_N13_CYINIT
    );
  rx_output_fifo_BU74 : X_MUX2
    port map (
      IA => rx_output_fifo_N11,
      IB => rx_output_fifo_N11_CYINIT,
      SEL => rx_output_fifo_N11_FROM,
      O => rx_output_fifo_N1944
    );
  rx_output_fifo_BU75 : X_XOR2
    port map (
      I0 => rx_output_fifo_N11_CYINIT,
      I1 => rx_output_fifo_N11_FROM,
      O => rx_output_fifo_N1910
    );
  rx_output_fifo_N11_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N11,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N11_FROM
    );
  rx_output_fifo_N10_rt_1009 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N10,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N10_rt
    );
  rx_output_fifo_BU80 : X_XOR2
    port map (
      I0 => rx_output_fifo_N1944,
      I1 => rx_output_fifo_N10_rt,
      O => rx_output_fifo_N1911
    );
  rx_output_fifo_N11_CYINIT_1010 : X_BUF
    port map (
      I => rx_output_fifo_N1939,
      O => rx_output_fifo_N11_CYINIT
    );
  tx_input_n0074_0_LOGIC_ONE_1011 : X_ONE
    port map (
      O => tx_input_n0074_0_LOGIC_ONE
    );
  tx_input_Msub_n0034_inst_cy_118_1012 : X_MUX2
    port map (
      IA => tx_input_CNT(0),
      IB => tx_input_n0074_0_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_95,
      O => tx_input_Msub_n0034_inst_cy_118
    );
  tx_input_Msub_n0034_inst_sum_111 : X_XOR2
    port map (
      I0 => tx_input_n0074_0_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_95,
      O => tx_input_n0074_0_XORF
    );
  tx_input_Msub_n0034_inst_lut2_951 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_95
    );
  tx_input_n0074_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_35,
      ADR1 => VCC,
      ADR2 => tx_input_CNT(1),
      ADR3 => VCC,
      O => tx_input_n0074_0_GROM
    );
  tx_input_n0074_0_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_0_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_119
    );
  tx_input_n0074_0_XUSED : X_BUF
    port map (
      I => tx_input_n0074_0_XORF,
      O => tx_input_n0074(0)
    );
  tx_input_n0074_0_YUSED : X_BUF
    port map (
      I => tx_input_n0074_0_XORG,
      O => tx_input_n0074(1)
    );
  tx_input_Msub_n0034_inst_cy_119_1013 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_35,
      IB => tx_input_Msub_n0034_inst_cy_118,
      SEL => tx_input_n0074_0_GROM,
      O => tx_input_n0074_0_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_112 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_118,
      I1 => tx_input_n0074_0_GROM,
      O => tx_input_n0074_0_XORG
    );
  tx_input_n0074_0_CYINIT_1014 : X_BUF
    port map (
      I => tx_input_n0074_0_LOGIC_ONE,
      O => tx_input_n0074_0_CYINIT
    );
  rx_input_fifo_fifo_BU53 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2805,
      CE => rx_input_fifo_fifo_N2362,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N21_FFX_RST,
      O => rx_input_fifo_fifo_N21
    );
  rx_input_fifo_fifo_N21_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N21_FFX_RST
    );
  tx_input_Msub_n0034_inst_cy_120_1015 : X_MUX2
    port map (
      IA => tx_input_CNT(2),
      IB => tx_input_n0074_2_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_97,
      O => tx_input_Msub_n0034_inst_cy_120
    );
  tx_input_Msub_n0034_inst_sum_113 : X_XOR2
    port map (
      I0 => tx_input_n0074_2_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_97,
      O => tx_input_n0074_2_XORF
    );
  tx_input_Msub_n0034_inst_lut2_971 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_97
    );
  tx_input_Msub_n0034_inst_lut2_981 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_98
    );
  tx_input_n0074_2_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_2_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_121
    );
  tx_input_n0074_2_XUSED : X_BUF
    port map (
      I => tx_input_n0074_2_XORF,
      O => tx_input_n0074(2)
    );
  tx_input_n0074_2_YUSED : X_BUF
    port map (
      I => tx_input_n0074_2_XORG,
      O => tx_input_n0074(3)
    );
  tx_input_Msub_n0034_inst_cy_121_1016 : X_MUX2
    port map (
      IA => tx_input_CNT(3),
      IB => tx_input_Msub_n0034_inst_cy_120,
      SEL => tx_input_Msub_n0034_inst_lut2_98,
      O => tx_input_n0074_2_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_114 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_120,
      I1 => tx_input_Msub_n0034_inst_lut2_98,
      O => tx_input_n0074_2_XORG
    );
  tx_input_n0074_2_CYINIT_1017 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_119,
      O => tx_input_n0074_2_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_122_1018 : X_MUX2
    port map (
      IA => tx_input_CNT(4),
      IB => tx_input_n0074_4_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_99,
      O => tx_input_Msub_n0034_inst_cy_122
    );
  tx_input_Msub_n0034_inst_sum_115 : X_XOR2
    port map (
      I0 => tx_input_n0074_4_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_99,
      O => tx_input_n0074_4_XORF
    );
  tx_input_Msub_n0034_inst_lut2_991 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_99
    );
  tx_input_Msub_n0034_inst_lut2_1001 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_100
    );
  tx_input_n0074_4_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_4_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_123
    );
  tx_input_n0074_4_XUSED : X_BUF
    port map (
      I => tx_input_n0074_4_XORF,
      O => tx_input_n0074(4)
    );
  tx_input_n0074_4_YUSED : X_BUF
    port map (
      I => tx_input_n0074_4_XORG,
      O => tx_input_n0074(5)
    );
  tx_input_Msub_n0034_inst_cy_123_1019 : X_MUX2
    port map (
      IA => tx_input_CNT(5),
      IB => tx_input_Msub_n0034_inst_cy_122,
      SEL => tx_input_Msub_n0034_inst_lut2_100,
      O => tx_input_n0074_4_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_116 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_122,
      I1 => tx_input_Msub_n0034_inst_lut2_100,
      O => tx_input_n0074_4_XORG
    );
  tx_input_n0074_4_CYINIT_1020 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_121,
      O => tx_input_n0074_4_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_124_1021 : X_MUX2
    port map (
      IA => tx_input_CNT(6),
      IB => tx_input_n0074_6_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_101,
      O => tx_input_Msub_n0034_inst_cy_124
    );
  tx_input_Msub_n0034_inst_sum_117 : X_XOR2
    port map (
      I0 => tx_input_n0074_6_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_101,
      O => tx_input_n0074_6_XORF
    );
  tx_input_Msub_n0034_inst_lut2_1011 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(6),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_101
    );
  tx_input_Msub_n0034_inst_lut2_1021 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(7),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_102
    );
  tx_input_n0074_6_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_6_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_125
    );
  tx_input_n0074_6_XUSED : X_BUF
    port map (
      I => tx_input_n0074_6_XORF,
      O => tx_input_n0074(6)
    );
  tx_input_n0074_6_YUSED : X_BUF
    port map (
      I => tx_input_n0074_6_XORG,
      O => tx_input_n0074(7)
    );
  tx_input_Msub_n0034_inst_cy_125_1022 : X_MUX2
    port map (
      IA => tx_input_CNT(7),
      IB => tx_input_Msub_n0034_inst_cy_124,
      SEL => tx_input_Msub_n0034_inst_lut2_102,
      O => tx_input_n0074_6_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_118 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_124,
      I1 => tx_input_Msub_n0034_inst_lut2_102,
      O => tx_input_n0074_6_XORG
    );
  tx_input_n0074_6_CYINIT_1023 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_123,
      O => tx_input_n0074_6_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_126_1024 : X_MUX2
    port map (
      IA => tx_input_CNT(8),
      IB => tx_input_n0074_8_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_103,
      O => tx_input_Msub_n0034_inst_cy_126
    );
  tx_input_Msub_n0034_inst_sum_119 : X_XOR2
    port map (
      I0 => tx_input_n0074_8_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_103,
      O => tx_input_n0074_8_XORF
    );
  tx_input_Msub_n0034_inst_lut2_1031 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_103
    );
  tx_input_Msub_n0034_inst_lut2_1041 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_104
    );
  tx_input_n0074_8_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_8_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_127
    );
  tx_input_n0074_8_XUSED : X_BUF
    port map (
      I => tx_input_n0074_8_XORF,
      O => tx_input_n0074(8)
    );
  tx_input_n0074_8_YUSED : X_BUF
    port map (
      I => tx_input_n0074_8_XORG,
      O => tx_input_n0074(9)
    );
  tx_input_Msub_n0034_inst_cy_127_1025 : X_MUX2
    port map (
      IA => tx_input_CNT(9),
      IB => tx_input_Msub_n0034_inst_cy_126,
      SEL => tx_input_Msub_n0034_inst_lut2_104,
      O => tx_input_n0074_8_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_120 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_126,
      I1 => tx_input_Msub_n0034_inst_lut2_104,
      O => tx_input_n0074_8_XORG
    );
  tx_input_n0074_8_CYINIT_1026 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_125,
      O => tx_input_n0074_8_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_128_1027 : X_MUX2
    port map (
      IA => tx_input_CNT(10),
      IB => tx_input_n0074_10_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_105,
      O => tx_input_Msub_n0034_inst_cy_128
    );
  tx_input_Msub_n0034_inst_sum_121 : X_XOR2
    port map (
      I0 => tx_input_n0074_10_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_105,
      O => tx_input_n0074_10_XORF
    );
  tx_input_Msub_n0034_inst_lut2_1051 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(10),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_105
    );
  tx_input_Msub_n0034_inst_lut2_1061 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(11),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_106
    );
  tx_input_n0074_10_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_10_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_129
    );
  tx_input_n0074_10_XUSED : X_BUF
    port map (
      I => tx_input_n0074_10_XORF,
      O => tx_input_n0074(10)
    );
  tx_input_n0074_10_YUSED : X_BUF
    port map (
      I => tx_input_n0074_10_XORG,
      O => tx_input_n0074(11)
    );
  tx_input_Msub_n0034_inst_cy_129_1028 : X_MUX2
    port map (
      IA => tx_input_CNT(11),
      IB => tx_input_Msub_n0034_inst_cy_128,
      SEL => tx_input_Msub_n0034_inst_lut2_106,
      O => tx_input_n0074_10_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_122 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_128,
      I1 => tx_input_Msub_n0034_inst_lut2_106,
      O => tx_input_n0074_10_XORG
    );
  tx_input_n0074_10_CYINIT_1029 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_127,
      O => tx_input_n0074_10_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_130_1030 : X_MUX2
    port map (
      IA => tx_input_CNT(12),
      IB => tx_input_n0074_12_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_107,
      O => tx_input_Msub_n0034_inst_cy_130
    );
  tx_input_Msub_n0034_inst_sum_123 : X_XOR2
    port map (
      I0 => tx_input_n0074_12_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_107,
      O => tx_input_n0074_12_XORF
    );
  tx_input_Msub_n0034_inst_lut2_1071 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(12),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_107
    );
  tx_input_Msub_n0034_inst_lut2_1081 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_108
    );
  tx_input_n0074_12_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_12_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_131
    );
  tx_input_n0074_12_XUSED : X_BUF
    port map (
      I => tx_input_n0074_12_XORF,
      O => tx_input_n0074(12)
    );
  tx_input_n0074_12_YUSED : X_BUF
    port map (
      I => tx_input_n0074_12_XORG,
      O => tx_input_n0074(13)
    );
  tx_input_Msub_n0034_inst_cy_131_1031 : X_MUX2
    port map (
      IA => tx_input_CNT(13),
      IB => tx_input_Msub_n0034_inst_cy_130,
      SEL => tx_input_Msub_n0034_inst_lut2_108,
      O => tx_input_n0074_12_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_124 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_130,
      I1 => tx_input_Msub_n0034_inst_lut2_108,
      O => tx_input_n0074_12_XORG
    );
  tx_input_n0074_12_CYINIT_1032 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_129,
      O => tx_input_n0074_12_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_132_1033 : X_MUX2
    port map (
      IA => tx_input_CNT(14),
      IB => tx_input_n0074_14_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_109,
      O => tx_input_Msub_n0034_inst_cy_132
    );
  tx_input_Msub_n0034_inst_sum_125 : X_XOR2
    port map (
      I0 => tx_input_n0074_14_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_109,
      O => tx_input_n0074_14_XORF
    );
  tx_input_Msub_n0034_inst_lut2_1091 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(14),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_109
    );
  tx_input_Msub_n0034_inst_lut2_1101 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(15),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_110
    );
  tx_input_n0074_14_XUSED : X_BUF
    port map (
      I => tx_input_n0074_14_XORF,
      O => tx_input_n0074(14)
    );
  tx_input_n0074_14_YUSED : X_BUF
    port map (
      I => tx_input_n0074_14_XORG,
      O => tx_input_n0074(15)
    );
  tx_input_Msub_n0034_inst_sum_126 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_132,
      I1 => tx_input_Msub_n0034_inst_lut2_110,
      O => tx_input_n0074_14_XORG
    );
  tx_input_n0074_14_CYINIT_1034 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_131,
      O => tx_input_n0074_14_CYINIT
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ONE_1035 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ZERO_1036 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_177_1037 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(32),
      ADR1 => rx_input_memio_addrchk_macaddrl(32),
      ADR2 => rx_input_memio_addrchk_datal(33),
      ADR3 => rx_input_memio_addrchk_macaddrl(33),
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(34),
      ADR1 => rx_input_memio_addrchk_datal(35),
      ADR2 => rx_input_memio_addrchk_macaddrl(35),
      ADR3 => rx_input_memio_addrchk_macaddrl(34),
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_1038 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_1_LOGIC_ZERO_1039 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_1_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_179_1040 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_1_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_1_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(37),
      ADR1 => rx_input_memio_addrchk_datal(36),
      ADR2 => rx_input_memio_addrchk_macaddrl(36),
      ADR3 => rx_input_memio_addrchk_macaddrl(37),
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(38),
      ADR1 => rx_input_memio_addrchk_datal(39),
      ADR2 => rx_input_memio_addrchk_macaddrl(39),
      ADR3 => rx_input_memio_addrchk_macaddrl(38),
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_1_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_1_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(1)
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_1_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_1_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_1_CYINIT_1041 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_1_CYINIT
    );
  mac_control_PHY_status_MII_Interface_mdccnt_32_LOGIC_ZERO_1042 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_mdccnt_32_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_187_1043 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_32,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_32_LOGIC_ZERO,
      SEL => mac_control_PHY_status_MII_Interface_cs_FFd5_rt,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_187
    );
  mac_control_PHY_status_MII_Interface_cs_FFd5_rt_1044 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_32,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_cs_FFd5_rt
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_341 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_17,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR2 => mac_control_PHY_status_MII_Interface_mdccnt_32,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_34
    );
  mac_control_PHY_status_MII_Interface_mdccnt_32_COUTUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_32_CYMUXG,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_188
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_188_1045 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_17,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_187,
      SEL => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_34,
      O => mac_control_PHY_status_MII_Interface_mdccnt_32_CYMUXG
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_165_1046 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_187,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_34,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_165
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_LOGIC_ZERO_1047 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_mdccnt_33_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_189_1048 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_mdccnt_33_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_33_CYINIT,
      SEL => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_35,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_189
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_166_1049 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_33_CYINIT,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_35,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_166
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_351 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => mac_control_PHY_status_MII_Interface_mdccnt_33,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_35
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_361 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR2 => mac_control_PHY_status_MII_Interface_mdccnt_34,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_36
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_COUTUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_33_CYMUXG,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_190
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_190_1050 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_mdccnt_33_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_189,
      SEL => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_36,
      O => mac_control_PHY_status_MII_Interface_mdccnt_33_CYMUXG
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_167_1051 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_189,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_36,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_167
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_CYINIT_1052 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_188,
      O => mac_control_PHY_status_MII_Interface_mdccnt_33_CYINIT
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_LOGIC_ZERO_1053 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_mdccnt_35_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_191_1054 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_mdccnt_35_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_35_CYINIT,
      SEL => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_37,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_191
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_168_1055 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_35_CYINIT,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_37,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_168
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_371 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_mdccnt_35,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_37
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_381 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR2 => mac_control_PHY_status_MII_Interface_mdccnt_36,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_38
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_COUTUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_35_CYMUXG,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_192
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_192_1056 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_mdccnt_35_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_191,
      SEL => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_38,
      O => mac_control_PHY_status_MII_Interface_mdccnt_35_CYMUXG
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_169_1057 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_191,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_38,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_169
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_CYINIT_1058 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_190,
      O => mac_control_PHY_status_MII_Interface_mdccnt_35_CYINIT
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_170_1059 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_37_CYINIT,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_39,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_170
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_391 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => mac_control_PHY_status_MII_Interface_mdccnt_37,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_39
    );
  mac_control_PHY_status_MII_Interface_n001124_SW0_2_1060 : X_LUT4
    generic map(
      INIT => X"FFAF"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_mdccnt_36,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_mdccnt_37,
      ADR3 => mac_control_PHY_status_MII_Interface_mdccnt_35,
      O => mac_control_PHY_status_MII_Interface_mdccnt_37_GROM
    );
  mac_control_PHY_status_MII_Interface_mdccnt_37_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_37_GROM,
      O => mac_control_PHY_status_MII_Interface_n001124_SW0_2
    );
  mac_control_PHY_status_MII_Interface_mdccnt_37_CYINIT_1061 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_192,
      O => mac_control_PHY_status_MII_Interface_mdccnt_37_CYINIT
    );
  rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ONE_1062 : X_ONE
    port map (
      O => rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ONE
    );
  rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ZERO_1063 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ZERO
    );
  rx_output_Mcompar_n0018_inst_cy_78_1064 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ONE,
      SEL => rx_output_Mcompar_n0018_inst_lut4_0,
      O => rx_output_Mcompar_n0018_inst_cy_78
    );
  rx_output_Mcompar_n0018_inst_lut4_01 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_output_bpl(0),
      ADR1 => addr3ext(0),
      ADR2 => addr3ext(1),
      ADR3 => rx_output_bpl(1),
      O => rx_output_Mcompar_n0018_inst_lut4_0
    );
  rx_output_Mcompar_n0018_inst_lut4_11 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_output_bpl(2),
      ADR1 => addr3ext(2),
      ADR2 => addr3ext(3),
      ADR3 => rx_output_bpl(3),
      O => rx_output_Mcompar_n0018_inst_lut4_1
    );
  rx_output_Mcompar_n0018_inst_cy_79_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_79_CYMUXG,
      O => rx_output_Mcompar_n0018_inst_cy_79
    );
  rx_output_Mcompar_n0018_inst_cy_79_1065 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_78,
      SEL => rx_output_Mcompar_n0018_inst_lut4_1,
      O => rx_output_Mcompar_n0018_inst_cy_79_CYMUXG
    );
  rx_output_Mcompar_n0018_inst_cy_81_LOGIC_ZERO_1066 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0018_inst_cy_81_LOGIC_ZERO
    );
  rx_output_Mcompar_n0018_inst_cy_80_1067 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_81_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_81_CYINIT,
      SEL => rx_output_Mcompar_n0018_inst_lut4_2,
      O => rx_output_Mcompar_n0018_inst_cy_80
    );
  rx_output_Mcompar_n0018_inst_lut4_21 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_output_bpl(5),
      ADR1 => rx_output_bpl(4),
      ADR2 => addr3ext(5),
      ADR3 => addr3ext(4),
      O => rx_output_Mcompar_n0018_inst_lut4_2
    );
  rx_output_Mcompar_n0018_inst_lut4_31 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_output_bpl(7),
      ADR1 => rx_output_bpl(6),
      ADR2 => addr3ext(7),
      ADR3 => addr3ext(6),
      O => rx_output_Mcompar_n0018_inst_lut4_3
    );
  rx_output_Mcompar_n0018_inst_cy_81_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_81_CYMUXG,
      O => rx_output_Mcompar_n0018_inst_cy_81
    );
  rx_output_Mcompar_n0018_inst_cy_81_1068 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_81_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_80,
      SEL => rx_output_Mcompar_n0018_inst_lut4_3,
      O => rx_output_Mcompar_n0018_inst_cy_81_CYMUXG
    );
  rx_output_Mcompar_n0018_inst_cy_81_CYINIT_1069 : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_79,
      O => rx_output_Mcompar_n0018_inst_cy_81_CYINIT
    );
  rx_output_Mcompar_n0018_inst_cy_83_LOGIC_ZERO_1070 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0018_inst_cy_83_LOGIC_ZERO
    );
  rx_output_Mcompar_n0018_inst_cy_82_1071 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_83_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_83_CYINIT,
      SEL => rx_output_Mcompar_n0018_inst_lut4_4,
      O => rx_output_Mcompar_n0018_inst_cy_82
    );
  rx_output_Mcompar_n0018_inst_lut4_41 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_output_bpl(8),
      ADR1 => addr3ext(9),
      ADR2 => addr3ext(8),
      ADR3 => rx_output_bpl(9),
      O => rx_output_Mcompar_n0018_inst_lut4_4
    );
  rx_output_Mcompar_n0018_inst_lut4_51 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_output_bpl(11),
      ADR1 => addr3ext(11),
      ADR2 => rx_output_bpl(10),
      ADR3 => addr3ext(10),
      O => rx_output_Mcompar_n0018_inst_lut4_5
    );
  rx_output_Mcompar_n0018_inst_cy_83_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_83_CYMUXG,
      O => rx_output_Mcompar_n0018_inst_cy_83
    );
  rx_output_Mcompar_n0018_inst_cy_83_1072 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_83_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_82,
      SEL => rx_output_Mcompar_n0018_inst_lut4_5,
      O => rx_output_Mcompar_n0018_inst_cy_83_CYMUXG
    );
  rx_output_Mcompar_n0018_inst_cy_83_CYINIT_1073 : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_81,
      O => rx_output_Mcompar_n0018_inst_cy_83_CYINIT
    );
  rx_output_n0018_LOGIC_ZERO_1074 : X_ZERO
    port map (
      O => rx_output_n0018_LOGIC_ZERO
    );
  rx_output_Mcompar_n0018_inst_cy_84_1075 : X_MUX2
    port map (
      IA => rx_output_n0018_LOGIC_ZERO,
      IB => rx_output_n0018_CYINIT,
      SEL => rx_output_Mcompar_n0018_inst_lut4_6,
      O => rx_output_Mcompar_n0018_inst_cy_84
    );
  rx_output_Mcompar_n0018_inst_lut4_61 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => addr3ext(13),
      ADR1 => rx_output_bpl(12),
      ADR2 => rx_output_bpl(13),
      ADR3 => addr3ext(12),
      O => rx_output_Mcompar_n0018_inst_lut4_6
    );
  rx_output_Mcompar_n0018_inst_lut4_71 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_output_bpl(15),
      ADR1 => addr3ext(15),
      ADR2 => addr3ext(14),
      ADR3 => rx_output_bpl(14),
      O => rx_output_Mcompar_n0018_inst_lut4_7
    );
  rx_output_n0018_COUTUSED : X_BUF
    port map (
      I => rx_output_n0018_CYMUXG,
      O => rx_output_n0018
    );
  rx_output_Mcompar_n0018_inst_cy_85 : X_MUX2
    port map (
      IA => rx_output_n0018_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_84,
      SEL => rx_output_Mcompar_n0018_inst_lut4_7,
      O => rx_output_n0018_CYMUXG
    );
  rx_output_n0018_CYINIT_1076 : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_83,
      O => rx_output_n0018_CYINIT
    );
  mac_control_txf_cnt_0_LOGIC_ZERO_1077 : X_ZERO
    port map (
      O => mac_control_txf_cnt_0_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_16_1078 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_0,
      IB => mac_control_txf_cnt_0_LOGIC_ZERO,
      SEL => mac_control_txf_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_txf_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_0,
      ADR1 => mac_control_txf_cnt(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_txf_cnt_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_56,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(1),
      O => mac_control_txf_cnt_0_GROM
    );
  mac_control_txf_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_0_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_17_1079 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_56,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_txf_cnt_0_GROM,
      O => mac_control_txf_cnt_0_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_txf_cnt_0_GROM,
      O => mac_control_txf_cnt_n0000(1)
    );
  mac_control_txf_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(3),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(3)
    );
  mac_control_txf_cnt_2_LOGIC_ZERO_1080 : X_ZERO
    port map (
      O => mac_control_txf_cnt_2_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_18_1081 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_2_LOGIC_ZERO,
      IB => mac_control_txf_cnt_2_CYINIT,
      SEL => mac_control_txf_cnt_2_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_2_CYINIT,
      I1 => mac_control_txf_cnt_2_FROM,
      O => mac_control_txf_cnt_n0000(2)
    );
  mac_control_txf_cnt_2_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_2_FROM
    );
  mac_control_txf_cnt_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(3),
      ADR3 => VCC,
      O => mac_control_txf_cnt_2_GROM
    );
  mac_control_txf_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_2_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_19_1082 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_2_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_txf_cnt_2_GROM,
      O => mac_control_txf_cnt_2_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_txf_cnt_2_GROM,
      O => mac_control_txf_cnt_n0000(3)
    );
  mac_control_txf_cnt_2_CYINIT_1083 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_txf_cnt_2_CYINIT
    );
  mac_control_txf_cnt_4_LOGIC_ZERO_1084 : X_ZERO
    port map (
      O => mac_control_txf_cnt_4_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_20_1085 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_4_LOGIC_ZERO,
      IB => mac_control_txf_cnt_4_CYINIT,
      SEL => mac_control_txf_cnt_4_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_4_CYINIT,
      I1 => mac_control_txf_cnt_4_FROM,
      O => mac_control_txf_cnt_n0000(4)
    );
  mac_control_txf_cnt_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_4_FROM
    );
  mac_control_txf_cnt_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(5),
      ADR3 => VCC,
      O => mac_control_txf_cnt_4_GROM
    );
  mac_control_txf_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_4_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_21_1086 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_4_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_txf_cnt_4_GROM,
      O => mac_control_txf_cnt_4_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_txf_cnt_4_GROM,
      O => mac_control_txf_cnt_n0000(5)
    );
  mac_control_txf_cnt_4_CYINIT_1087 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_txf_cnt_4_CYINIT
    );
  mac_control_txf_cnt_6_LOGIC_ZERO_1088 : X_ZERO
    port map (
      O => mac_control_txf_cnt_6_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_22_1089 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_6_LOGIC_ZERO,
      IB => mac_control_txf_cnt_6_CYINIT,
      SEL => mac_control_txf_cnt_6_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_6_CYINIT,
      I1 => mac_control_txf_cnt_6_FROM,
      O => mac_control_txf_cnt_n0000(6)
    );
  mac_control_txf_cnt_6_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txf_cnt(6),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_6_FROM
    );
  mac_control_txf_cnt_6_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(7),
      ADR3 => VCC,
      O => mac_control_txf_cnt_6_GROM
    );
  mac_control_txf_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_6_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_23_1090 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_6_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_txf_cnt_6_GROM,
      O => mac_control_txf_cnt_6_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_txf_cnt_6_GROM,
      O => mac_control_txf_cnt_n0000(7)
    );
  mac_control_txf_cnt_6_CYINIT_1091 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_txf_cnt_6_CYINIT
    );
  rx_input_fifo_control_dinl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(8),
      CE => rx_input_fifo_control_dinl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_9_FFY_RST,
      O => rx_input_fifo_control_dinl(8)
    );
  rx_input_fifo_control_dinl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_9_FFY_RST
    );
  mac_control_txf_cnt_8_LOGIC_ZERO_1092 : X_ZERO
    port map (
      O => mac_control_txf_cnt_8_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_24_1093 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_8_LOGIC_ZERO,
      IB => mac_control_txf_cnt_8_CYINIT,
      SEL => mac_control_txf_cnt_8_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_8_CYINIT,
      I1 => mac_control_txf_cnt_8_FROM,
      O => mac_control_txf_cnt_n0000(8)
    );
  mac_control_txf_cnt_8_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txf_cnt(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_8_FROM
    );
  mac_control_txf_cnt_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(9),
      ADR3 => VCC,
      O => mac_control_txf_cnt_8_GROM
    );
  mac_control_txf_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_8_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_25_1094 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_8_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_txf_cnt_8_GROM,
      O => mac_control_txf_cnt_8_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_txf_cnt_8_GROM,
      O => mac_control_txf_cnt_n0000(9)
    );
  mac_control_txf_cnt_8_CYINIT_1095 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_txf_cnt_8_CYINIT
    );
  mac_control_txf_cnt_10_LOGIC_ZERO_1096 : X_ZERO
    port map (
      O => mac_control_txf_cnt_10_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_26_1097 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_10_LOGIC_ZERO,
      IB => mac_control_txf_cnt_10_CYINIT,
      SEL => mac_control_txf_cnt_10_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_10_CYINIT,
      I1 => mac_control_txf_cnt_10_FROM,
      O => mac_control_txf_cnt_n0000(10)
    );
  mac_control_txf_cnt_10_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_10_FROM
    );
  mac_control_txf_cnt_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(11),
      ADR3 => VCC,
      O => mac_control_txf_cnt_10_GROM
    );
  mac_control_txf_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_10_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_27_1098 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_10_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_txf_cnt_10_GROM,
      O => mac_control_txf_cnt_10_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_txf_cnt_10_GROM,
      O => mac_control_txf_cnt_n0000(11)
    );
  mac_control_txf_cnt_10_CYINIT_1099 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_txf_cnt_10_CYINIT
    );
  mac_control_txf_cnt_12_LOGIC_ZERO_1100 : X_ZERO
    port map (
      O => mac_control_txf_cnt_12_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_28_1101 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_12_LOGIC_ZERO,
      IB => mac_control_txf_cnt_12_CYINIT,
      SEL => mac_control_txf_cnt_12_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_12_CYINIT,
      I1 => mac_control_txf_cnt_12_FROM,
      O => mac_control_txf_cnt_n0000(12)
    );
  mac_control_txf_cnt_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_12_FROM
    );
  mac_control_txf_cnt_12_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(13),
      ADR3 => VCC,
      O => mac_control_txf_cnt_12_GROM
    );
  mac_control_txf_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_12_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_29_1102 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_12_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_txf_cnt_12_GROM,
      O => mac_control_txf_cnt_12_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_txf_cnt_12_GROM,
      O => mac_control_txf_cnt_n0000(13)
    );
  mac_control_txf_cnt_12_CYINIT_1103 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_txf_cnt_12_CYINIT
    );
  mac_control_txf_cnt_14_LOGIC_ZERO_1104 : X_ZERO
    port map (
      O => mac_control_txf_cnt_14_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_30_1105 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_14_LOGIC_ZERO,
      IB => mac_control_txf_cnt_14_CYINIT,
      SEL => mac_control_txf_cnt_14_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_14_CYINIT,
      I1 => mac_control_txf_cnt_14_FROM,
      O => mac_control_txf_cnt_n0000(14)
    );
  mac_control_txf_cnt_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_14_FROM
    );
  mac_control_txf_cnt_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(15),
      ADR3 => VCC,
      O => mac_control_txf_cnt_14_GROM
    );
  mac_control_txf_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_14_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_31_1106 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_14_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_txf_cnt_14_GROM,
      O => mac_control_txf_cnt_14_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_txf_cnt_14_GROM,
      O => mac_control_txf_cnt_n0000(15)
    );
  mac_control_txf_cnt_14_CYINIT_1107 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_txf_cnt_14_CYINIT
    );
  mac_control_txf_cnt_16_LOGIC_ZERO_1108 : X_ZERO
    port map (
      O => mac_control_txf_cnt_16_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_32_1109 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_16_LOGIC_ZERO,
      IB => mac_control_txf_cnt_16_CYINIT,
      SEL => mac_control_txf_cnt_16_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_16_CYINIT,
      I1 => mac_control_txf_cnt_16_FROM,
      O => mac_control_txf_cnt_n0000(16)
    );
  mac_control_txf_cnt_16_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_16_FROM
    );
  mac_control_txf_cnt_16_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txf_cnt(17),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_16_GROM
    );
  mac_control_txf_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_16_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_33_1110 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_16_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_txf_cnt_16_GROM,
      O => mac_control_txf_cnt_16_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_txf_cnt_16_GROM,
      O => mac_control_txf_cnt_n0000(17)
    );
  mac_control_txf_cnt_16_CYINIT_1111 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_txf_cnt_16_CYINIT
    );
  rx_input_fifo_fifo_BU187 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2485,
      CE => rx_input_fifo_fifo_N2364,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2505_FFX_RST,
      O => rx_input_fifo_fifo_N2505
    );
  rx_input_fifo_fifo_N2505_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2505_FFX_RST
    );
  mac_control_txf_cnt_18_LOGIC_ZERO_1112 : X_ZERO
    port map (
      O => mac_control_txf_cnt_18_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_34_1113 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_18_LOGIC_ZERO,
      IB => mac_control_txf_cnt_18_CYINIT,
      SEL => mac_control_txf_cnt_18_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_18_CYINIT,
      I1 => mac_control_txf_cnt_18_FROM,
      O => mac_control_txf_cnt_n0000(18)
    );
  mac_control_txf_cnt_18_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txf_cnt(18),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_18_FROM
    );
  mac_control_txf_cnt_18_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txf_cnt(19),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_18_GROM
    );
  mac_control_txf_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_18_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_35_1114 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_18_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_txf_cnt_18_GROM,
      O => mac_control_txf_cnt_18_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_txf_cnt_18_GROM,
      O => mac_control_txf_cnt_n0000(19)
    );
  mac_control_txf_cnt_18_CYINIT_1115 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_txf_cnt_18_CYINIT
    );
  mac_control_txf_cnt_20_LOGIC_ZERO_1116 : X_ZERO
    port map (
      O => mac_control_txf_cnt_20_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_36_1117 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_20_LOGIC_ZERO,
      IB => mac_control_txf_cnt_20_CYINIT,
      SEL => mac_control_txf_cnt_20_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_20_CYINIT,
      I1 => mac_control_txf_cnt_20_FROM,
      O => mac_control_txf_cnt_n0000(20)
    );
  mac_control_txf_cnt_20_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(20),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_20_FROM
    );
  mac_control_txf_cnt_20_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txf_cnt(21),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_20_GROM
    );
  mac_control_txf_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_20_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_37_1118 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_20_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_txf_cnt_20_GROM,
      O => mac_control_txf_cnt_20_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_txf_cnt_20_GROM,
      O => mac_control_txf_cnt_n0000(21)
    );
  mac_control_txf_cnt_20_CYINIT_1119 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_txf_cnt_20_CYINIT
    );
  mac_control_txf_cnt_22_LOGIC_ZERO_1120 : X_ZERO
    port map (
      O => mac_control_txf_cnt_22_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_38_1121 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_22_LOGIC_ZERO,
      IB => mac_control_txf_cnt_22_CYINIT,
      SEL => mac_control_txf_cnt_22_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_22_CYINIT,
      I1 => mac_control_txf_cnt_22_FROM,
      O => mac_control_txf_cnt_n0000(22)
    );
  mac_control_txf_cnt_22_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txf_cnt(22),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_22_FROM
    );
  mac_control_txf_cnt_22_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(23),
      ADR3 => VCC,
      O => mac_control_txf_cnt_22_GROM
    );
  mac_control_txf_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_22_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_39_1122 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_22_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_txf_cnt_22_GROM,
      O => mac_control_txf_cnt_22_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_txf_cnt_22_GROM,
      O => mac_control_txf_cnt_n0000(23)
    );
  mac_control_txf_cnt_22_CYINIT_1123 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_txf_cnt_22_CYINIT
    );
  mac_control_txf_cnt_24_LOGIC_ZERO_1124 : X_ZERO
    port map (
      O => mac_control_txf_cnt_24_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_40_1125 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_24_LOGIC_ZERO,
      IB => mac_control_txf_cnt_24_CYINIT,
      SEL => mac_control_txf_cnt_24_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_24_CYINIT,
      I1 => mac_control_txf_cnt_24_FROM,
      O => mac_control_txf_cnt_n0000(24)
    );
  mac_control_txf_cnt_24_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(24),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_24_FROM
    );
  mac_control_txf_cnt_24_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txf_cnt(25),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_24_GROM
    );
  mac_control_txf_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_24_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_41_1126 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_24_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_txf_cnt_24_GROM,
      O => mac_control_txf_cnt_24_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_txf_cnt_24_GROM,
      O => mac_control_txf_cnt_n0000(25)
    );
  mac_control_txf_cnt_24_CYINIT_1127 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_txf_cnt_24_CYINIT
    );
  mac_control_txf_cnt_26_LOGIC_ZERO_1128 : X_ZERO
    port map (
      O => mac_control_txf_cnt_26_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_42_1129 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_26_LOGIC_ZERO,
      IB => mac_control_txf_cnt_26_CYINIT,
      SEL => mac_control_txf_cnt_26_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_26_CYINIT,
      I1 => mac_control_txf_cnt_26_FROM,
      O => mac_control_txf_cnt_n0000(26)
    );
  mac_control_txf_cnt_26_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(26),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_26_FROM
    );
  mac_control_txf_cnt_26_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(27),
      ADR3 => VCC,
      O => mac_control_txf_cnt_26_GROM
    );
  mac_control_txf_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_26_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_43_1130 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_26_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_txf_cnt_26_GROM,
      O => mac_control_txf_cnt_26_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_txf_cnt_26_GROM,
      O => mac_control_txf_cnt_n0000(27)
    );
  mac_control_txf_cnt_26_CYINIT_1131 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_txf_cnt_26_CYINIT
    );
  mac_control_txf_cnt_28_LOGIC_ZERO_1132 : X_ZERO
    port map (
      O => mac_control_txf_cnt_28_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_44_1133 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_28_LOGIC_ZERO,
      IB => mac_control_txf_cnt_28_CYINIT,
      SEL => mac_control_txf_cnt_28_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_28_CYINIT,
      I1 => mac_control_txf_cnt_28_FROM,
      O => mac_control_txf_cnt_n0000(28)
    );
  mac_control_txf_cnt_28_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(28),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_28_FROM
    );
  mac_control_txf_cnt_28_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(29),
      ADR3 => VCC,
      O => mac_control_txf_cnt_28_GROM
    );
  mac_control_txf_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_28_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_45_1134 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_28_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_txf_cnt_28_GROM,
      O => mac_control_txf_cnt_28_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_txf_cnt_28_GROM,
      O => mac_control_txf_cnt_n0000(29)
    );
  mac_control_txf_cnt_28_CYINIT_1135 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_txf_cnt_28_CYINIT
    );
  mac_control_txf_cnt_30_LOGIC_ZERO_1136 : X_ZERO
    port map (
      O => mac_control_txf_cnt_30_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_46_1137 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_30_LOGIC_ZERO,
      IB => mac_control_txf_cnt_30_CYINIT,
      SEL => mac_control_txf_cnt_30_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_30_CYINIT,
      I1 => mac_control_txf_cnt_30_FROM,
      O => mac_control_txf_cnt_n0000(30)
    );
  mac_control_txf_cnt_30_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(30),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_30_FROM
    );
  mac_control_txf_cnt_31_rt_1138 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(31),
      ADR3 => VCC,
      O => mac_control_txf_cnt_31_rt
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_txf_cnt_31_rt,
      O => mac_control_txf_cnt_n0000(31)
    );
  mac_control_txf_cnt_30_CYINIT_1139 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_txf_cnt_30_CYINIT
    );
  addr3ext_0_LOGIC_ZERO_1140 : X_ZERO
    port map (
      O => addr3ext_0_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_101_1141 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_15,
      IB => addr3ext_0_LOGIC_ZERO,
      SEL => rx_output_cs_FFd19_rt,
      O => rx_output_macnt_inst_cy_101
    );
  rx_output_cs_FFd19_rt_1142 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_15,
      ADR1 => rx_output_cs_FFd19,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_cs_FFd19_rt
    );
  rx_output_macnt_inst_lut3_01 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_39,
      ADR1 => rx_output_bp(0),
      ADR2 => addr3ext(0),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_0
    );
  addr3ext_0_COUTUSED : X_BUF
    port map (
      I => addr3ext_0_CYMUXG,
      O => rx_output_macnt_inst_cy_102
    );
  rx_output_macnt_inst_cy_102_1143 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_39,
      IB => rx_output_macnt_inst_cy_101,
      SEL => rx_output_macnt_inst_lut3_0,
      O => addr3ext_0_CYMUXG
    );
  rx_output_macnt_inst_sum_95_1144 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_101,
      I1 => rx_output_macnt_inst_lut3_0,
      O => rx_output_macnt_inst_sum_95
    );
  addr3ext_1_LOGIC_ZERO_1145 : X_ZERO
    port map (
      O => addr3ext_1_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_103_1146 : X_MUX2
    port map (
      IA => addr3ext_1_LOGIC_ZERO,
      IB => addr3ext_1_CYINIT,
      SEL => rx_output_macnt_inst_lut3_1,
      O => rx_output_macnt_inst_cy_103
    );
  rx_output_macnt_inst_sum_96_1147 : X_XOR2
    port map (
      I0 => addr3ext_1_CYINIT,
      I1 => rx_output_macnt_inst_lut3_1,
      O => rx_output_macnt_inst_sum_96
    );
  rx_output_macnt_inst_lut3_16 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(1),
      ADR2 => rx_output_bp(1),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_1
    );
  rx_output_macnt_inst_lut3_21 : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => rx_output_bp(2),
      ADR1 => addr3ext(2),
      ADR2 => VCC,
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_2
    );
  addr3ext_1_COUTUSED : X_BUF
    port map (
      I => addr3ext_1_CYMUXG,
      O => rx_output_macnt_inst_cy_104
    );
  rx_output_macnt_inst_cy_104_1148 : X_MUX2
    port map (
      IA => addr3ext_1_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_103,
      SEL => rx_output_macnt_inst_lut3_2,
      O => addr3ext_1_CYMUXG
    );
  rx_output_macnt_inst_sum_97_1149 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_103,
      I1 => rx_output_macnt_inst_lut3_2,
      O => rx_output_macnt_inst_sum_97
    );
  addr3ext_1_CYINIT_1150 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_102,
      O => addr3ext_1_CYINIT
    );
  addr3ext_3_LOGIC_ZERO_1151 : X_ZERO
    port map (
      O => addr3ext_3_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_105_1152 : X_MUX2
    port map (
      IA => addr3ext_3_LOGIC_ZERO,
      IB => addr3ext_3_CYINIT,
      SEL => rx_output_macnt_inst_lut3_3,
      O => rx_output_macnt_inst_cy_105
    );
  rx_output_macnt_inst_sum_98_1153 : X_XOR2
    port map (
      I0 => addr3ext_3_CYINIT,
      I1 => rx_output_macnt_inst_lut3_3,
      O => rx_output_macnt_inst_sum_98
    );
  rx_output_macnt_inst_lut3_31 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => VCC,
      ADR2 => rx_output_bp(3),
      ADR3 => addr3ext(3),
      O => rx_output_macnt_inst_lut3_3
    );
  rx_output_macnt_inst_lut3_41 : X_LUT4
    generic map(
      INIT => X"D8D8"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => rx_output_bp(4),
      ADR2 => addr3ext(4),
      ADR3 => VCC,
      O => rx_output_macnt_inst_lut3_4
    );
  addr3ext_3_COUTUSED : X_BUF
    port map (
      I => addr3ext_3_CYMUXG,
      O => rx_output_macnt_inst_cy_106
    );
  rx_output_macnt_inst_cy_106_1154 : X_MUX2
    port map (
      IA => addr3ext_3_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_105,
      SEL => rx_output_macnt_inst_lut3_4,
      O => addr3ext_3_CYMUXG
    );
  rx_output_macnt_inst_sum_99_1155 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_105,
      I1 => rx_output_macnt_inst_lut3_4,
      O => rx_output_macnt_inst_sum_99
    );
  addr3ext_3_CYINIT_1156 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_104,
      O => addr3ext_3_CYINIT
    );
  addr3ext_5_LOGIC_ZERO_1157 : X_ZERO
    port map (
      O => addr3ext_5_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_107_1158 : X_MUX2
    port map (
      IA => addr3ext_5_LOGIC_ZERO,
      IB => addr3ext_5_CYINIT,
      SEL => rx_output_macnt_inst_lut3_5,
      O => rx_output_macnt_inst_cy_107
    );
  rx_output_macnt_inst_sum_100_1159 : X_XOR2
    port map (
      I0 => addr3ext_5_CYINIT,
      I1 => rx_output_macnt_inst_lut3_5,
      O => rx_output_macnt_inst_sum_100
    );
  rx_output_macnt_inst_lut3_51 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => VCC,
      ADR2 => rx_output_bp(5),
      ADR3 => addr3ext(5),
      O => rx_output_macnt_inst_lut3_5
    );
  rx_output_macnt_inst_lut3_61 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(6),
      ADR2 => rx_output_bp(6),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_6
    );
  addr3ext_5_COUTUSED : X_BUF
    port map (
      I => addr3ext_5_CYMUXG,
      O => rx_output_macnt_inst_cy_108
    );
  rx_output_macnt_inst_cy_108_1160 : X_MUX2
    port map (
      IA => addr3ext_5_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_107,
      SEL => rx_output_macnt_inst_lut3_6,
      O => addr3ext_5_CYMUXG
    );
  rx_output_macnt_inst_sum_101_1161 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_107,
      I1 => rx_output_macnt_inst_lut3_6,
      O => rx_output_macnt_inst_sum_101
    );
  addr3ext_5_CYINIT_1162 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_106,
      O => addr3ext_5_CYINIT
    );
  addr3ext_7_LOGIC_ZERO_1163 : X_ZERO
    port map (
      O => addr3ext_7_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_109_1164 : X_MUX2
    port map (
      IA => addr3ext_7_LOGIC_ZERO,
      IB => addr3ext_7_CYINIT,
      SEL => rx_output_macnt_inst_lut3_7,
      O => rx_output_macnt_inst_cy_109
    );
  rx_output_macnt_inst_sum_102_1165 : X_XOR2
    port map (
      I0 => addr3ext_7_CYINIT,
      I1 => rx_output_macnt_inst_lut3_7,
      O => rx_output_macnt_inst_sum_102
    );
  rx_output_macnt_inst_lut3_71 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => addr3ext(7),
      ADR1 => rx_output_bp(7),
      ADR2 => VCC,
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_7
    );
  rx_output_macnt_inst_lut3_81 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => addr3ext(8),
      ADR2 => rx_output_bp(8),
      ADR3 => VCC,
      O => rx_output_macnt_inst_lut3_8
    );
  addr3ext_7_COUTUSED : X_BUF
    port map (
      I => addr3ext_7_CYMUXG,
      O => rx_output_macnt_inst_cy_110
    );
  rx_output_macnt_inst_cy_110_1166 : X_MUX2
    port map (
      IA => addr3ext_7_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_109,
      SEL => rx_output_macnt_inst_lut3_8,
      O => addr3ext_7_CYMUXG
    );
  rx_output_macnt_inst_sum_103_1167 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_109,
      I1 => rx_output_macnt_inst_lut3_8,
      O => rx_output_macnt_inst_sum_103
    );
  addr3ext_7_CYINIT_1168 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_108,
      O => addr3ext_7_CYINIT
    );
  addr3ext_9_LOGIC_ZERO_1169 : X_ZERO
    port map (
      O => addr3ext_9_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_111_1170 : X_MUX2
    port map (
      IA => addr3ext_9_LOGIC_ZERO,
      IB => addr3ext_9_CYINIT,
      SEL => rx_output_macnt_inst_lut3_9,
      O => rx_output_macnt_inst_cy_111
    );
  rx_output_macnt_inst_sum_104_1171 : X_XOR2
    port map (
      I0 => addr3ext_9_CYINIT,
      I1 => rx_output_macnt_inst_lut3_9,
      O => rx_output_macnt_inst_sum_104
    );
  rx_output_macnt_inst_lut3_91 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => addr3ext(9),
      ADR1 => rx_output_cs_FFd19,
      ADR2 => rx_output_bp(9),
      ADR3 => VCC,
      O => rx_output_macnt_inst_lut3_9
    );
  rx_output_macnt_inst_lut3_101 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_output_bp(10),
      ADR1 => VCC,
      ADR2 => addr3ext(10),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_10
    );
  addr3ext_9_COUTUSED : X_BUF
    port map (
      I => addr3ext_9_CYMUXG,
      O => rx_output_macnt_inst_cy_112
    );
  rx_output_macnt_inst_cy_112_1172 : X_MUX2
    port map (
      IA => addr3ext_9_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_111,
      SEL => rx_output_macnt_inst_lut3_10,
      O => addr3ext_9_CYMUXG
    );
  rx_output_macnt_inst_sum_105_1173 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_111,
      I1 => rx_output_macnt_inst_lut3_10,
      O => rx_output_macnt_inst_sum_105
    );
  addr3ext_9_CYINIT_1174 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_110,
      O => addr3ext_9_CYINIT
    );
  addr3ext_11_LOGIC_ZERO_1175 : X_ZERO
    port map (
      O => addr3ext_11_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_113_1176 : X_MUX2
    port map (
      IA => addr3ext_11_LOGIC_ZERO,
      IB => addr3ext_11_CYINIT,
      SEL => rx_output_macnt_inst_lut3_11,
      O => rx_output_macnt_inst_cy_113
    );
  rx_output_macnt_inst_sum_106_1177 : X_XOR2
    port map (
      I0 => addr3ext_11_CYINIT,
      I1 => rx_output_macnt_inst_lut3_11,
      O => rx_output_macnt_inst_sum_106
    );
  rx_output_macnt_inst_lut3_111 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => addr3ext(11),
      ADR1 => rx_output_cs_FFd19,
      ADR2 => rx_output_bp(11),
      ADR3 => VCC,
      O => rx_output_macnt_inst_lut3_11
    );
  rx_output_macnt_inst_lut3_121 : X_LUT4
    generic map(
      INIT => X"D8D8"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => rx_output_bp(12),
      ADR2 => addr3ext(12),
      ADR3 => VCC,
      O => rx_output_macnt_inst_lut3_12
    );
  addr3ext_11_COUTUSED : X_BUF
    port map (
      I => addr3ext_11_CYMUXG,
      O => rx_output_macnt_inst_cy_114
    );
  rx_output_macnt_inst_cy_114_1178 : X_MUX2
    port map (
      IA => addr3ext_11_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_113,
      SEL => rx_output_macnt_inst_lut3_12,
      O => addr3ext_11_CYMUXG
    );
  rx_output_macnt_inst_sum_107_1179 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_113,
      I1 => rx_output_macnt_inst_lut3_12,
      O => rx_output_macnt_inst_sum_107
    );
  addr3ext_11_CYINIT_1180 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_112,
      O => addr3ext_11_CYINIT
    );
  addr3ext_13_LOGIC_ZERO_1181 : X_ZERO
    port map (
      O => addr3ext_13_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_115_1182 : X_MUX2
    port map (
      IA => addr3ext_13_LOGIC_ZERO,
      IB => addr3ext_13_CYINIT,
      SEL => rx_output_macnt_inst_lut3_13,
      O => rx_output_macnt_inst_cy_115
    );
  rx_output_macnt_inst_sum_108_1183 : X_XOR2
    port map (
      I0 => addr3ext_13_CYINIT,
      I1 => rx_output_macnt_inst_lut3_13,
      O => rx_output_macnt_inst_sum_108
    );
  rx_output_macnt_inst_lut3_131 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(13),
      ADR2 => rx_output_bp(13),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_13
    );
  rx_output_macnt_inst_lut3_141 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => addr3ext(14),
      ADR1 => rx_output_cs_FFd19,
      ADR2 => rx_output_bp(14),
      ADR3 => VCC,
      O => rx_output_macnt_inst_lut3_14
    );
  addr3ext_13_COUTUSED : X_BUF
    port map (
      I => addr3ext_13_CYMUXG,
      O => rx_output_macnt_inst_cy_116
    );
  rx_output_macnt_inst_cy_116_1184 : X_MUX2
    port map (
      IA => addr3ext_13_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_115,
      SEL => rx_output_macnt_inst_lut3_14,
      O => addr3ext_13_CYMUXG
    );
  rx_output_macnt_inst_sum_109_1185 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_115,
      I1 => rx_output_macnt_inst_lut3_14,
      O => rx_output_macnt_inst_sum_109
    );
  addr3ext_13_CYINIT_1186 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_114,
      O => addr3ext_13_CYINIT
    );
  rx_output_macnt_inst_sum_110_1187 : X_XOR2
    port map (
      I0 => addr3ext_15_CYINIT,
      I1 => rx_output_macnt_inst_lut3_15,
      O => rx_output_macnt_inst_sum_110
    );
  rx_output_macnt_inst_lut3_151 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => addr3ext(15),
      ADR2 => rx_output_bp(15),
      ADR3 => VCC,
      O => rx_output_macnt_inst_lut3_15
    );
  rx_output_cs_FFd18_In_2_1188 : X_LUT4
    generic map(
      INIT => X"F5FF"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => VCC,
      ADR2 => rx_output_nfl,
      ADR3 => rx_output_nf,
      O => addr3ext_15_GROM
    );
  addr3ext_15_YUSED : X_BUF
    port map (
      I => addr3ext_15_GROM,
      O => rx_output_cs_FFd18_In_2
    );
  addr3ext_15_CYINIT_1189 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_116,
      O => addr3ext_15_CYINIT
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE_1190 : X_ONE
    port map (
      O => rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO_1191 : X_ZERO
    port map (
      O => rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_151_1192 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE,
      SEL => rx_fifocheck_diff_0_rt,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_151
    );
  rx_fifocheck_diff_0_rt_1193 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_fifocheck_diff(0),
      ADR3 => VCC,
      O => rx_fifocheck_diff_0_rt
    );
  rx_fifocheck_BEL_2 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_fifocheck_diff(0),
      ADR3 => VCC,
      O => rx_fifocheck_SIG_27
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_152_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_152
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_152_1194 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_151,
      SEL => rx_fifocheck_SIG_27,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE_1195 : X_ONE
    port map (
      O => rx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_153_1196 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut4_8,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_153
    );
  rx_fifocheck_Mcompar_n0003_inst_lut4_81 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(4),
      ADR1 => rx_fifocheck_diff(2),
      ADR2 => rx_fifocheck_diff(3),
      ADR3 => rx_fifocheck_diff(1),
      O => rx_fifocheck_Mcompar_n0003_inst_lut4_8
    );
  rx_fifocheck_Mcompar_n0003_inst_lut4_91 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(2),
      ADR1 => rx_fifocheck_diff(1),
      ADR2 => rx_fifocheck_diff(4),
      ADR3 => rx_fifocheck_diff(3),
      O => rx_fifocheck_Mcompar_n0003_inst_lut4_9
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_154_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_154
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_154_1197 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_153,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut4_9,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT_1198 : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_152,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT
    );
  tx_input_dh_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(10),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_11_FFY_RST,
      O => tx_input_dh(10)
    );
  tx_input_dh_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_11_FFY_RST
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE_1199 : X_ONE
    port map (
      O => rx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_155_1200 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut4_10,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_155
    );
  rx_fifocheck_Mcompar_n0003_inst_lut4_101 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(5),
      ADR1 => rx_fifocheck_diff(7),
      ADR2 => rx_fifocheck_diff(6),
      ADR3 => rx_fifocheck_diff(8),
      O => rx_fifocheck_Mcompar_n0003_inst_lut4_10
    );
  rx_fifocheck_Mcompar_n0003_inst_lut4_111 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(11),
      ADR1 => rx_fifocheck_diff(12),
      ADR2 => rx_fifocheck_diff(10),
      ADR3 => rx_fifocheck_diff(9),
      O => rx_fifocheck_Mcompar_n0003_inst_lut4_11
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_156_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_156
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_156_1201 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_155,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut4_11,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT_1202 : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_154,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO_1203 : X_ZERO
    port map (
      O => rx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_157_1204 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT,
      SEL => rx_fifocheck_diff_13_rt,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_157
    );
  rx_fifocheck_diff_13_rt_1205 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_fifocheck_diff(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_diff_13_rt
    );
  rx_fifocheck_BEL_3 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_fifocheck_diff(13),
      ADR3 => VCC,
      O => rx_fifocheck_SIG_28
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_158_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_158
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_158_1206 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_157,
      SEL => rx_fifocheck_SIG_28,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT_1207 : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_156,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT
    );
  rx_input_fifo_control_dinl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_dout(9),
      CE => rx_input_fifo_control_dinl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_9_FFX_RST,
      O => rx_input_fifo_control_dinl(9)
    );
  rx_input_fifo_control_dinl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_9_FFX_RST
    );
  rx_fifocheck_n0003_LOGIC_ONE_1208 : X_ONE
    port map (
      O => rx_fifocheck_n0003_LOGIC_ONE
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_159_1209 : X_MUX2
    port map (
      IA => rx_fifocheck_n0003_LOGIC_ONE,
      IB => rx_fifocheck_n0003_CYINIT,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut3_32,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_159
    );
  rx_fifocheck_Mcompar_n0003_inst_lut3_321 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => rx_fifocheck_diff(15),
      ADR1 => rx_fifocheck_diff(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_Mcompar_n0003_inst_lut3_32
    );
  rx_fifocheck_Mcompar_n0003_inst_lut3_331 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => rx_fifocheck_diff(15),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_diff(14),
      ADR3 => VCC,
      O => rx_fifocheck_Mcompar_n0003_inst_lut3_33
    );
  rx_fifocheck_n0003_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_n0003_CYMUXG,
      O => rx_fifocheck_n0003
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_160 : X_MUX2
    port map (
      IA => rx_fifocheck_n0003_LOGIC_ONE,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_159,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut3_33,
      O => rx_fifocheck_n0003_CYMUXG
    );
  rx_fifocheck_n0003_CYINIT_1210 : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_158,
      O => rx_fifocheck_n0003_CYINIT
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE_1211 : X_ONE
    port map (
      O => tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO_1212 : X_ZERO
    port map (
      O => tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_151_1213 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE,
      SEL => tx_fifocheck_diff_0_rt,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_151
    );
  tx_fifocheck_diff_0_rt_1214 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => tx_fifocheck_diff(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_diff_0_rt
    );
  tx_fifocheck_BEL_4 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_fifocheck_diff(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_SIG_29
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_152_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_152
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_152_1215 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_151,
      SEL => tx_fifocheck_SIG_29,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE_1216 : X_ONE
    port map (
      O => tx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_153_1217 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut4_8,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_153
    );
  tx_fifocheck_Mcompar_n0003_inst_lut4_81 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(2),
      ADR1 => tx_fifocheck_diff(3),
      ADR2 => tx_fifocheck_diff(1),
      ADR3 => tx_fifocheck_diff(4),
      O => tx_fifocheck_Mcompar_n0003_inst_lut4_8
    );
  tx_fifocheck_Mcompar_n0003_inst_lut4_91 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(2),
      ADR1 => tx_fifocheck_diff(3),
      ADR2 => tx_fifocheck_diff(1),
      ADR3 => tx_fifocheck_diff(4),
      O => tx_fifocheck_Mcompar_n0003_inst_lut4_9
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_154_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_154
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_154_1218 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_153,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut4_9,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT_1219 : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_152,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE_1220 : X_ONE
    port map (
      O => tx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_155_1221 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut4_10,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_155
    );
  tx_fifocheck_Mcompar_n0003_inst_lut4_101 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(8),
      ADR1 => tx_fifocheck_diff(5),
      ADR2 => tx_fifocheck_diff(7),
      ADR3 => tx_fifocheck_diff(6),
      O => tx_fifocheck_Mcompar_n0003_inst_lut4_10
    );
  tx_fifocheck_Mcompar_n0003_inst_lut4_111 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(11),
      ADR1 => tx_fifocheck_diff(10),
      ADR2 => tx_fifocheck_diff(12),
      ADR3 => tx_fifocheck_diff(9),
      O => tx_fifocheck_Mcompar_n0003_inst_lut4_11
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_156_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_156
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_156_1222 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_155,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut4_11,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT_1223 : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_154,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO_1224 : X_ZERO
    port map (
      O => tx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_157_1225 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT,
      SEL => tx_fifocheck_diff_13_rt,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_157
    );
  tx_fifocheck_diff_13_rt_1226 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_diff(13),
      O => tx_fifocheck_diff_13_rt
    );
  tx_fifocheck_BEL_5 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_diff(13),
      O => tx_fifocheck_SIG_30
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_158_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_158
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_158_1227 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_157,
      SEL => tx_fifocheck_SIG_30,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT_1228 : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_156,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT
    );
  tx_fifocheck_n0003_LOGIC_ONE_1229 : X_ONE
    port map (
      O => tx_fifocheck_n0003_LOGIC_ONE
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_159_1230 : X_MUX2
    port map (
      IA => tx_fifocheck_n0003_LOGIC_ONE,
      IB => tx_fifocheck_n0003_CYINIT,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut3_32,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_159
    );
  tx_fifocheck_Mcompar_n0003_inst_lut3_321 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => tx_fifocheck_diff(15),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_diff(14),
      O => tx_fifocheck_Mcompar_n0003_inst_lut3_32
    );
  tx_fifocheck_Mcompar_n0003_inst_lut3_331 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_fifocheck_diff(14),
      ADR3 => tx_fifocheck_diff(15),
      O => tx_fifocheck_Mcompar_n0003_inst_lut3_33
    );
  tx_fifocheck_n0003_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_n0003_CYMUXG,
      O => tx_fifocheck_n0003
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_160 : X_MUX2
    port map (
      IA => tx_fifocheck_n0003_LOGIC_ONE,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_159,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut3_33,
      O => tx_fifocheck_n0003_CYMUXG
    );
  tx_fifocheck_n0003_CYINIT_1231 : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_158,
      O => tx_fifocheck_n0003_CYINIT
    );
  mac_control_phyrstcnt_110_LOGIC_ONE_1232 : X_ONE
    port map (
      O => mac_control_phyrstcnt_110_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_294_1233 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_10,
      IB => mac_control_phyrstcnt_110_LOGIC_ONE,
      SEL => mac_control_N52153_rt,
      O => mac_control_phyrstcnt_inst_cy_294
    );
  mac_control_N52153_rt_1234 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_10,
      ADR1 => VCC,
      ADR2 => mac_control_N52153,
      ADR3 => VCC,
      O => mac_control_N52153_rt
    );
  mac_control_phyrstcnt_inst_lut3_1921 : X_LUT4
    generic map(
      INIT => X"FF0F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_35,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_110,
      ADR3 => mac_control_N52153,
      O => mac_control_phyrstcnt_inst_lut3_192
    );
  mac_control_phyrstcnt_110_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_110_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_295
    );
  mac_control_phyrstcnt_inst_cy_295_1235 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_35,
      IB => mac_control_phyrstcnt_inst_cy_294,
      SEL => mac_control_phyrstcnt_inst_lut3_192,
      O => mac_control_phyrstcnt_110_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_257_1236 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_294,
      I1 => mac_control_phyrstcnt_inst_lut3_192,
      O => mac_control_phyrstcnt_inst_sum_257
    );
  mac_control_phyrstcnt_111_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_111_FFY_RST
    );
  mac_control_phyrstcnt_112_1237 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_259,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_111_FFY_RST,
      O => mac_control_phyrstcnt_112
    );
  mac_control_phyrstcnt_111_LOGIC_ONE_1238 : X_ONE
    port map (
      O => mac_control_phyrstcnt_111_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_296_1239 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_111_LOGIC_ONE,
      IB => mac_control_phyrstcnt_111_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_193,
      O => mac_control_phyrstcnt_inst_cy_296
    );
  mac_control_phyrstcnt_inst_sum_258_1240 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_111_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_193,
      O => mac_control_phyrstcnt_inst_sum_258
    );
  mac_control_phyrstcnt_inst_lut3_1931 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_111,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_193
    );
  mac_control_phyrstcnt_inst_lut3_1941 : X_LUT4
    generic map(
      INIT => X"AAFF"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_112,
      O => mac_control_phyrstcnt_inst_lut3_194
    );
  mac_control_phyrstcnt_111_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_111_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_297
    );
  mac_control_phyrstcnt_inst_cy_297_1241 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_111_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_296,
      SEL => mac_control_phyrstcnt_inst_lut3_194,
      O => mac_control_phyrstcnt_111_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_259_1242 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_296,
      I1 => mac_control_phyrstcnt_inst_lut3_194,
      O => mac_control_phyrstcnt_inst_sum_259
    );
  mac_control_phyrstcnt_111_CYINIT_1243 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_295,
      O => mac_control_phyrstcnt_111_CYINIT
    );
  mac_control_phyrstcnt_113_LOGIC_ONE_1244 : X_ONE
    port map (
      O => mac_control_phyrstcnt_113_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_298_1245 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_113_LOGIC_ONE,
      IB => mac_control_phyrstcnt_113_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_195,
      O => mac_control_phyrstcnt_inst_cy_298
    );
  mac_control_phyrstcnt_inst_sum_260_1246 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_113_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_195,
      O => mac_control_phyrstcnt_inst_sum_260
    );
  mac_control_phyrstcnt_inst_lut3_1951 : X_LUT4
    generic map(
      INIT => X"BBBB"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => mac_control_phyrstcnt_113,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_195
    );
  mac_control_phyrstcnt_inst_lut3_1961 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_114,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_196
    );
  mac_control_phyrstcnt_113_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_113_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_299
    );
  mac_control_phyrstcnt_inst_cy_299_1247 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_113_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_298,
      SEL => mac_control_phyrstcnt_inst_lut3_196,
      O => mac_control_phyrstcnt_113_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_261_1248 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_298,
      I1 => mac_control_phyrstcnt_inst_lut3_196,
      O => mac_control_phyrstcnt_inst_sum_261
    );
  mac_control_phyrstcnt_113_CYINIT_1249 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_297,
      O => mac_control_phyrstcnt_113_CYINIT
    );
  mac_control_phyrstcnt_115_LOGIC_ONE_1250 : X_ONE
    port map (
      O => mac_control_phyrstcnt_115_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_300_1251 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_115_LOGIC_ONE,
      IB => mac_control_phyrstcnt_115_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_197,
      O => mac_control_phyrstcnt_inst_cy_300
    );
  mac_control_phyrstcnt_inst_sum_262_1252 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_115_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_197,
      O => mac_control_phyrstcnt_inst_sum_262
    );
  mac_control_phyrstcnt_inst_lut3_1971 : X_LUT4
    generic map(
      INIT => X"DDDD"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_115,
      ADR1 => mac_control_N52153,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_197
    );
  mac_control_phyrstcnt_inst_lut3_1981 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N52153,
      ADR2 => mac_control_phyrstcnt_116,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_198
    );
  mac_control_phyrstcnt_115_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_115_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_301
    );
  mac_control_phyrstcnt_inst_cy_301_1253 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_115_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_300,
      SEL => mac_control_phyrstcnt_inst_lut3_198,
      O => mac_control_phyrstcnt_115_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_263_1254 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_300,
      I1 => mac_control_phyrstcnt_inst_lut3_198,
      O => mac_control_phyrstcnt_inst_sum_263
    );
  mac_control_phyrstcnt_115_CYINIT_1255 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_299,
      O => mac_control_phyrstcnt_115_CYINIT
    );
  mac_control_phyrstcnt_117_LOGIC_ONE_1256 : X_ONE
    port map (
      O => mac_control_phyrstcnt_117_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_302_1257 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_117_LOGIC_ONE,
      IB => mac_control_phyrstcnt_117_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_199,
      O => mac_control_phyrstcnt_inst_cy_302
    );
  mac_control_phyrstcnt_inst_sum_264_1258 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_117_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_199,
      O => mac_control_phyrstcnt_inst_sum_264
    );
  mac_control_phyrstcnt_inst_lut3_1991 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyrstcnt_117,
      ADR2 => mac_control_N52153,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_199
    );
  mac_control_phyrstcnt_inst_lut3_2001 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_118,
      ADR1 => VCC,
      ADR2 => mac_control_N52153,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_200
    );
  mac_control_phyrstcnt_117_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_117_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_303
    );
  mac_control_phyrstcnt_inst_cy_303_1259 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_117_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_302,
      SEL => mac_control_phyrstcnt_inst_lut3_200,
      O => mac_control_phyrstcnt_117_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_265_1260 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_302,
      I1 => mac_control_phyrstcnt_inst_lut3_200,
      O => mac_control_phyrstcnt_inst_sum_265
    );
  mac_control_phyrstcnt_117_CYINIT_1261 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_301,
      O => mac_control_phyrstcnt_117_CYINIT
    );
  mac_control_phyrstcnt_119_LOGIC_ONE_1262 : X_ONE
    port map (
      O => mac_control_phyrstcnt_119_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_304_1263 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_119_LOGIC_ONE,
      IB => mac_control_phyrstcnt_119_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_201,
      O => mac_control_phyrstcnt_inst_cy_304
    );
  mac_control_phyrstcnt_inst_sum_266_1264 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_119_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_201,
      O => mac_control_phyrstcnt_inst_sum_266
    );
  mac_control_phyrstcnt_inst_lut3_2011 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyrstcnt_119,
      ADR2 => mac_control_N52153,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_201
    );
  mac_control_phyrstcnt_inst_lut3_2021 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_N52153,
      ADR3 => mac_control_phyrstcnt_120,
      O => mac_control_phyrstcnt_inst_lut3_202
    );
  mac_control_phyrstcnt_119_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_119_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_305
    );
  mac_control_phyrstcnt_inst_cy_305_1265 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_119_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_304,
      SEL => mac_control_phyrstcnt_inst_lut3_202,
      O => mac_control_phyrstcnt_119_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_267_1266 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_304,
      I1 => mac_control_phyrstcnt_inst_lut3_202,
      O => mac_control_phyrstcnt_inst_sum_267
    );
  mac_control_phyrstcnt_119_CYINIT_1267 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_303,
      O => mac_control_phyrstcnt_119_CYINIT
    );
  mac_control_phyrstcnt_121_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_121_FFX_RST
    );
  mac_control_phyrstcnt_121_1268 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_268,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_121_FFX_RST,
      O => mac_control_phyrstcnt_121
    );
  mac_control_phyrstcnt_121_LOGIC_ONE_1269 : X_ONE
    port map (
      O => mac_control_phyrstcnt_121_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_306_1270 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_121_LOGIC_ONE,
      IB => mac_control_phyrstcnt_121_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_203,
      O => mac_control_phyrstcnt_inst_cy_306
    );
  mac_control_phyrstcnt_inst_sum_268_1271 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_121_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_203,
      O => mac_control_phyrstcnt_inst_sum_268
    );
  mac_control_phyrstcnt_inst_lut3_2031 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_121,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_203
    );
  mac_control_phyrstcnt_inst_lut3_2041 : X_LUT4
    generic map(
      INIT => X"AAFF"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_122,
      O => mac_control_phyrstcnt_inst_lut3_204
    );
  mac_control_phyrstcnt_121_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_121_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_307
    );
  mac_control_phyrstcnt_inst_cy_307_1272 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_121_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_306,
      SEL => mac_control_phyrstcnt_inst_lut3_204,
      O => mac_control_phyrstcnt_121_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_269_1273 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_306,
      I1 => mac_control_phyrstcnt_inst_lut3_204,
      O => mac_control_phyrstcnt_inst_sum_269
    );
  mac_control_phyrstcnt_121_CYINIT_1274 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_305,
      O => mac_control_phyrstcnt_121_CYINIT
    );
  tx_input_dh_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(11),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_11_FFX_RST,
      O => tx_input_dh(11)
    );
  tx_input_dh_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_11_FFX_RST
    );
  mac_control_phyrstcnt_123_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_123_FFX_RST
    );
  mac_control_phyrstcnt_123_1275 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_270,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_123_FFX_RST,
      O => mac_control_phyrstcnt_123
    );
  mac_control_phyrstcnt_123_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_123_FFY_RST
    );
  mac_control_phyrstcnt_124_1276 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_271,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_123_FFY_RST,
      O => mac_control_phyrstcnt_124
    );
  mac_control_phyrstcnt_123_LOGIC_ONE_1277 : X_ONE
    port map (
      O => mac_control_phyrstcnt_123_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_308_1278 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_123_LOGIC_ONE,
      IB => mac_control_phyrstcnt_123_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_205,
      O => mac_control_phyrstcnt_inst_cy_308
    );
  mac_control_phyrstcnt_inst_sum_270_1279 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_123_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_205,
      O => mac_control_phyrstcnt_inst_sum_270
    );
  mac_control_phyrstcnt_inst_lut3_2051 : X_LUT4
    generic map(
      INIT => X"F5F5"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_123,
      ADR1 => VCC,
      ADR2 => mac_control_N52153,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_205
    );
  mac_control_phyrstcnt_inst_lut3_2061 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_124,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_206
    );
  mac_control_phyrstcnt_123_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_123_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_309
    );
  mac_control_phyrstcnt_inst_cy_309_1280 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_123_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_308,
      SEL => mac_control_phyrstcnt_inst_lut3_206,
      O => mac_control_phyrstcnt_123_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_271_1281 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_308,
      I1 => mac_control_phyrstcnt_inst_lut3_206,
      O => mac_control_phyrstcnt_inst_sum_271
    );
  mac_control_phyrstcnt_123_CYINIT_1282 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_307,
      O => mac_control_phyrstcnt_123_CYINIT
    );
  mac_control_phyrstcnt_125_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_125_FFX_RST
    );
  mac_control_phyrstcnt_125_1283 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_272,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_125_FFX_RST,
      O => mac_control_phyrstcnt_125
    );
  mac_control_phyrstcnt_125_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_125_FFY_RST
    );
  mac_control_phyrstcnt_126_1284 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_273,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_125_FFY_RST,
      O => mac_control_phyrstcnt_126
    );
  mac_control_phyrstcnt_125_LOGIC_ONE_1285 : X_ONE
    port map (
      O => mac_control_phyrstcnt_125_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_310_1286 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_125_LOGIC_ONE,
      IB => mac_control_phyrstcnt_125_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_207,
      O => mac_control_phyrstcnt_inst_cy_310
    );
  mac_control_phyrstcnt_inst_sum_272_1287 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_125_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_207,
      O => mac_control_phyrstcnt_inst_sum_272
    );
  mac_control_phyrstcnt_inst_lut3_2071 : X_LUT4
    generic map(
      INIT => X"CFCF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N52153,
      ADR2 => mac_control_phyrstcnt_125,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_207
    );
  mac_control_phyrstcnt_inst_lut3_2081 : X_LUT4
    generic map(
      INIT => X"AAFF"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_126,
      O => mac_control_phyrstcnt_inst_lut3_208
    );
  mac_control_phyrstcnt_125_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_125_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_311
    );
  mac_control_phyrstcnt_inst_cy_311_1288 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_125_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_310,
      SEL => mac_control_phyrstcnt_inst_lut3_208,
      O => mac_control_phyrstcnt_125_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_273_1289 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_310,
      I1 => mac_control_phyrstcnt_inst_lut3_208,
      O => mac_control_phyrstcnt_inst_sum_273
    );
  mac_control_phyrstcnt_125_CYINIT_1290 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_309,
      O => mac_control_phyrstcnt_125_CYINIT
    );
  mac_control_phyrstcnt_127_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_127_FFY_RST
    );
  mac_control_phyrstcnt_128_1291 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_275,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_127_FFY_RST,
      O => mac_control_phyrstcnt_128
    );
  mac_control_phyrstcnt_127_LOGIC_ONE_1292 : X_ONE
    port map (
      O => mac_control_phyrstcnt_127_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_312_1293 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_127_LOGIC_ONE,
      IB => mac_control_phyrstcnt_127_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_209,
      O => mac_control_phyrstcnt_inst_cy_312
    );
  mac_control_phyrstcnt_inst_sum_274_1294 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_127_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_209,
      O => mac_control_phyrstcnt_inst_sum_274
    );
  mac_control_phyrstcnt_inst_lut3_2091 : X_LUT4
    generic map(
      INIT => X"F5F5"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_127,
      ADR1 => VCC,
      ADR2 => mac_control_N52153,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_209
    );
  mac_control_phyrstcnt_inst_lut3_2101 : X_LUT4
    generic map(
      INIT => X"CCFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N52153,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_128,
      O => mac_control_phyrstcnt_inst_lut3_210
    );
  mac_control_phyrstcnt_127_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_127_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_313
    );
  mac_control_phyrstcnt_inst_cy_313_1295 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_127_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_312,
      SEL => mac_control_phyrstcnt_inst_lut3_210,
      O => mac_control_phyrstcnt_127_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_275_1296 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_312,
      I1 => mac_control_phyrstcnt_inst_lut3_210,
      O => mac_control_phyrstcnt_inst_sum_275
    );
  mac_control_phyrstcnt_127_CYINIT_1297 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_311,
      O => mac_control_phyrstcnt_127_CYINIT
    );
  mac_control_phyrstcnt_129_LOGIC_ONE_1298 : X_ONE
    port map (
      O => mac_control_phyrstcnt_129_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_314_1299 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_129_LOGIC_ONE,
      IB => mac_control_phyrstcnt_129_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_211,
      O => mac_control_phyrstcnt_inst_cy_314
    );
  mac_control_phyrstcnt_inst_sum_276_1300 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_129_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_211,
      O => mac_control_phyrstcnt_inst_sum_276
    );
  mac_control_phyrstcnt_inst_lut3_2111 : X_LUT4
    generic map(
      INIT => X"AAFF"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_129,
      O => mac_control_phyrstcnt_inst_lut3_211
    );
  mac_control_phyrstcnt_inst_lut3_2121 : X_LUT4
    generic map(
      INIT => X"AAFF"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_130,
      O => mac_control_phyrstcnt_inst_lut3_212
    );
  mac_control_phyrstcnt_129_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_129_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_315
    );
  mac_control_phyrstcnt_inst_cy_315_1301 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_129_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_314,
      SEL => mac_control_phyrstcnt_inst_lut3_212,
      O => mac_control_phyrstcnt_129_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_277_1302 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_314,
      I1 => mac_control_phyrstcnt_inst_lut3_212,
      O => mac_control_phyrstcnt_inst_sum_277
    );
  mac_control_phyrstcnt_129_CYINIT_1303 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_313,
      O => mac_control_phyrstcnt_129_CYINIT
    );
  mac_control_phyrstcnt_131_LOGIC_ONE_1304 : X_ONE
    port map (
      O => mac_control_phyrstcnt_131_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_316_1305 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_131_LOGIC_ONE,
      IB => mac_control_phyrstcnt_131_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_213,
      O => mac_control_phyrstcnt_inst_cy_316
    );
  mac_control_phyrstcnt_inst_sum_278_1306 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_131_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_213,
      O => mac_control_phyrstcnt_inst_sum_278
    );
  mac_control_phyrstcnt_inst_lut3_2131 : X_LUT4
    generic map(
      INIT => X"DDDD"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_131,
      ADR1 => mac_control_N52153,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_213
    );
  mac_control_phyrstcnt_inst_lut3_2141 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_132,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_214
    );
  mac_control_phyrstcnt_131_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_131_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_317
    );
  mac_control_phyrstcnt_inst_cy_317_1307 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_131_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_316,
      SEL => mac_control_phyrstcnt_inst_lut3_214,
      O => mac_control_phyrstcnt_131_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_279_1308 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_316,
      I1 => mac_control_phyrstcnt_inst_lut3_214,
      O => mac_control_phyrstcnt_inst_sum_279
    );
  mac_control_phyrstcnt_131_CYINIT_1309 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_315,
      O => mac_control_phyrstcnt_131_CYINIT
    );
  mac_control_phyrstcnt_133_LOGIC_ONE_1310 : X_ONE
    port map (
      O => mac_control_phyrstcnt_133_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_318_1311 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_133_LOGIC_ONE,
      IB => mac_control_phyrstcnt_133_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_215,
      O => mac_control_phyrstcnt_inst_cy_318
    );
  mac_control_phyrstcnt_inst_sum_280_1312 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_133_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_215,
      O => mac_control_phyrstcnt_inst_sum_280
    );
  mac_control_phyrstcnt_inst_lut3_2151 : X_LUT4
    generic map(
      INIT => X"DDDD"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_133,
      ADR1 => mac_control_N52153,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_215
    );
  mac_control_phyrstcnt_inst_lut3_2161 : X_LUT4
    generic map(
      INIT => X"CCFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N52153,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_134,
      O => mac_control_phyrstcnt_inst_lut3_216
    );
  mac_control_phyrstcnt_133_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_133_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_319
    );
  mac_control_phyrstcnt_inst_cy_319_1313 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_133_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_318,
      SEL => mac_control_phyrstcnt_inst_lut3_216,
      O => mac_control_phyrstcnt_133_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_281_1314 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_318,
      I1 => mac_control_phyrstcnt_inst_lut3_216,
      O => mac_control_phyrstcnt_inst_sum_281
    );
  mac_control_phyrstcnt_133_CYINIT_1315 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_317,
      O => mac_control_phyrstcnt_133_CYINIT
    );
  mac_control_phyrstcnt_135_LOGIC_ONE_1316 : X_ONE
    port map (
      O => mac_control_phyrstcnt_135_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_320_1317 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_135_LOGIC_ONE,
      IB => mac_control_phyrstcnt_135_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_217,
      O => mac_control_phyrstcnt_inst_cy_320
    );
  mac_control_phyrstcnt_inst_sum_282_1318 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_135_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_217,
      O => mac_control_phyrstcnt_inst_sum_282
    );
  mac_control_phyrstcnt_inst_lut3_2171 : X_LUT4
    generic map(
      INIT => X"FF55"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_135,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_N52153,
      O => mac_control_phyrstcnt_inst_lut3_217
    );
  mac_control_phyrstcnt_inst_lut3_2181 : X_LUT4
    generic map(
      INIT => X"AAFF"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_136,
      O => mac_control_phyrstcnt_inst_lut3_218
    );
  mac_control_phyrstcnt_135_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_135_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_321
    );
  mac_control_phyrstcnt_inst_cy_321_1319 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_135_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_320,
      SEL => mac_control_phyrstcnt_inst_lut3_218,
      O => mac_control_phyrstcnt_135_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_283_1320 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_320,
      I1 => mac_control_phyrstcnt_inst_lut3_218,
      O => mac_control_phyrstcnt_inst_sum_283
    );
  mac_control_phyrstcnt_135_CYINIT_1321 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_319,
      O => mac_control_phyrstcnt_135_CYINIT
    );
  mac_control_phyrstcnt_137_LOGIC_ONE_1322 : X_ONE
    port map (
      O => mac_control_phyrstcnt_137_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_322_1323 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_137_LOGIC_ONE,
      IB => mac_control_phyrstcnt_137_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_219,
      O => mac_control_phyrstcnt_inst_cy_322
    );
  mac_control_phyrstcnt_inst_sum_284_1324 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_137_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_219,
      O => mac_control_phyrstcnt_inst_sum_284
    );
  mac_control_phyrstcnt_inst_lut3_2191 : X_LUT4
    generic map(
      INIT => X"CFCF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N52153,
      ADR2 => mac_control_phyrstcnt_137,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_219
    );
  mac_control_phyrstcnt_inst_lut3_2201 : X_LUT4
    generic map(
      INIT => X"BBBB"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => mac_control_phyrstcnt_138,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_220
    );
  mac_control_phyrstcnt_137_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_137_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_323
    );
  mac_control_phyrstcnt_inst_cy_323_1325 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_137_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_322,
      SEL => mac_control_phyrstcnt_inst_lut3_220,
      O => mac_control_phyrstcnt_137_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_285_1326 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_322,
      I1 => mac_control_phyrstcnt_inst_lut3_220,
      O => mac_control_phyrstcnt_inst_sum_285
    );
  mac_control_phyrstcnt_137_CYINIT_1327 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_321,
      O => mac_control_phyrstcnt_137_CYINIT
    );
  mac_control_phyrstcnt_139_LOGIC_ONE_1328 : X_ONE
    port map (
      O => mac_control_phyrstcnt_139_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_324_1329 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_139_LOGIC_ONE,
      IB => mac_control_phyrstcnt_139_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_221,
      O => mac_control_phyrstcnt_inst_cy_324
    );
  mac_control_phyrstcnt_inst_sum_286_1330 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_139_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_221,
      O => mac_control_phyrstcnt_inst_sum_286
    );
  mac_control_phyrstcnt_inst_lut3_2211 : X_LUT4
    generic map(
      INIT => X"CCFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N52153,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_139,
      O => mac_control_phyrstcnt_inst_lut3_221
    );
  mac_control_phyrstcnt_inst_lut3_2221 : X_LUT4
    generic map(
      INIT => X"CCFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N52153,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_140,
      O => mac_control_phyrstcnt_inst_lut3_222
    );
  mac_control_phyrstcnt_139_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_139_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_325
    );
  mac_control_phyrstcnt_inst_cy_325_1331 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_139_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_324,
      SEL => mac_control_phyrstcnt_inst_lut3_222,
      O => mac_control_phyrstcnt_139_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_287_1332 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_324,
      I1 => mac_control_phyrstcnt_inst_lut3_222,
      O => mac_control_phyrstcnt_inst_sum_287
    );
  mac_control_phyrstcnt_139_CYINIT_1333 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_323,
      O => mac_control_phyrstcnt_139_CYINIT
    );
  mac_control_phyrstcnt_inst_sum_288_1334 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_141_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_223,
      O => mac_control_phyrstcnt_inst_sum_288
    );
  mac_control_phyrstcnt_inst_lut3_2231 : X_LUT4
    generic map(
      INIT => X"FF55"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_141,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_N52153,
      O => mac_control_phyrstcnt_inst_lut3_223
    );
  mac_control_phyrstcnt_141_CYINIT_1335 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_325,
      O => mac_control_phyrstcnt_141_CYINIT
    );
  rx_input_memio_macnt_70_LOGIC_ZERO_1336 : X_ZERO
    port map (
      O => rx_input_memio_macnt_70_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_253_1337 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_37,
      IB => rx_input_memio_macnt_70_LOGIC_ZERO,
      SEL => rx_input_memio_SIG_31,
      O => rx_input_memio_macnt_inst_cy_253
    );
  rx_input_memio_BEL_6 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_37,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_SIG_31
    );
  rx_input_memio_macnt_inst_lut3_561 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_1,
      ADR1 => rx_input_memio_bp(0),
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => rx_input_memio_macnt_70,
      O => rx_input_memio_macnt_inst_lut3_56
    );
  rx_input_memio_macnt_70_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_70_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_254
    );
  rx_input_memio_macnt_inst_cy_254_1338 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_1,
      IB => rx_input_memio_macnt_inst_cy_253,
      SEL => rx_input_memio_macnt_inst_lut3_56,
      O => rx_input_memio_macnt_70_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_219_1339 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_253,
      I1 => rx_input_memio_macnt_inst_lut3_56,
      O => rx_input_memio_macnt_inst_sum_219
    );
  tx_input_dh_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(13),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_13_FFX_RST,
      O => tx_input_dh(13)
    );
  tx_input_dh_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_13_FFX_RST
    );
  rx_input_memio_macnt_71_LOGIC_ZERO_1340 : X_ZERO
    port map (
      O => rx_input_memio_macnt_71_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_255_1341 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_71_LOGIC_ZERO,
      IB => rx_input_memio_macnt_71_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_57,
      O => rx_input_memio_macnt_inst_cy_255
    );
  rx_input_memio_macnt_inst_sum_220_1342 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_71_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_57,
      O => rx_input_memio_macnt_inst_sum_220
    );
  rx_input_memio_macnt_inst_lut3_571 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bp(1),
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_71,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_macnt_inst_lut3_57
    );
  rx_input_memio_macnt_inst_lut3_581 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bp(2),
      ADR2 => rx_input_memio_macnt_72,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_macnt_inst_lut3_58
    );
  rx_input_memio_macnt_71_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_71_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_256
    );
  rx_input_memio_macnt_inst_cy_256_1343 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_71_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_255,
      SEL => rx_input_memio_macnt_inst_lut3_58,
      O => rx_input_memio_macnt_71_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_221_1344 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_255,
      I1 => rx_input_memio_macnt_inst_lut3_58,
      O => rx_input_memio_macnt_inst_sum_221
    );
  rx_input_memio_macnt_71_CYINIT_1345 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_254,
      O => rx_input_memio_macnt_71_CYINIT
    );
  rx_input_memio_macnt_73_LOGIC_ZERO_1346 : X_ZERO
    port map (
      O => rx_input_memio_macnt_73_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_257_1347 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_73_LOGIC_ZERO,
      IB => rx_input_memio_macnt_73_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_59,
      O => rx_input_memio_macnt_inst_cy_257
    );
  rx_input_memio_macnt_inst_sum_222_1348 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_73_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_59,
      O => rx_input_memio_macnt_inst_sum_222
    );
  rx_input_memio_macnt_inst_lut3_591 : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_macnt_73,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => rx_input_memio_bp(3),
      O => rx_input_memio_macnt_inst_lut3_59
    );
  rx_input_memio_macnt_inst_lut3_601 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bp(4),
      ADR2 => rx_input_memio_macnt_74,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_macnt_inst_lut3_60
    );
  rx_input_memio_macnt_73_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_73_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_258
    );
  rx_input_memio_macnt_inst_cy_258_1349 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_73_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_257,
      SEL => rx_input_memio_macnt_inst_lut3_60,
      O => rx_input_memio_macnt_73_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_223_1350 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_257,
      I1 => rx_input_memio_macnt_inst_lut3_60,
      O => rx_input_memio_macnt_inst_sum_223
    );
  rx_input_memio_macnt_73_CYINIT_1351 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_256,
      O => rx_input_memio_macnt_73_CYINIT
    );
  rx_input_memio_macnt_75_LOGIC_ZERO_1352 : X_ZERO
    port map (
      O => rx_input_memio_macnt_75_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_259_1353 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_75_LOGIC_ZERO,
      IB => rx_input_memio_macnt_75_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_61,
      O => rx_input_memio_macnt_inst_cy_259
    );
  rx_input_memio_macnt_inst_sum_224_1354 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_75_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_61,
      O => rx_input_memio_macnt_inst_sum_224
    );
  rx_input_memio_macnt_inst_lut3_611 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_macnt_75,
      ADR2 => rx_input_memio_bp(5),
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_macnt_inst_lut3_61
    );
  rx_input_memio_macnt_inst_lut3_621 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bp(6),
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => rx_input_memio_macnt_76,
      O => rx_input_memio_macnt_inst_lut3_62
    );
  rx_input_memio_macnt_75_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_75_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_260
    );
  rx_input_memio_macnt_inst_cy_260_1355 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_75_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_259,
      SEL => rx_input_memio_macnt_inst_lut3_62,
      O => rx_input_memio_macnt_75_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_225_1356 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_259,
      I1 => rx_input_memio_macnt_inst_lut3_62,
      O => rx_input_memio_macnt_inst_sum_225
    );
  rx_input_memio_macnt_75_CYINIT_1357 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_258,
      O => rx_input_memio_macnt_75_CYINIT
    );
  rx_input_memio_macnt_77_LOGIC_ZERO_1358 : X_ZERO
    port map (
      O => rx_input_memio_macnt_77_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_261_1359 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_77_LOGIC_ZERO,
      IB => rx_input_memio_macnt_77_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_63,
      O => rx_input_memio_macnt_inst_cy_261
    );
  rx_input_memio_macnt_inst_sum_226_1360 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_77_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_63,
      O => rx_input_memio_macnt_inst_sum_226
    );
  rx_input_memio_macnt_inst_lut3_631 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => rx_input_memio_bp(7),
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => rx_input_memio_macnt_77,
      O => rx_input_memio_macnt_inst_lut3_63
    );
  rx_input_memio_macnt_inst_lut3_641 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => rx_input_memio_macnt_78,
      ADR3 => rx_input_memio_bp(8),
      O => rx_input_memio_macnt_inst_lut3_64
    );
  rx_input_memio_macnt_77_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_77_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_262
    );
  rx_input_memio_macnt_inst_cy_262_1361 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_77_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_261,
      SEL => rx_input_memio_macnt_inst_lut3_64,
      O => rx_input_memio_macnt_77_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_227_1362 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_261,
      I1 => rx_input_memio_macnt_inst_lut3_64,
      O => rx_input_memio_macnt_inst_sum_227
    );
  rx_input_memio_macnt_77_CYINIT_1363 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_260,
      O => rx_input_memio_macnt_77_CYINIT
    );
  rx_input_memio_macnt_79_LOGIC_ZERO_1364 : X_ZERO
    port map (
      O => rx_input_memio_macnt_79_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_263_1365 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_79_LOGIC_ZERO,
      IB => rx_input_memio_macnt_79_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_65,
      O => rx_input_memio_macnt_inst_cy_263
    );
  rx_input_memio_macnt_inst_sum_228_1366 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_79_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_65,
      O => rx_input_memio_macnt_inst_sum_228
    );
  rx_input_memio_macnt_inst_lut3_651 : X_LUT4
    generic map(
      INIT => X"D8D8"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => rx_input_memio_bp(9),
      ADR2 => rx_input_memio_macnt_79,
      ADR3 => VCC,
      O => rx_input_memio_macnt_inst_lut3_65
    );
  rx_input_memio_macnt_inst_lut3_661 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => rx_input_memio_macnt_80,
      ADR3 => rx_input_memio_bp(10),
      O => rx_input_memio_macnt_inst_lut3_66
    );
  rx_input_memio_macnt_79_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_79_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_264
    );
  rx_input_memio_macnt_inst_cy_264_1367 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_79_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_263,
      SEL => rx_input_memio_macnt_inst_lut3_66,
      O => rx_input_memio_macnt_79_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_229_1368 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_263,
      I1 => rx_input_memio_macnt_inst_lut3_66,
      O => rx_input_memio_macnt_inst_sum_229
    );
  rx_input_memio_macnt_79_CYINIT_1369 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_262,
      O => rx_input_memio_macnt_79_CYINIT
    );
  rx_input_memio_macnt_81_LOGIC_ZERO_1370 : X_ZERO
    port map (
      O => rx_input_memio_macnt_81_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_265_1371 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_81_LOGIC_ZERO,
      IB => rx_input_memio_macnt_81_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_67,
      O => rx_input_memio_macnt_inst_cy_265
    );
  rx_input_memio_macnt_inst_sum_230_1372 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_81_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_67,
      O => rx_input_memio_macnt_inst_sum_230
    );
  rx_input_memio_macnt_inst_lut3_671 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bp(11),
      ADR3 => rx_input_memio_macnt_81,
      O => rx_input_memio_macnt_inst_lut3_67
    );
  rx_input_memio_macnt_inst_lut3_681 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => rx_input_memio_macnt_82,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bp(12),
      O => rx_input_memio_macnt_inst_lut3_68
    );
  rx_input_memio_macnt_81_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_81_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_266
    );
  rx_input_memio_macnt_inst_cy_266_1373 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_81_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_265,
      SEL => rx_input_memio_macnt_inst_lut3_68,
      O => rx_input_memio_macnt_81_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_231_1374 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_265,
      I1 => rx_input_memio_macnt_inst_lut3_68,
      O => rx_input_memio_macnt_inst_sum_231
    );
  rx_input_memio_macnt_81_CYINIT_1375 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_264,
      O => rx_input_memio_macnt_81_CYINIT
    );
  rx_input_memio_macnt_83_LOGIC_ZERO_1376 : X_ZERO
    port map (
      O => rx_input_memio_macnt_83_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_267_1377 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_83_LOGIC_ZERO,
      IB => rx_input_memio_macnt_83_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_69,
      O => rx_input_memio_macnt_inst_cy_267
    );
  rx_input_memio_macnt_inst_sum_232_1378 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_83_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_69,
      O => rx_input_memio_macnt_inst_sum_232
    );
  rx_input_memio_macnt_inst_lut3_691 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => rx_input_memio_macnt_83,
      ADR2 => rx_input_memio_bp(13),
      ADR3 => VCC,
      O => rx_input_memio_macnt_inst_lut3_69
    );
  rx_input_memio_macnt_inst_lut3_701 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_84,
      ADR3 => rx_input_memio_bp(14),
      O => rx_input_memio_macnt_inst_lut3_70
    );
  rx_input_memio_macnt_83_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_83_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_268
    );
  rx_input_memio_macnt_inst_cy_268_1379 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_83_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_267,
      SEL => rx_input_memio_macnt_inst_lut3_70,
      O => rx_input_memio_macnt_83_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_233_1380 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_267,
      I1 => rx_input_memio_macnt_inst_lut3_70,
      O => rx_input_memio_macnt_inst_sum_233
    );
  rx_input_memio_macnt_83_CYINIT_1381 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_266,
      O => rx_input_memio_macnt_83_CYINIT
    );
  rx_input_memio_macnt_inst_sum_234_1382 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_85_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_71,
      O => rx_input_memio_macnt_inst_sum_234
    );
  rx_input_memio_macnt_inst_lut3_711 : X_LUT4
    generic map(
      INIT => X"F3C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => rx_input_memio_bp(15),
      ADR3 => rx_input_memio_macnt_85,
      O => rx_input_memio_macnt_inst_lut3_71
    );
  rx_input_memio_macnt_85_CYINIT_1383 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_268,
      O => rx_input_memio_macnt_85_CYINIT
    );
  rx_output_n0070_2_LOGIC_ZERO_1384 : X_ZERO
    port map (
      O => rx_output_n0070_2_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_63_1385 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_19,
      IB => rx_output_n0070_2_LOGIC_ZERO,
      SEL => rx_output_Madd_n0047_inst_lut2_64,
      O => rx_output_Madd_n0047_inst_cy_63
    );
  rx_output_Madd_n0047_inst_lut2_641 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_19,
      ADR1 => rx_output_len(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_Madd_n0047_inst_lut2_64
    );
  rx_output_n0070_2_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_34,
      ADR1 => rx_output_len(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_2_GROM
    );
  rx_output_n0070_2_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_2_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_64
    );
  rx_output_n0070_2_YUSED : X_BUF
    port map (
      I => rx_output_n0070_2_XORG,
      O => rx_output_n0070(2)
    );
  rx_output_Madd_n0047_inst_cy_64_1386 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_34,
      IB => rx_output_Madd_n0047_inst_cy_63,
      SEL => rx_output_n0070_2_GROM,
      O => rx_output_n0070_2_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_65 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_63,
      I1 => rx_output_n0070_2_GROM,
      O => rx_output_n0070_2_XORG
    );
  rx_output_n0070_3_LOGIC_ZERO_1387 : X_ZERO
    port map (
      O => rx_output_n0070_3_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_65_1388 : X_MUX2
    port map (
      IA => rx_output_n0070_3_LOGIC_ZERO,
      IB => rx_output_n0070_3_CYINIT,
      SEL => rx_output_n0070_3_FROM,
      O => rx_output_Madd_n0047_inst_cy_65
    );
  rx_output_Madd_n0047_inst_sum_66 : X_XOR2
    port map (
      I0 => rx_output_n0070_3_CYINIT,
      I1 => rx_output_n0070_3_FROM,
      O => rx_output_n0070_3_XORF
    );
  rx_output_n0070_3_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_3_FROM
    );
  rx_output_n0070_3_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(4),
      O => rx_output_n0070_3_GROM
    );
  rx_output_n0070_3_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_3_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_66
    );
  rx_output_n0070_3_XUSED : X_BUF
    port map (
      I => rx_output_n0070_3_XORF,
      O => rx_output_n0070(3)
    );
  rx_output_n0070_3_YUSED : X_BUF
    port map (
      I => rx_output_n0070_3_XORG,
      O => rx_output_n0070(4)
    );
  rx_output_Madd_n0047_inst_cy_66_1389 : X_MUX2
    port map (
      IA => rx_output_n0070_3_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_65,
      SEL => rx_output_n0070_3_GROM,
      O => rx_output_n0070_3_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_67 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_65,
      I1 => rx_output_n0070_3_GROM,
      O => rx_output_n0070_3_XORG
    );
  rx_output_n0070_3_CYINIT_1390 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_64,
      O => rx_output_n0070_3_CYINIT
    );
  rx_output_n0070_5_LOGIC_ZERO_1391 : X_ZERO
    port map (
      O => rx_output_n0070_5_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_67_1392 : X_MUX2
    port map (
      IA => rx_output_n0070_5_LOGIC_ZERO,
      IB => rx_output_n0070_5_CYINIT,
      SEL => rx_output_n0070_5_FROM,
      O => rx_output_Madd_n0047_inst_cy_67
    );
  rx_output_Madd_n0047_inst_sum_68 : X_XOR2
    port map (
      I0 => rx_output_n0070_5_CYINIT,
      I1 => rx_output_n0070_5_FROM,
      O => rx_output_n0070_5_XORF
    );
  rx_output_n0070_5_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_5_FROM
    );
  rx_output_n0070_5_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(6),
      O => rx_output_n0070_5_GROM
    );
  rx_output_n0070_5_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_5_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_68
    );
  rx_output_n0070_5_XUSED : X_BUF
    port map (
      I => rx_output_n0070_5_XORF,
      O => rx_output_n0070(5)
    );
  rx_output_n0070_5_YUSED : X_BUF
    port map (
      I => rx_output_n0070_5_XORG,
      O => rx_output_n0070(6)
    );
  rx_output_Madd_n0047_inst_cy_68_1393 : X_MUX2
    port map (
      IA => rx_output_n0070_5_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_67,
      SEL => rx_output_n0070_5_GROM,
      O => rx_output_n0070_5_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_69 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_67,
      I1 => rx_output_n0070_5_GROM,
      O => rx_output_n0070_5_XORG
    );
  rx_output_n0070_5_CYINIT_1394 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_66,
      O => rx_output_n0070_5_CYINIT
    );
  tx_input_dh_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(15),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_15_FFX_RST,
      O => tx_input_dh(15)
    );
  tx_input_dh_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_15_FFX_RST
    );
  rx_output_n0070_7_LOGIC_ZERO_1395 : X_ZERO
    port map (
      O => rx_output_n0070_7_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_69_1396 : X_MUX2
    port map (
      IA => rx_output_n0070_7_LOGIC_ZERO,
      IB => rx_output_n0070_7_CYINIT,
      SEL => rx_output_n0070_7_FROM,
      O => rx_output_Madd_n0047_inst_cy_69
    );
  rx_output_Madd_n0047_inst_sum_70 : X_XOR2
    port map (
      I0 => rx_output_n0070_7_CYINIT,
      I1 => rx_output_n0070_7_FROM,
      O => rx_output_n0070_7_XORF
    );
  rx_output_n0070_7_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_7_FROM
    );
  rx_output_n0070_7_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_7_GROM
    );
  rx_output_n0070_7_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_7_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_70
    );
  rx_output_n0070_7_XUSED : X_BUF
    port map (
      I => rx_output_n0070_7_XORF,
      O => rx_output_n0070(7)
    );
  rx_output_n0070_7_YUSED : X_BUF
    port map (
      I => rx_output_n0070_7_XORG,
      O => rx_output_n0070(8)
    );
  rx_output_Madd_n0047_inst_cy_70_1397 : X_MUX2
    port map (
      IA => rx_output_n0070_7_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_69,
      SEL => rx_output_n0070_7_GROM,
      O => rx_output_n0070_7_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_71 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_69,
      I1 => rx_output_n0070_7_GROM,
      O => rx_output_n0070_7_XORG
    );
  rx_output_n0070_7_CYINIT_1398 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_68,
      O => rx_output_n0070_7_CYINIT
    );
  rx_output_n0070_9_LOGIC_ZERO_1399 : X_ZERO
    port map (
      O => rx_output_n0070_9_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_71_1400 : X_MUX2
    port map (
      IA => rx_output_n0070_9_LOGIC_ZERO,
      IB => rx_output_n0070_9_CYINIT,
      SEL => rx_output_n0070_9_FROM,
      O => rx_output_Madd_n0047_inst_cy_71
    );
  rx_output_Madd_n0047_inst_sum_72 : X_XOR2
    port map (
      I0 => rx_output_n0070_9_CYINIT,
      I1 => rx_output_n0070_9_FROM,
      O => rx_output_n0070_9_XORF
    );
  rx_output_n0070_9_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(9),
      ADR3 => VCC,
      O => rx_output_n0070_9_FROM
    );
  rx_output_n0070_9_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_9_GROM
    );
  rx_output_n0070_9_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_9_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_72
    );
  rx_output_n0070_9_XUSED : X_BUF
    port map (
      I => rx_output_n0070_9_XORF,
      O => rx_output_n0070(9)
    );
  rx_output_n0070_9_YUSED : X_BUF
    port map (
      I => rx_output_n0070_9_XORG,
      O => rx_output_n0070(10)
    );
  rx_output_Madd_n0047_inst_cy_72_1401 : X_MUX2
    port map (
      IA => rx_output_n0070_9_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_71,
      SEL => rx_output_n0070_9_GROM,
      O => rx_output_n0070_9_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_73 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_71,
      I1 => rx_output_n0070_9_GROM,
      O => rx_output_n0070_9_XORG
    );
  rx_output_n0070_9_CYINIT_1402 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_70,
      O => rx_output_n0070_9_CYINIT
    );
  rx_output_n0070_11_LOGIC_ZERO_1403 : X_ZERO
    port map (
      O => rx_output_n0070_11_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_73_1404 : X_MUX2
    port map (
      IA => rx_output_n0070_11_LOGIC_ZERO,
      IB => rx_output_n0070_11_CYINIT,
      SEL => rx_output_n0070_11_FROM,
      O => rx_output_Madd_n0047_inst_cy_73
    );
  rx_output_Madd_n0047_inst_sum_74 : X_XOR2
    port map (
      I0 => rx_output_n0070_11_CYINIT,
      I1 => rx_output_n0070_11_FROM,
      O => rx_output_n0070_11_XORF
    );
  rx_output_n0070_11_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(11),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_11_FROM
    );
  rx_output_n0070_11_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(12),
      O => rx_output_n0070_11_GROM
    );
  rx_output_n0070_11_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_11_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_74
    );
  rx_output_n0070_11_XUSED : X_BUF
    port map (
      I => rx_output_n0070_11_XORF,
      O => rx_output_n0070(11)
    );
  rx_output_n0070_11_YUSED : X_BUF
    port map (
      I => rx_output_n0070_11_XORG,
      O => rx_output_n0070(12)
    );
  rx_output_Madd_n0047_inst_cy_74_1405 : X_MUX2
    port map (
      IA => rx_output_n0070_11_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_73,
      SEL => rx_output_n0070_11_GROM,
      O => rx_output_n0070_11_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_75 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_73,
      I1 => rx_output_n0070_11_GROM,
      O => rx_output_n0070_11_XORG
    );
  rx_output_n0070_11_CYINIT_1406 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_72,
      O => rx_output_n0070_11_CYINIT
    );
  rx_output_n0070_13_LOGIC_ZERO_1407 : X_ZERO
    port map (
      O => rx_output_n0070_13_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_75_1408 : X_MUX2
    port map (
      IA => rx_output_n0070_13_LOGIC_ZERO,
      IB => rx_output_n0070_13_CYINIT,
      SEL => rx_output_n0070_13_FROM,
      O => rx_output_Madd_n0047_inst_cy_75
    );
  rx_output_Madd_n0047_inst_sum_76 : X_XOR2
    port map (
      I0 => rx_output_n0070_13_CYINIT,
      I1 => rx_output_n0070_13_FROM,
      O => rx_output_n0070_13_XORF
    );
  rx_output_n0070_13_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_13_FROM
    );
  rx_output_n0070_13_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(14),
      O => rx_output_n0070_13_GROM
    );
  rx_output_n0070_13_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_13_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_76
    );
  rx_output_n0070_13_XUSED : X_BUF
    port map (
      I => rx_output_n0070_13_XORF,
      O => rx_output_n0070(13)
    );
  rx_output_n0070_13_YUSED : X_BUF
    port map (
      I => rx_output_n0070_13_XORG,
      O => rx_output_n0070(14)
    );
  rx_output_Madd_n0047_inst_cy_76_1409 : X_MUX2
    port map (
      IA => rx_output_n0070_13_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_75,
      SEL => rx_output_n0070_13_GROM,
      O => rx_output_n0070_13_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_77 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_75,
      I1 => rx_output_n0070_13_GROM,
      O => rx_output_n0070_13_XORG
    );
  rx_output_n0070_13_CYINIT_1410 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_74,
      O => rx_output_n0070_13_CYINIT
    );
  rx_output_Madd_n0047_inst_sum_78 : X_XOR2
    port map (
      I0 => rx_output_n0070_15_CYINIT,
      I1 => rx_output_SIG_45,
      O => rx_output_n0070_15_XORF
    );
  rx_output_BEL_20 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(15),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_SIG_45
    );
  rx_output_n0070_15_XUSED : X_BUF
    port map (
      I => rx_output_n0070_15_XORF,
      O => rx_output_n0070(15)
    );
  rx_output_n0070_15_CYINIT_1411 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_76,
      O => rx_output_n0070_15_CYINIT
    );
  tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ONE_1412 : X_ONE
    port map (
      O => tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ONE
    );
  tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ZERO_1413 : X_ZERO
    port map (
      O => tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ZERO
    );
  tx_output_Mcompar_n0006_inst_cy_78_1414 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ONE,
      SEL => tx_output_Mcompar_n0006_inst_lut4_0,
      O => tx_output_Mcompar_n0006_inst_cy_78
    );
  tx_output_Mcompar_n0006_inst_lut4_01 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => tx_output_addrl(0),
      ADR1 => tx_output_bpl(1),
      ADR2 => tx_output_addrl(1),
      ADR3 => tx_output_bpl(0),
      O => tx_output_Mcompar_n0006_inst_lut4_0
    );
  tx_output_Mcompar_n0006_inst_lut4_11 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => tx_output_addrl(2),
      ADR1 => tx_output_addrl(3),
      ADR2 => tx_output_bpl(3),
      ADR3 => tx_output_bpl(2),
      O => tx_output_Mcompar_n0006_inst_lut4_1
    );
  tx_output_Mcompar_n0006_inst_cy_79_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_79_CYMUXG,
      O => tx_output_Mcompar_n0006_inst_cy_79
    );
  tx_output_Mcompar_n0006_inst_cy_79_1415 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_78,
      SEL => tx_output_Mcompar_n0006_inst_lut4_1,
      O => tx_output_Mcompar_n0006_inst_cy_79_CYMUXG
    );
  tx_output_Mcompar_n0006_inst_cy_81_LOGIC_ZERO_1416 : X_ZERO
    port map (
      O => tx_output_Mcompar_n0006_inst_cy_81_LOGIC_ZERO
    );
  tx_output_Mcompar_n0006_inst_cy_80_1417 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_81_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_81_CYINIT,
      SEL => tx_output_Mcompar_n0006_inst_lut4_2,
      O => tx_output_Mcompar_n0006_inst_cy_80
    );
  tx_output_Mcompar_n0006_inst_lut4_21 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => tx_output_addrl(4),
      ADR1 => tx_output_addrl(5),
      ADR2 => tx_output_bpl(5),
      ADR3 => tx_output_bpl(4),
      O => tx_output_Mcompar_n0006_inst_lut4_2
    );
  tx_output_Mcompar_n0006_inst_lut4_31 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => tx_output_addrl(6),
      ADR1 => tx_output_addrl(7),
      ADR2 => tx_output_bpl(6),
      ADR3 => tx_output_bpl(7),
      O => tx_output_Mcompar_n0006_inst_lut4_3
    );
  tx_output_Mcompar_n0006_inst_cy_81_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_81_CYMUXG,
      O => tx_output_Mcompar_n0006_inst_cy_81
    );
  tx_output_Mcompar_n0006_inst_cy_81_1418 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_81_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_80,
      SEL => tx_output_Mcompar_n0006_inst_lut4_3,
      O => tx_output_Mcompar_n0006_inst_cy_81_CYMUXG
    );
  tx_output_Mcompar_n0006_inst_cy_81_CYINIT_1419 : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_79,
      O => tx_output_Mcompar_n0006_inst_cy_81_CYINIT
    );
  tx_output_Mcompar_n0006_inst_cy_83_LOGIC_ZERO_1420 : X_ZERO
    port map (
      O => tx_output_Mcompar_n0006_inst_cy_83_LOGIC_ZERO
    );
  tx_output_Mcompar_n0006_inst_cy_82_1421 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_83_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_83_CYINIT,
      SEL => tx_output_Mcompar_n0006_inst_lut4_4,
      O => tx_output_Mcompar_n0006_inst_cy_82
    );
  tx_output_Mcompar_n0006_inst_lut4_41 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => tx_output_bpl(9),
      ADR1 => tx_output_bpl(8),
      ADR2 => tx_output_addrl(8),
      ADR3 => tx_output_addrl(9),
      O => tx_output_Mcompar_n0006_inst_lut4_4
    );
  tx_output_Mcompar_n0006_inst_lut4_51 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => tx_output_addrl(10),
      ADR1 => tx_output_bpl(11),
      ADR2 => tx_output_bpl(10),
      ADR3 => tx_output_addrl(11),
      O => tx_output_Mcompar_n0006_inst_lut4_5
    );
  tx_output_Mcompar_n0006_inst_cy_83_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_83_CYMUXG,
      O => tx_output_Mcompar_n0006_inst_cy_83
    );
  tx_output_Mcompar_n0006_inst_cy_83_1422 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_83_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_82,
      SEL => tx_output_Mcompar_n0006_inst_lut4_5,
      O => tx_output_Mcompar_n0006_inst_cy_83_CYMUXG
    );
  tx_output_Mcompar_n0006_inst_cy_83_CYINIT_1423 : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_81,
      O => tx_output_Mcompar_n0006_inst_cy_83_CYINIT
    );
  rx_input_GMII_INCE : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_lince,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_ince_FFX_RST,
      O => rx_input_ince
    );
  rx_input_ince_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_ince_FFX_RST
    );
  tx_output_n0006_LOGIC_ZERO_1424 : X_ZERO
    port map (
      O => tx_output_n0006_LOGIC_ZERO
    );
  tx_output_Mcompar_n0006_inst_cy_84_1425 : X_MUX2
    port map (
      IA => tx_output_n0006_LOGIC_ZERO,
      IB => tx_output_n0006_CYINIT,
      SEL => tx_output_Mcompar_n0006_inst_lut4_6,
      O => tx_output_Mcompar_n0006_inst_cy_84
    );
  tx_output_Mcompar_n0006_inst_lut4_61 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => tx_output_addrl(12),
      ADR1 => tx_output_addrl(13),
      ADR2 => tx_output_bpl(13),
      ADR3 => tx_output_bpl(12),
      O => tx_output_Mcompar_n0006_inst_lut4_6
    );
  tx_output_Mcompar_n0006_inst_lut4_71 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => tx_output_addrl(14),
      ADR1 => tx_output_addrl(15),
      ADR2 => tx_output_bpl(14),
      ADR3 => tx_output_bpl(15),
      O => tx_output_Mcompar_n0006_inst_lut4_7
    );
  tx_output_n0006_COUTUSED : X_BUF
    port map (
      I => tx_output_n0006_CYMUXG,
      O => tx_output_n0006
    );
  tx_output_Mcompar_n0006_inst_cy_85 : X_MUX2
    port map (
      IA => tx_output_n0006_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_84,
      SEL => tx_output_Mcompar_n0006_inst_lut4_7,
      O => tx_output_n0006_CYMUXG
    );
  tx_output_n0006_CYINIT_1426 : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_83,
      O => tx_output_n0006_CYINIT
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ONE_1427 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ZERO_1428 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_177_1429 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(41),
      ADR1 => rx_input_memio_addrchk_datal(40),
      ADR2 => rx_input_memio_addrchk_datal(41),
      ADR3 => rx_input_memio_addrchk_macaddrl(40),
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(42),
      ADR1 => rx_input_memio_addrchk_macaddrl(43),
      ADR2 => rx_input_memio_addrchk_datal(43),
      ADR3 => rx_input_memio_addrchk_datal(42),
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_1430 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_0_LOGIC_ZERO_1431 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_0_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_179_1432 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_0_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_0_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(44),
      ADR1 => rx_input_memio_addrchk_macaddrl(45),
      ADR2 => rx_input_memio_addrchk_datal(45),
      ADR3 => rx_input_memio_addrchk_datal(44),
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(46),
      ADR1 => rx_input_memio_addrchk_macaddrl(47),
      ADR2 => rx_input_memio_addrchk_datal(47),
      ADR3 => rx_input_memio_addrchk_datal(46),
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_0_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_0_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(0)
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_0_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_0_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_0_CYINIT_1433 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_0_CYINIT
    );
  rx_input_memio_bcntl_0_LOGIC_ONE_1434 : X_ONE
    port map (
      O => rx_input_memio_bcntl_0_LOGIC_ONE
    );
  rx_input_memio_Msub_n0042_inst_cy_237_1435 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_86,
      IB => rx_input_memio_bcntl_0_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_149,
      O => rx_input_memio_Msub_n0042_inst_cy_237
    );
  rx_input_memio_Msub_n0042_inst_sum_203 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_0_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_149,
      O => rx_input_memio_n0042(0)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1491 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_86,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_149
    );
  rx_input_memio_Msub_n0042_inst_lut2_1501 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_87,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_150
    );
  rx_input_memio_bcntl_0_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_0_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_238
    );
  rx_input_memio_Msub_n0042_inst_cy_238_1436 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_87,
      IB => rx_input_memio_Msub_n0042_inst_cy_237,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_150,
      O => rx_input_memio_bcntl_0_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_204 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_237,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_150,
      O => rx_input_memio_n0042(1)
    );
  rx_input_memio_bcntl_0_CYINIT_1437 : X_BUF
    port map (
      I => rx_input_memio_bcntl_0_LOGIC_ONE,
      O => rx_input_memio_bcntl_0_CYINIT
    );
  rx_input_memio_bcntl_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_2_FFY_RST
    );
  rx_input_memio_bcntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(3),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_2_FFY_RST,
      O => rx_input_memio_bcntl(3)
    );
  rx_input_memio_Msub_n0042_inst_cy_239_1438 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_7,
      IB => rx_input_memio_bcntl_2_CYINIT,
      SEL => rx_input_memio_bcntl_2_FROM,
      O => rx_input_memio_Msub_n0042_inst_cy_239
    );
  rx_input_memio_Msub_n0042_inst_sum_205 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_2_CYINIT,
      I1 => rx_input_memio_bcntl_2_FROM,
      O => rx_input_memio_n0042(2)
    );
  rx_input_memio_bcntl_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_7,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bcnt_88,
      O => rx_input_memio_bcntl_2_FROM
    );
  rx_input_memio_Msub_n0042_inst_lut2_1521 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_89,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_152
    );
  rx_input_memio_bcntl_2_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_2_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_240
    );
  rx_input_memio_Msub_n0042_inst_cy_240_1439 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_89,
      IB => rx_input_memio_Msub_n0042_inst_cy_239,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_152,
      O => rx_input_memio_bcntl_2_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_206 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_239,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_152,
      O => rx_input_memio_n0042(3)
    );
  rx_input_memio_bcntl_2_CYINIT_1440 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_238,
      O => rx_input_memio_bcntl_2_CYINIT
    );
  rx_input_memio_bcntl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_4_FFY_RST
    );
  rx_input_memio_bcntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(5),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_4_FFY_RST,
      O => rx_input_memio_bcntl(5)
    );
  rx_input_memio_Msub_n0042_inst_cy_241_1441 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_90,
      IB => rx_input_memio_bcntl_4_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_153,
      O => rx_input_memio_Msub_n0042_inst_cy_241
    );
  rx_input_memio_Msub_n0042_inst_sum_207 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_4_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_153,
      O => rx_input_memio_n0042(4)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1531 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_90,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_153
    );
  rx_input_memio_Msub_n0042_inst_lut2_1541 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_91,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_154
    );
  rx_input_memio_bcntl_4_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_4_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_242
    );
  rx_input_memio_Msub_n0042_inst_cy_242_1442 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_91,
      IB => rx_input_memio_Msub_n0042_inst_cy_241,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_154,
      O => rx_input_memio_bcntl_4_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_208 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_241,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_154,
      O => rx_input_memio_n0042(5)
    );
  rx_input_memio_bcntl_4_CYINIT_1443 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_240,
      O => rx_input_memio_bcntl_4_CYINIT
    );
  rx_input_memio_bcntl_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_6_FFY_RST
    );
  rx_input_memio_bcntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(7),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_6_FFY_RST,
      O => rx_input_memio_bcntl(7)
    );
  rx_input_memio_Msub_n0042_inst_cy_243_1444 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_92,
      IB => rx_input_memio_bcntl_6_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_155,
      O => rx_input_memio_Msub_n0042_inst_cy_243
    );
  rx_input_memio_Msub_n0042_inst_sum_209 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_6_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_155,
      O => rx_input_memio_n0042(6)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1551 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_92,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_155
    );
  rx_input_memio_Msub_n0042_inst_lut2_1561 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_93,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_156
    );
  rx_input_memio_bcntl_6_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_6_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_244
    );
  rx_input_memio_Msub_n0042_inst_cy_244_1445 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_93,
      IB => rx_input_memio_Msub_n0042_inst_cy_243,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_156,
      O => rx_input_memio_bcntl_6_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_210 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_243,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_156,
      O => rx_input_memio_n0042(7)
    );
  rx_input_memio_bcntl_6_CYINIT_1446 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_242,
      O => rx_input_memio_bcntl_6_CYINIT
    );
  rx_input_memio_bcntl_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_8_FFY_RST
    );
  rx_input_memio_bcntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(9),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_8_FFY_RST,
      O => rx_input_memio_bcntl(9)
    );
  rx_input_memio_Msub_n0042_inst_cy_245_1447 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_94,
      IB => rx_input_memio_bcntl_8_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_157,
      O => rx_input_memio_Msub_n0042_inst_cy_245
    );
  rx_input_memio_Msub_n0042_inst_sum_211 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_8_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_157,
      O => rx_input_memio_n0042(8)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1571 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_94,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_157
    );
  rx_input_memio_Msub_n0042_inst_lut2_1581 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_95,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_158
    );
  rx_input_memio_bcntl_8_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_8_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_246
    );
  rx_input_memio_Msub_n0042_inst_cy_246_1448 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_95,
      IB => rx_input_memio_Msub_n0042_inst_cy_245,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_158,
      O => rx_input_memio_bcntl_8_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_212 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_245,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_158,
      O => rx_input_memio_n0042(9)
    );
  rx_input_memio_bcntl_8_CYINIT_1449 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_244,
      O => rx_input_memio_bcntl_8_CYINIT
    );
  rx_input_memio_bcntl_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_10_FFY_RST
    );
  rx_input_memio_bcntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(11),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_10_FFY_RST,
      O => rx_input_memio_bcntl(11)
    );
  rx_input_memio_Msub_n0042_inst_cy_247_1450 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_96,
      IB => rx_input_memio_bcntl_10_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_159,
      O => rx_input_memio_Msub_n0042_inst_cy_247
    );
  rx_input_memio_Msub_n0042_inst_sum_213 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_10_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_159,
      O => rx_input_memio_n0042(10)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1591 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_96,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_159
    );
  rx_input_memio_Msub_n0042_inst_lut2_1601 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_97,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_160
    );
  rx_input_memio_bcntl_10_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_10_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_248
    );
  rx_input_memio_Msub_n0042_inst_cy_248_1451 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_97,
      IB => rx_input_memio_Msub_n0042_inst_cy_247,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_160,
      O => rx_input_memio_bcntl_10_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_214 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_247,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_160,
      O => rx_input_memio_n0042(11)
    );
  rx_input_memio_bcntl_10_CYINIT_1452 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_246,
      O => rx_input_memio_bcntl_10_CYINIT
    );
  tx_input_dl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(10),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_11_FFY_RST,
      O => tx_input_dl(10)
    );
  tx_input_dl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_11_FFY_RST
    );
  rx_input_memio_bcntl_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_12_FFY_RST
    );
  rx_input_memio_bcntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(13),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_12_FFY_RST,
      O => rx_input_memio_bcntl(13)
    );
  rx_input_memio_Msub_n0042_inst_cy_249_1453 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_98,
      IB => rx_input_memio_bcntl_12_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_161,
      O => rx_input_memio_Msub_n0042_inst_cy_249
    );
  rx_input_memio_Msub_n0042_inst_sum_215 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_12_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_161,
      O => rx_input_memio_n0042(12)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1611 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_98,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_161
    );
  rx_input_memio_Msub_n0042_inst_lut2_1621 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_99,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_162
    );
  rx_input_memio_bcntl_12_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_12_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_250
    );
  rx_input_memio_Msub_n0042_inst_cy_250_1454 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_99,
      IB => rx_input_memio_Msub_n0042_inst_cy_249,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_162,
      O => rx_input_memio_bcntl_12_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_216 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_249,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_162,
      O => rx_input_memio_n0042(13)
    );
  rx_input_memio_bcntl_12_CYINIT_1455 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_248,
      O => rx_input_memio_bcntl_12_CYINIT
    );
  rx_input_memio_bcntl_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_14_FFY_RST
    );
  rx_input_memio_bcntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(15),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_14_FFY_RST,
      O => rx_input_memio_bcntl(15)
    );
  rx_input_memio_Msub_n0042_inst_cy_251_1456 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_100,
      IB => rx_input_memio_bcntl_14_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_163,
      O => rx_input_memio_Msub_n0042_inst_cy_251
    );
  rx_input_memio_Msub_n0042_inst_sum_217 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_14_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_163,
      O => rx_input_memio_n0042(14)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1631 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_100,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_163
    );
  rx_input_memio_Msub_n0042_inst_lut2_1641 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_101,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_164
    );
  rx_input_memio_Msub_n0042_inst_sum_218 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_251,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_164,
      O => rx_input_memio_n0042(15)
    );
  rx_input_memio_bcntl_14_CYINIT_1457 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_250,
      O => rx_input_memio_bcntl_14_CYINIT
    );
  tx_input_addr_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_16_FFY_RST
    );
  tx_input_addr_16_1458 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_127,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_16_FFY_RST,
      O => tx_input_addr_16
    );
  tx_input_addr_16_LOGIC_ZERO_1459 : X_ZERO
    port map (
      O => tx_input_addr_16_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_134_1460 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_13,
      IB => tx_input_addr_16_LOGIC_ZERO,
      SEL => tx_input_cs_FFd12_rt,
      O => tx_input_addr_inst_cy_134
    );
  tx_input_cs_FFd12_rt_1461 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_13,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_cs_FFd12_rt
    );
  tx_input_addr_inst_lut3_161 : X_LUT4
    generic map(
      INIT => X"F3C0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_5,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => txbp(0),
      ADR3 => tx_input_addr_16,
      O => tx_input_addr_inst_lut3_16
    );
  tx_input_addr_16_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_16_CYMUXG,
      O => tx_input_addr_inst_cy_135
    );
  tx_input_addr_inst_cy_135_1462 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_5,
      IB => tx_input_addr_inst_cy_134,
      SEL => tx_input_addr_inst_lut3_16,
      O => tx_input_addr_16_CYMUXG
    );
  tx_input_addr_inst_sum_127_1463 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_134,
      I1 => tx_input_addr_inst_lut3_16,
      O => tx_input_addr_inst_sum_127
    );
  tx_input_addr_17_LOGIC_ZERO_1464 : X_ZERO
    port map (
      O => tx_input_addr_17_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_136_1465 : X_MUX2
    port map (
      IA => tx_input_addr_17_LOGIC_ZERO,
      IB => tx_input_addr_17_CYINIT,
      SEL => tx_input_addr_inst_lut3_17,
      O => tx_input_addr_inst_cy_136
    );
  tx_input_addr_inst_sum_128_1466 : X_XOR2
    port map (
      I0 => tx_input_addr_17_CYINIT,
      I1 => tx_input_addr_inst_lut3_17,
      O => tx_input_addr_inst_sum_128
    );
  tx_input_addr_inst_lut3_171 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => txbp(1),
      ADR1 => VCC,
      ADR2 => tx_input_cs_FFd12,
      ADR3 => tx_input_addr_17,
      O => tx_input_addr_inst_lut3_17
    );
  tx_input_addr_inst_lut3_181 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_addr_18,
      ADR2 => txbp(2),
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_addr_inst_lut3_18
    );
  tx_input_addr_17_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_17_CYMUXG,
      O => tx_input_addr_inst_cy_137
    );
  tx_input_addr_inst_cy_137_1467 : X_MUX2
    port map (
      IA => tx_input_addr_17_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_136,
      SEL => tx_input_addr_inst_lut3_18,
      O => tx_input_addr_17_CYMUXG
    );
  tx_input_addr_inst_sum_129_1468 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_136,
      I1 => tx_input_addr_inst_lut3_18,
      O => tx_input_addr_inst_sum_129
    );
  tx_input_addr_17_CYINIT_1469 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_135,
      O => tx_input_addr_17_CYINIT
    );
  tx_input_addr_19_LOGIC_ZERO_1470 : X_ZERO
    port map (
      O => tx_input_addr_19_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_138_1471 : X_MUX2
    port map (
      IA => tx_input_addr_19_LOGIC_ZERO,
      IB => tx_input_addr_19_CYINIT,
      SEL => tx_input_addr_inst_lut3_19,
      O => tx_input_addr_inst_cy_138
    );
  tx_input_addr_inst_sum_130_1472 : X_XOR2
    port map (
      I0 => tx_input_addr_19_CYINIT,
      I1 => tx_input_addr_inst_lut3_19,
      O => tx_input_addr_inst_sum_130
    );
  tx_input_addr_inst_lut3_191 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => txbp(3),
      ADR2 => VCC,
      ADR3 => tx_input_addr_19,
      O => tx_input_addr_inst_lut3_19
    );
  tx_input_addr_inst_lut3_201 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => txbp(4),
      ADR1 => VCC,
      ADR2 => tx_input_addr_20,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_addr_inst_lut3_20
    );
  tx_input_addr_19_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_19_CYMUXG,
      O => tx_input_addr_inst_cy_139
    );
  tx_input_addr_inst_cy_139_1473 : X_MUX2
    port map (
      IA => tx_input_addr_19_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_138,
      SEL => tx_input_addr_inst_lut3_20,
      O => tx_input_addr_19_CYMUXG
    );
  tx_input_addr_inst_sum_131_1474 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_138,
      I1 => tx_input_addr_inst_lut3_20,
      O => tx_input_addr_inst_sum_131
    );
  tx_input_addr_19_CYINIT_1475 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_137,
      O => tx_input_addr_19_CYINIT
    );
  tx_input_addr_21_LOGIC_ZERO_1476 : X_ZERO
    port map (
      O => tx_input_addr_21_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_140_1477 : X_MUX2
    port map (
      IA => tx_input_addr_21_LOGIC_ZERO,
      IB => tx_input_addr_21_CYINIT,
      SEL => tx_input_addr_inst_lut3_21,
      O => tx_input_addr_inst_cy_140
    );
  tx_input_addr_inst_sum_132_1478 : X_XOR2
    port map (
      I0 => tx_input_addr_21_CYINIT,
      I1 => tx_input_addr_inst_lut3_21,
      O => tx_input_addr_inst_sum_132
    );
  tx_input_addr_inst_lut3_211 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => VCC,
      ADR2 => tx_input_addr_21,
      ADR3 => txbp(5),
      O => tx_input_addr_inst_lut3_21
    );
  tx_input_addr_inst_lut3_221 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => txbp(6),
      ADR2 => tx_input_addr_22,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_addr_inst_lut3_22
    );
  tx_input_addr_21_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_21_CYMUXG,
      O => tx_input_addr_inst_cy_141
    );
  tx_input_addr_inst_cy_141_1479 : X_MUX2
    port map (
      IA => tx_input_addr_21_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_140,
      SEL => tx_input_addr_inst_lut3_22,
      O => tx_input_addr_21_CYMUXG
    );
  tx_input_addr_inst_sum_133_1480 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_140,
      I1 => tx_input_addr_inst_lut3_22,
      O => tx_input_addr_inst_sum_133
    );
  tx_input_addr_21_CYINIT_1481 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_139,
      O => tx_input_addr_21_CYINIT
    );
  tx_input_addr_23_LOGIC_ZERO_1482 : X_ZERO
    port map (
      O => tx_input_addr_23_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_142_1483 : X_MUX2
    port map (
      IA => tx_input_addr_23_LOGIC_ZERO,
      IB => tx_input_addr_23_CYINIT,
      SEL => tx_input_addr_inst_lut3_23,
      O => tx_input_addr_inst_cy_142
    );
  tx_input_addr_inst_sum_134_1484 : X_XOR2
    port map (
      I0 => tx_input_addr_23_CYINIT,
      I1 => tx_input_addr_inst_lut3_23,
      O => tx_input_addr_inst_sum_134
    );
  tx_input_addr_inst_lut3_231 : X_LUT4
    generic map(
      INIT => X"F3C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => txbp(7),
      ADR3 => tx_input_addr_23,
      O => tx_input_addr_inst_lut3_23
    );
  tx_input_addr_inst_lut3_241 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => txbp(8),
      ADR1 => tx_input_addr_24,
      ADR2 => tx_input_cs_FFd12,
      ADR3 => VCC,
      O => tx_input_addr_inst_lut3_24
    );
  tx_input_addr_23_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_23_CYMUXG,
      O => tx_input_addr_inst_cy_143
    );
  tx_input_addr_inst_cy_143_1485 : X_MUX2
    port map (
      IA => tx_input_addr_23_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_142,
      SEL => tx_input_addr_inst_lut3_24,
      O => tx_input_addr_23_CYMUXG
    );
  tx_input_addr_inst_sum_135_1486 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_142,
      I1 => tx_input_addr_inst_lut3_24,
      O => tx_input_addr_inst_sum_135
    );
  tx_input_addr_23_CYINIT_1487 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_141,
      O => tx_input_addr_23_CYINIT
    );
  tx_input_addr_25_LOGIC_ZERO_1488 : X_ZERO
    port map (
      O => tx_input_addr_25_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_144_1489 : X_MUX2
    port map (
      IA => tx_input_addr_25_LOGIC_ZERO,
      IB => tx_input_addr_25_CYINIT,
      SEL => tx_input_addr_inst_lut3_25,
      O => tx_input_addr_inst_cy_144
    );
  tx_input_addr_inst_sum_136_1490 : X_XOR2
    port map (
      I0 => tx_input_addr_25_CYINIT,
      I1 => tx_input_addr_inst_lut3_25,
      O => tx_input_addr_inst_sum_136
    );
  tx_input_addr_inst_lut3_251 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => txbp(9),
      ADR2 => tx_input_cs_FFd12,
      ADR3 => tx_input_addr_25,
      O => tx_input_addr_inst_lut3_25
    );
  tx_input_addr_inst_lut3_261 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => txbp(10),
      ADR1 => VCC,
      ADR2 => tx_input_addr_26,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_addr_inst_lut3_26
    );
  tx_input_addr_25_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_25_CYMUXG,
      O => tx_input_addr_inst_cy_145
    );
  tx_input_addr_inst_cy_145_1491 : X_MUX2
    port map (
      IA => tx_input_addr_25_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_144,
      SEL => tx_input_addr_inst_lut3_26,
      O => tx_input_addr_25_CYMUXG
    );
  tx_input_addr_inst_sum_137_1492 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_144,
      I1 => tx_input_addr_inst_lut3_26,
      O => tx_input_addr_inst_sum_137
    );
  tx_input_addr_25_CYINIT_1493 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_143,
      O => tx_input_addr_25_CYINIT
    );
  tx_input_addr_27_LOGIC_ZERO_1494 : X_ZERO
    port map (
      O => tx_input_addr_27_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_146_1495 : X_MUX2
    port map (
      IA => tx_input_addr_27_LOGIC_ZERO,
      IB => tx_input_addr_27_CYINIT,
      SEL => tx_input_addr_inst_lut3_27,
      O => tx_input_addr_inst_cy_146
    );
  tx_input_addr_inst_sum_138_1496 : X_XOR2
    port map (
      I0 => tx_input_addr_27_CYINIT,
      I1 => tx_input_addr_inst_lut3_27,
      O => tx_input_addr_inst_sum_138
    );
  tx_input_addr_inst_lut3_271 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => tx_input_addr_27,
      ADR3 => txbp(11),
      O => tx_input_addr_inst_lut3_27
    );
  tx_input_addr_inst_lut3_281 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => tx_input_addr_28,
      ADR3 => txbp(12),
      O => tx_input_addr_inst_lut3_28
    );
  tx_input_addr_27_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_27_CYMUXG,
      O => tx_input_addr_inst_cy_147
    );
  tx_input_addr_inst_cy_147_1497 : X_MUX2
    port map (
      IA => tx_input_addr_27_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_146,
      SEL => tx_input_addr_inst_lut3_28,
      O => tx_input_addr_27_CYMUXG
    );
  tx_input_addr_inst_sum_139_1498 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_146,
      I1 => tx_input_addr_inst_lut3_28,
      O => tx_input_addr_inst_sum_139
    );
  tx_input_addr_27_CYINIT_1499 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_145,
      O => tx_input_addr_27_CYINIT
    );
  tx_input_addr_29_LOGIC_ZERO_1500 : X_ZERO
    port map (
      O => tx_input_addr_29_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_148_1501 : X_MUX2
    port map (
      IA => tx_input_addr_29_LOGIC_ZERO,
      IB => tx_input_addr_29_CYINIT,
      SEL => tx_input_addr_inst_lut3_29,
      O => tx_input_addr_inst_cy_148
    );
  tx_input_addr_inst_sum_140_1502 : X_XOR2
    port map (
      I0 => tx_input_addr_29_CYINIT,
      I1 => tx_input_addr_inst_lut3_29,
      O => tx_input_addr_inst_sum_140
    );
  tx_input_addr_inst_lut3_291 : X_LUT4
    generic map(
      INIT => X"F3C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => txbp(13),
      ADR3 => tx_input_addr_29,
      O => tx_input_addr_inst_lut3_29
    );
  tx_input_addr_inst_lut3_301 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => tx_input_addr_30,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => VCC,
      ADR3 => txbp(14),
      O => tx_input_addr_inst_lut3_30
    );
  tx_input_addr_29_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_29_CYMUXG,
      O => tx_input_addr_inst_cy_149
    );
  tx_input_addr_inst_cy_149_1503 : X_MUX2
    port map (
      IA => tx_input_addr_29_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_148,
      SEL => tx_input_addr_inst_lut3_30,
      O => tx_input_addr_29_CYMUXG
    );
  tx_input_addr_inst_sum_141_1504 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_148,
      I1 => tx_input_addr_inst_lut3_30,
      O => tx_input_addr_inst_sum_141
    );
  tx_input_addr_29_CYINIT_1505 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_147,
      O => tx_input_addr_29_CYINIT
    );
  tx_input_addr_inst_sum_142_1506 : X_XOR2
    port map (
      I0 => tx_input_addr_31_CYINIT,
      I1 => tx_input_addr_inst_lut3_31,
      O => tx_input_addr_inst_sum_142
    );
  tx_input_addr_inst_lut3_311 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_addr_31,
      ADR2 => txbp(15),
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_addr_inst_lut3_31
    );
  tx_input_addr_31_CYINIT_1507 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_149,
      O => tx_input_addr_31_CYINIT
    );
  mac_control_rxf_cnt_0_LOGIC_ZERO_1508 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_0_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_16_1509 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_1,
      IB => mac_control_rxf_cnt_0_LOGIC_ZERO,
      SEL => mac_control_rxf_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_rxf_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(0),
      O => mac_control_rxf_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_rxf_cnt_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_56,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(1),
      O => mac_control_rxf_cnt_0_GROM
    );
  mac_control_rxf_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_0_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_17_1510 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_56,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_rxf_cnt_0_GROM,
      O => mac_control_rxf_cnt_0_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_rxf_cnt_0_GROM,
      O => mac_control_rxf_cnt_n0000(1)
    );
  mac_control_rxf_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(3),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(3)
    );
  mac_control_rxf_cnt_2_LOGIC_ZERO_1511 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_2_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_18_1512 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_2_CYINIT,
      SEL => mac_control_rxf_cnt_2_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_2_CYINIT,
      I1 => mac_control_rxf_cnt_2_FROM,
      O => mac_control_rxf_cnt_n0000(2)
    );
  mac_control_rxf_cnt_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(2),
      O => mac_control_rxf_cnt_2_FROM
    );
  mac_control_rxf_cnt_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(3),
      O => mac_control_rxf_cnt_2_GROM
    );
  mac_control_rxf_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_2_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_19_1513 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_rxf_cnt_2_GROM,
      O => mac_control_rxf_cnt_2_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_rxf_cnt_2_GROM,
      O => mac_control_rxf_cnt_n0000(3)
    );
  mac_control_rxf_cnt_2_CYINIT_1514 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_rxf_cnt_2_CYINIT
    );
  mac_control_rxf_cnt_4_LOGIC_ZERO_1515 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_4_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_20_1516 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_4_CYINIT,
      SEL => mac_control_rxf_cnt_4_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_4_CYINIT,
      I1 => mac_control_rxf_cnt_4_FROM,
      O => mac_control_rxf_cnt_n0000(4)
    );
  mac_control_rxf_cnt_4_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(4),
      O => mac_control_rxf_cnt_4_FROM
    );
  mac_control_rxf_cnt_4_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxf_cnt(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxf_cnt_4_GROM
    );
  mac_control_rxf_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_4_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_21_1517 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_rxf_cnt_4_GROM,
      O => mac_control_rxf_cnt_4_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_rxf_cnt_4_GROM,
      O => mac_control_rxf_cnt_n0000(5)
    );
  mac_control_rxf_cnt_4_CYINIT_1518 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_rxf_cnt_4_CYINIT
    );
  mac_control_rxf_cnt_6_LOGIC_ZERO_1519 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_6_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_22_1520 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_6_CYINIT,
      SEL => mac_control_rxf_cnt_6_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_6_CYINIT,
      I1 => mac_control_rxf_cnt_6_FROM,
      O => mac_control_rxf_cnt_n0000(6)
    );
  mac_control_rxf_cnt_6_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(6),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_6_FROM
    );
  mac_control_rxf_cnt_6_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(7),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_6_GROM
    );
  mac_control_rxf_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_6_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_23_1521 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_rxf_cnt_6_GROM,
      O => mac_control_rxf_cnt_6_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_rxf_cnt_6_GROM,
      O => mac_control_rxf_cnt_n0000(7)
    );
  mac_control_rxf_cnt_6_CYINIT_1522 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_rxf_cnt_6_CYINIT
    );
  mac_control_rxf_cnt_8_LOGIC_ZERO_1523 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_8_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_24_1524 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_8_CYINIT,
      SEL => mac_control_rxf_cnt_8_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_8_CYINIT,
      I1 => mac_control_rxf_cnt_8_FROM,
      O => mac_control_rxf_cnt_n0000(8)
    );
  mac_control_rxf_cnt_8_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(8),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_8_FROM
    );
  mac_control_rxf_cnt_8_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(9),
      O => mac_control_rxf_cnt_8_GROM
    );
  mac_control_rxf_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_8_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_25_1525 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_rxf_cnt_8_GROM,
      O => mac_control_rxf_cnt_8_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_rxf_cnt_8_GROM,
      O => mac_control_rxf_cnt_n0000(9)
    );
  mac_control_rxf_cnt_8_CYINIT_1526 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_rxf_cnt_8_CYINIT
    );
  tx_input_dl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(11),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_11_FFX_RST,
      O => tx_input_dl(11)
    );
  tx_input_dl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_11_FFX_RST
    );
  mac_control_rxf_cnt_10_LOGIC_ZERO_1527 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_10_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_26_1528 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_10_CYINIT,
      SEL => mac_control_rxf_cnt_10_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_10_CYINIT,
      I1 => mac_control_rxf_cnt_10_FROM,
      O => mac_control_rxf_cnt_n0000(10)
    );
  mac_control_rxf_cnt_10_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(10),
      O => mac_control_rxf_cnt_10_FROM
    );
  mac_control_rxf_cnt_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(11),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_10_GROM
    );
  mac_control_rxf_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_10_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_27_1529 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_rxf_cnt_10_GROM,
      O => mac_control_rxf_cnt_10_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_rxf_cnt_10_GROM,
      O => mac_control_rxf_cnt_n0000(11)
    );
  mac_control_rxf_cnt_10_CYINIT_1530 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_rxf_cnt_10_CYINIT
    );
  mac_control_rxf_cnt_12_LOGIC_ZERO_1531 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_12_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_28_1532 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_12_CYINIT,
      SEL => mac_control_rxf_cnt_12_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_12_CYINIT,
      I1 => mac_control_rxf_cnt_12_FROM,
      O => mac_control_rxf_cnt_n0000(12)
    );
  mac_control_rxf_cnt_12_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(12),
      O => mac_control_rxf_cnt_12_FROM
    );
  mac_control_rxf_cnt_12_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxf_cnt(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxf_cnt_12_GROM
    );
  mac_control_rxf_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_12_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_29_1533 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_rxf_cnt_12_GROM,
      O => mac_control_rxf_cnt_12_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_rxf_cnt_12_GROM,
      O => mac_control_rxf_cnt_n0000(13)
    );
  mac_control_rxf_cnt_12_CYINIT_1534 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_rxf_cnt_12_CYINIT
    );
  mac_control_rxf_cnt_14_LOGIC_ZERO_1535 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_14_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_30_1536 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_14_CYINIT,
      SEL => mac_control_rxf_cnt_14_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_14_CYINIT,
      I1 => mac_control_rxf_cnt_14_FROM,
      O => mac_control_rxf_cnt_n0000(14)
    );
  mac_control_rxf_cnt_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxf_cnt(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxf_cnt_14_FROM
    );
  mac_control_rxf_cnt_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(15),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_14_GROM
    );
  mac_control_rxf_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_14_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_31_1537 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_rxf_cnt_14_GROM,
      O => mac_control_rxf_cnt_14_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_rxf_cnt_14_GROM,
      O => mac_control_rxf_cnt_n0000(15)
    );
  mac_control_rxf_cnt_14_CYINIT_1538 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_rxf_cnt_14_CYINIT
    );
  mac_control_rxf_cnt_16_LOGIC_ZERO_1539 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_16_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_32_1540 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_16_CYINIT,
      SEL => mac_control_rxf_cnt_16_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_16_CYINIT,
      I1 => mac_control_rxf_cnt_16_FROM,
      O => mac_control_rxf_cnt_n0000(16)
    );
  mac_control_rxf_cnt_16_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(16),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_16_FROM
    );
  mac_control_rxf_cnt_16_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(17),
      O => mac_control_rxf_cnt_16_GROM
    );
  mac_control_rxf_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_16_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_33_1541 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_rxf_cnt_16_GROM,
      O => mac_control_rxf_cnt_16_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_rxf_cnt_16_GROM,
      O => mac_control_rxf_cnt_n0000(17)
    );
  mac_control_rxf_cnt_16_CYINIT_1542 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_rxf_cnt_16_CYINIT
    );
  mac_control_rxf_cnt_18_LOGIC_ZERO_1543 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_18_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_34_1544 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_18_CYINIT,
      SEL => mac_control_rxf_cnt_18_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_18_CYINIT,
      I1 => mac_control_rxf_cnt_18_FROM,
      O => mac_control_rxf_cnt_n0000(18)
    );
  mac_control_rxf_cnt_18_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(18),
      O => mac_control_rxf_cnt_18_FROM
    );
  mac_control_rxf_cnt_18_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(19),
      O => mac_control_rxf_cnt_18_GROM
    );
  mac_control_rxf_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_18_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_35_1545 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_rxf_cnt_18_GROM,
      O => mac_control_rxf_cnt_18_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_rxf_cnt_18_GROM,
      O => mac_control_rxf_cnt_n0000(19)
    );
  mac_control_rxf_cnt_18_CYINIT_1546 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_rxf_cnt_18_CYINIT
    );
  mac_control_rxf_cnt_20_LOGIC_ZERO_1547 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_20_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_36_1548 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_20_CYINIT,
      SEL => mac_control_rxf_cnt_20_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_20_CYINIT,
      I1 => mac_control_rxf_cnt_20_FROM,
      O => mac_control_rxf_cnt_n0000(20)
    );
  mac_control_rxf_cnt_20_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(20),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_20_FROM
    );
  mac_control_rxf_cnt_20_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(21),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxf_cnt_20_GROM
    );
  mac_control_rxf_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_20_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_37_1549 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_rxf_cnt_20_GROM,
      O => mac_control_rxf_cnt_20_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_rxf_cnt_20_GROM,
      O => mac_control_rxf_cnt_n0000(21)
    );
  mac_control_rxf_cnt_20_CYINIT_1550 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_rxf_cnt_20_CYINIT
    );
  mac_control_rxf_cnt_22_LOGIC_ZERO_1551 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_22_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_38_1552 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_22_CYINIT,
      SEL => mac_control_rxf_cnt_22_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_22_CYINIT,
      I1 => mac_control_rxf_cnt_22_FROM,
      O => mac_control_rxf_cnt_n0000(22)
    );
  mac_control_rxf_cnt_22_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(22),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_22_FROM
    );
  mac_control_rxf_cnt_22_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(23),
      O => mac_control_rxf_cnt_22_GROM
    );
  mac_control_rxf_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_22_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_39_1553 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_rxf_cnt_22_GROM,
      O => mac_control_rxf_cnt_22_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_rxf_cnt_22_GROM,
      O => mac_control_rxf_cnt_n0000(23)
    );
  mac_control_rxf_cnt_22_CYINIT_1554 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_rxf_cnt_22_CYINIT
    );
  mac_control_rxf_cnt_24_LOGIC_ZERO_1555 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_24_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_40_1556 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_24_CYINIT,
      SEL => mac_control_rxf_cnt_24_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_24_CYINIT,
      I1 => mac_control_rxf_cnt_24_FROM,
      O => mac_control_rxf_cnt_n0000(24)
    );
  mac_control_rxf_cnt_24_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(24),
      O => mac_control_rxf_cnt_24_FROM
    );
  mac_control_rxf_cnt_24_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(25),
      O => mac_control_rxf_cnt_24_GROM
    );
  mac_control_rxf_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_24_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_41_1557 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_rxf_cnt_24_GROM,
      O => mac_control_rxf_cnt_24_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_rxf_cnt_24_GROM,
      O => mac_control_rxf_cnt_n0000(25)
    );
  mac_control_rxf_cnt_24_CYINIT_1558 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_rxf_cnt_24_CYINIT
    );
  mac_control_rxf_cnt_26_LOGIC_ZERO_1559 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_26_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_42_1560 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_26_CYINIT,
      SEL => mac_control_rxf_cnt_26_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_26_CYINIT,
      I1 => mac_control_rxf_cnt_26_FROM,
      O => mac_control_rxf_cnt_n0000(26)
    );
  mac_control_rxf_cnt_26_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxf_cnt(26),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxf_cnt_26_FROM
    );
  mac_control_rxf_cnt_26_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxf_cnt(27),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxf_cnt_26_GROM
    );
  mac_control_rxf_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_26_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_43_1561 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_rxf_cnt_26_GROM,
      O => mac_control_rxf_cnt_26_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_rxf_cnt_26_GROM,
      O => mac_control_rxf_cnt_n0000(27)
    );
  mac_control_rxf_cnt_26_CYINIT_1562 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_rxf_cnt_26_CYINIT
    );
  mac_control_rxf_cnt_28_LOGIC_ZERO_1563 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_28_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_44_1564 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_28_CYINIT,
      SEL => mac_control_rxf_cnt_28_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_28_CYINIT,
      I1 => mac_control_rxf_cnt_28_FROM,
      O => mac_control_rxf_cnt_n0000(28)
    );
  mac_control_rxf_cnt_28_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(28),
      O => mac_control_rxf_cnt_28_FROM
    );
  mac_control_rxf_cnt_28_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(29),
      O => mac_control_rxf_cnt_28_GROM
    );
  mac_control_rxf_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_28_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_45_1565 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_rxf_cnt_28_GROM,
      O => mac_control_rxf_cnt_28_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_rxf_cnt_28_GROM,
      O => mac_control_rxf_cnt_n0000(29)
    );
  mac_control_rxf_cnt_28_CYINIT_1566 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_rxf_cnt_28_CYINIT
    );
  mac_control_rxf_cnt_30_LOGIC_ZERO_1567 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_30_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_46_1568 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_30_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_30_CYINIT,
      SEL => mac_control_rxf_cnt_30_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_30_CYINIT,
      I1 => mac_control_rxf_cnt_30_FROM,
      O => mac_control_rxf_cnt_n0000(30)
    );
  mac_control_rxf_cnt_30_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(30),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_30_FROM
    );
  mac_control_rxf_cnt_31_rt_1569 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(31),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_31_rt
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_rxf_cnt_31_rt,
      O => mac_control_rxf_cnt_n0000(31)
    );
  mac_control_rxf_cnt_30_CYINIT_1570 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_rxf_cnt_30_CYINIT
    );
  tx_input_bp_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_27,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_11_FFX_RST,
      O => txbp(11)
    );
  txbp_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_11_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_n0078_1_LOGIC_ZERO_1571 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_n0078_1_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_181_1572 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_34,
      IB => mac_control_PHY_status_MII_Interface_n0078_1_LOGIC_ZERO,
      SEL => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_lut2_127,
      O => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_181
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_lut2_1271 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_34,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_lut2_127
    );
  mac_control_PHY_status_MII_Interface_n0078_1_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_15,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(1),
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_n0078_1_GROM
    );
  mac_control_PHY_status_MII_Interface_n0078_1_COUTUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0078_1_CYMUXG,
      O => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_182
    );
  mac_control_PHY_status_MII_Interface_n0078_1_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0078_1_XORG,
      O => mac_control_PHY_status_MII_Interface_n0078(1)
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_182_1573 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_15,
      IB => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_181,
      SEL => mac_control_PHY_status_MII_Interface_n0078_1_GROM,
      O => mac_control_PHY_status_MII_Interface_n0078_1_CYMUXG
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_sum_160 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_181,
      I1 => mac_control_PHY_status_MII_Interface_n0078_1_GROM,
      O => mac_control_PHY_status_MII_Interface_n0078_1_XORG
    );
  mac_control_PHY_status_MII_Interface_n0078_2_LOGIC_ZERO_1574 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_n0078_2_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_183_1575 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_n0078_2_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_n0078_2_CYINIT,
      SEL => mac_control_PHY_status_MII_Interface_n0078_2_FROM,
      O => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_183
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_sum_161 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_n0078_2_CYINIT,
      I1 => mac_control_PHY_status_MII_Interface_n0078_2_FROM,
      O => mac_control_PHY_status_MII_Interface_n0078_2_XORF
    );
  mac_control_PHY_status_MII_Interface_n0078_2_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_n0078_2_FROM
    );
  mac_control_PHY_status_MII_Interface_n0078_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_n0078_2_GROM
    );
  mac_control_PHY_status_MII_Interface_n0078_2_COUTUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0078_2_CYMUXG,
      O => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_184
    );
  mac_control_PHY_status_MII_Interface_n0078_2_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0078_2_XORF,
      O => mac_control_PHY_status_MII_Interface_n0078(2)
    );
  mac_control_PHY_status_MII_Interface_n0078_2_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0078_2_XORG,
      O => mac_control_PHY_status_MII_Interface_n0078(3)
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_184_1576 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_n0078_2_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_183,
      SEL => mac_control_PHY_status_MII_Interface_n0078_2_GROM,
      O => mac_control_PHY_status_MII_Interface_n0078_2_CYMUXG
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_sum_162 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_183,
      I1 => mac_control_PHY_status_MII_Interface_n0078_2_GROM,
      O => mac_control_PHY_status_MII_Interface_n0078_2_XORG
    );
  mac_control_PHY_status_MII_Interface_n0078_2_CYINIT_1577 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_182,
      O => mac_control_PHY_status_MII_Interface_n0078_2_CYINIT
    );
  mac_control_PHY_status_MII_Interface_n0078_4_LOGIC_ZERO_1578 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_n0078_4_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_185_1579 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_n0078_4_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_n0078_4_CYINIT,
      SEL => mac_control_PHY_status_MII_Interface_n0078_4_FROM,
      O => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_185
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_sum_163 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_n0078_4_CYINIT,
      I1 => mac_control_PHY_status_MII_Interface_n0078_4_FROM,
      O => mac_control_PHY_status_MII_Interface_n0078_4_XORF
    );
  mac_control_PHY_status_MII_Interface_n0078_4_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_n0078_4_FROM
    );
  mac_control_PHY_status_MII_Interface_statecnt_5_rt_1580 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(5),
      O => mac_control_PHY_status_MII_Interface_statecnt_5_rt
    );
  mac_control_PHY_status_MII_Interface_n0078_4_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0078_4_XORF,
      O => mac_control_PHY_status_MII_Interface_n0078(4)
    );
  mac_control_PHY_status_MII_Interface_n0078_4_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0078_4_XORG,
      O => mac_control_PHY_status_MII_Interface_n0078(5)
    );
  mac_control_PHY_status_MII_Interface_Madd_n0078_inst_sum_164 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_185,
      I1 => mac_control_PHY_status_MII_Interface_statecnt_5_rt,
      O => mac_control_PHY_status_MII_Interface_n0078_4_XORG
    );
  mac_control_PHY_status_MII_Interface_n0078_4_CYINIT_1581 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_Madd_n0078_inst_cy_184,
      O => mac_control_PHY_status_MII_Interface_n0078_4_CYINIT
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ONE_1582 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ZERO_1583 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_177_1584 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(0),
      ADR1 => rx_input_memio_addrchk_datal(1),
      ADR2 => rx_input_memio_addrchk_macaddrl(0),
      ADR3 => rx_input_memio_addrchk_macaddrl(1),
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(3),
      ADR1 => rx_input_memio_addrchk_macaddrl(2),
      ADR2 => rx_input_memio_addrchk_macaddrl(3),
      ADR3 => rx_input_memio_addrchk_datal(2),
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_1585 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_5_LOGIC_ZERO_1586 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_5_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_179_1587 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_5_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_5_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(4),
      ADR1 => rx_input_memio_addrchk_datal(5),
      ADR2 => rx_input_memio_addrchk_macaddrl(4),
      ADR3 => rx_input_memio_addrchk_macaddrl(5),
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(6),
      ADR1 => rx_input_memio_addrchk_datal(7),
      ADR2 => rx_input_memio_addrchk_macaddrl(7),
      ADR3 => rx_input_memio_addrchk_macaddrl(6),
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_5_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_5_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(5)
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_5_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_5_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_5_CYINIT_1588 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_5_CYINIT
    );
  rx_output_fifo_N9_LOGIC_ZERO_1589 : X_ZERO
    port map (
      O => rx_output_fifo_N9_LOGIC_ZERO
    );
  rx_output_fifo_BU199 : X_MUX2
    port map (
      IA => rx_output_fifo_N9,
      IB => rx_output_fifo_N9_CYINIT,
      SEL => rx_output_fifo_N2840,
      O => rx_output_fifo_N2842
    );
  rx_output_fifo_BU200 : X_XOR2
    port map (
      I0 => rx_output_fifo_N9_CYINIT,
      I1 => rx_output_fifo_N2840,
      O => rx_output_fifo_N2832
    );
  rx_output_fifo_BU198 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_output_fifo_N9,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N2840
    );
  rx_output_fifo_N9_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N8,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N9_GROM
    );
  rx_output_fifo_N9_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N9_CYMUXG,
      O => rx_output_fifo_N2847
    );
  rx_output_fifo_BU205 : X_MUX2
    port map (
      IA => rx_output_fifo_N8,
      IB => rx_output_fifo_N2842,
      SEL => rx_output_fifo_N9_GROM,
      O => rx_output_fifo_N9_CYMUXG
    );
  rx_output_fifo_BU206 : X_XOR2
    port map (
      I0 => rx_output_fifo_N2842,
      I1 => rx_output_fifo_N9_GROM,
      O => rx_output_fifo_N2833
    );
  rx_output_fifo_N9_CYINIT_1590 : X_BUF
    port map (
      I => rx_output_fifo_N9_LOGIC_ZERO,
      O => rx_output_fifo_N9_CYINIT
    );
  rx_output_fifo_BU211 : X_MUX2
    port map (
      IA => rx_output_fifo_N7,
      IB => rx_output_fifo_N7_CYINIT,
      SEL => rx_output_fifo_N7_FROM,
      O => rx_output_fifo_N2852
    );
  rx_output_fifo_BU212 : X_XOR2
    port map (
      I0 => rx_output_fifo_N7_CYINIT,
      I1 => rx_output_fifo_N7_FROM,
      O => rx_output_fifo_N2834
    );
  rx_output_fifo_N7_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N7,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N7_FROM
    );
  rx_output_fifo_N7_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N6,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N7_GROM
    );
  rx_output_fifo_N7_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N7_CYMUXG,
      O => rx_output_fifo_N2857
    );
  rx_output_fifo_BU217 : X_MUX2
    port map (
      IA => rx_output_fifo_N6,
      IB => rx_output_fifo_N2852,
      SEL => rx_output_fifo_N7_GROM,
      O => rx_output_fifo_N7_CYMUXG
    );
  rx_output_fifo_BU218 : X_XOR2
    port map (
      I0 => rx_output_fifo_N2852,
      I1 => rx_output_fifo_N7_GROM,
      O => rx_output_fifo_N2835
    );
  rx_output_fifo_N7_CYINIT_1591 : X_BUF
    port map (
      I => rx_output_fifo_N2847,
      O => rx_output_fifo_N7_CYINIT
    );
  rx_output_fifo_BU223 : X_MUX2
    port map (
      IA => rx_output_fifo_N5,
      IB => rx_output_fifo_N5_CYINIT,
      SEL => rx_output_fifo_N5_FROM,
      O => rx_output_fifo_N2862
    );
  rx_output_fifo_BU224 : X_XOR2
    port map (
      I0 => rx_output_fifo_N5_CYINIT,
      I1 => rx_output_fifo_N5_FROM,
      O => rx_output_fifo_N2836
    );
  rx_output_fifo_N5_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N5,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N5_FROM
    );
  rx_output_fifo_N5_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N4,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N5_GROM
    );
  rx_output_fifo_N5_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N5_CYMUXG,
      O => rx_output_fifo_N2867
    );
  rx_output_fifo_BU229 : X_MUX2
    port map (
      IA => rx_output_fifo_N4,
      IB => rx_output_fifo_N2862,
      SEL => rx_output_fifo_N5_GROM,
      O => rx_output_fifo_N5_CYMUXG
    );
  rx_output_fifo_BU230 : X_XOR2
    port map (
      I0 => rx_output_fifo_N2862,
      I1 => rx_output_fifo_N5_GROM,
      O => rx_output_fifo_N2837
    );
  rx_output_fifo_N5_CYINIT_1592 : X_BUF
    port map (
      I => rx_output_fifo_N2857,
      O => rx_output_fifo_N5_CYINIT
    );
  rx_output_fifo_BU235 : X_MUX2
    port map (
      IA => rx_output_fifo_N3,
      IB => rx_output_fifo_N3_CYINIT,
      SEL => rx_output_fifo_N3_FROM,
      O => rx_output_fifo_N2872
    );
  rx_output_fifo_BU236 : X_XOR2
    port map (
      I0 => rx_output_fifo_N3_CYINIT,
      I1 => rx_output_fifo_N3_FROM,
      O => rx_output_fifo_N2838
    );
  rx_output_fifo_N3_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N3_FROM
    );
  rx_output_fifo_N2_rt_1593 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N2_rt
    );
  rx_output_fifo_BU241 : X_XOR2
    port map (
      I0 => rx_output_fifo_N2872,
      I1 => rx_output_fifo_N2_rt,
      O => rx_output_fifo_N2839
    );
  rx_output_fifo_N3_CYINIT_1594 : X_BUF
    port map (
      I => rx_output_fifo_N2867,
      O => rx_output_fifo_N3_CYINIT
    );
  rx_output_fifo_N2576_LOGIC_ONE_1595 : X_ONE
    port map (
      O => rx_output_fifo_N2576_LOGIC_ONE
    );
  rx_output_fifo_N2576_LOGIC_ZERO_1596 : X_ZERO
    port map (
      O => rx_output_fifo_N2576_LOGIC_ZERO
    );
  rx_output_fifo_BU151 : X_MUX2
    port map (
      IA => rx_output_fifo_N2576_LOGIC_ZERO,
      IB => rx_output_fifo_N2576_LOGIC_ONE,
      SEL => rx_output_fifo_N2569,
      O => rx_output_fifo_N2577
    );
  rx_output_fifo_BU150 : X_LUT4
    generic map(
      INIT => X"E21D"
    )
    port map (
      ADR0 => rx_output_fifo_N1633,
      ADR1 => rx_output_fifo_empty,
      ADR2 => rx_output_fifo_N1617,
      ADR3 => rx_output_fifo_N1553,
      O => rx_output_fifo_N2569
    );
  rx_output_fifo_BU153 : X_LUT4
    generic map(
      INIT => X"B847"
    )
    port map (
      ADR0 => rx_output_fifo_N1616,
      ADR1 => rx_output_fifo_empty,
      ADR2 => rx_output_fifo_N1632,
      ADR3 => rx_output_fifo_N1552,
      O => rx_output_fifo_N2568
    );
  rx_output_fifo_N2576_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N2576_CYMUXG,
      O => rx_output_fifo_N2576
    );
  rx_output_fifo_BU154 : X_MUX2
    port map (
      IA => rx_output_fifo_N2576_LOGIC_ZERO,
      IB => rx_output_fifo_N2577,
      SEL => rx_output_fifo_N2568,
      O => rx_output_fifo_N2576_CYMUXG
    );
  rx_output_fifo_N2574_LOGIC_ZERO_1597 : X_ZERO
    port map (
      O => rx_output_fifo_N2574_LOGIC_ZERO
    );
  rx_output_fifo_BU157 : X_MUX2
    port map (
      IA => rx_output_fifo_N2574_LOGIC_ZERO,
      IB => rx_output_fifo_N2574_CYINIT,
      SEL => rx_output_fifo_N2567,
      O => rx_output_fifo_N2575
    );
  rx_output_fifo_BU156 : X_LUT4
    generic map(
      INIT => X"C3A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1631,
      ADR1 => rx_output_fifo_N1615,
      ADR2 => rx_output_fifo_N1551,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N2567
    );
  rx_output_fifo_BU159 : X_LUT4
    generic map(
      INIT => X"99A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1550,
      ADR1 => rx_output_fifo_N1614,
      ADR2 => rx_output_fifo_N1630,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N2566
    );
  rx_output_fifo_N2574_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N2574_CYMUXG,
      O => rx_output_fifo_N2574
    );
  rx_output_fifo_BU160 : X_MUX2
    port map (
      IA => rx_output_fifo_N2574_LOGIC_ZERO,
      IB => rx_output_fifo_N2575,
      SEL => rx_output_fifo_N2566,
      O => rx_output_fifo_N2574_CYMUXG
    );
  rx_output_fifo_N2574_CYINIT_1598 : X_BUF
    port map (
      I => rx_output_fifo_N2576,
      O => rx_output_fifo_N2574_CYINIT
    );
  tx_input_dl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(13),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_13_FFX_RST,
      O => tx_input_dl(13)
    );
  tx_input_dl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_13_FFX_RST
    );
  rx_output_fifo_N2572_LOGIC_ZERO_1599 : X_ZERO
    port map (
      O => rx_output_fifo_N2572_LOGIC_ZERO
    );
  rx_output_fifo_BU163 : X_MUX2
    port map (
      IA => rx_output_fifo_N2572_LOGIC_ZERO,
      IB => rx_output_fifo_N2572_CYINIT,
      SEL => rx_output_fifo_N2565,
      O => rx_output_fifo_N2573
    );
  rx_output_fifo_BU162 : X_LUT4
    generic map(
      INIT => X"CA35"
    )
    port map (
      ADR0 => rx_output_fifo_N1629,
      ADR1 => rx_output_fifo_N1613,
      ADR2 => rx_output_fifo_empty,
      ADR3 => rx_output_fifo_N1549,
      O => rx_output_fifo_N2565
    );
  rx_output_fifo_BU165 : X_LUT4
    generic map(
      INIT => X"99A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1548,
      ADR1 => rx_output_fifo_N1612,
      ADR2 => rx_output_fifo_N1628,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N2564
    );
  rx_output_fifo_N2572_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N2572_CYMUXG,
      O => rx_output_fifo_N2572
    );
  rx_output_fifo_BU166 : X_MUX2
    port map (
      IA => rx_output_fifo_N2572_LOGIC_ZERO,
      IB => rx_output_fifo_N2573,
      SEL => rx_output_fifo_N2564,
      O => rx_output_fifo_N2572_CYMUXG
    );
  rx_output_fifo_N2572_CYINIT_1600 : X_BUF
    port map (
      I => rx_output_fifo_N2574,
      O => rx_output_fifo_N2572_CYINIT
    );
  rx_output_fifo_BU172_O_LOGIC_ZERO_1601 : X_ZERO
    port map (
      O => rx_output_fifo_BU172_O_LOGIC_ZERO
    );
  rx_output_fifo_BU169 : X_MUX2
    port map (
      IA => rx_output_fifo_BU172_O_LOGIC_ZERO,
      IB => rx_output_fifo_BU172_O_CYINIT,
      SEL => rx_output_fifo_N2563,
      O => rx_output_fifo_N2571
    );
  rx_output_fifo_BU168 : X_LUT4
    generic map(
      INIT => X"D827"
    )
    port map (
      ADR0 => rx_output_fifo_empty,
      ADR1 => rx_output_fifo_N1611,
      ADR2 => rx_output_fifo_N1627,
      ADR3 => rx_output_fifo_N1547,
      O => rx_output_fifo_N2563
    );
  rx_output_fifo_BU171 : X_LUT4
    generic map(
      INIT => X"A599"
    )
    port map (
      ADR0 => rx_output_fifo_N1546,
      ADR1 => rx_output_fifo_N1626,
      ADR2 => rx_output_fifo_N1610,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N2562
    );
  rx_output_fifo_BU172_O_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_BU172_O_CYMUXG,
      O => rx_output_fifo_BU172_O
    );
  rx_output_fifo_BU172 : X_MUX2
    port map (
      IA => rx_output_fifo_BU172_O_LOGIC_ZERO,
      IB => rx_output_fifo_N2571,
      SEL => rx_output_fifo_N2562,
      O => rx_output_fifo_BU172_O_CYMUXG
    );
  rx_output_fifo_BU172_O_CYINIT_1602 : X_BUF
    port map (
      I => rx_output_fifo_N2572,
      O => rx_output_fifo_BU172_O_CYINIT
    );
  rx_output_fifo_BU175 : X_XOR2
    port map (
      I0 => rx_output_fifo_empty_CYINIT,
      I1 => rx_output_fifo_empty_FROM,
      O => rx_output_fifo_N2580
    );
  rx_output_fifo_empty_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_empty_FROM
    );
  rx_output_fifo_empty_CYINIT_1603 : X_BUF
    port map (
      I => rx_output_fifo_BU172_O,
      O => rx_output_fifo_empty_CYINIT
    );
  rx_output_fifo_N3614_LOGIC_ONE_1604 : X_ONE
    port map (
      O => rx_output_fifo_N3614_LOGIC_ONE
    );
  rx_output_fifo_N3614_LOGIC_ZERO_1605 : X_ZERO
    port map (
      O => rx_output_fifo_N3614_LOGIC_ZERO
    );
  rx_output_fifo_BU330 : X_MUX2
    port map (
      IA => rx_output_fifo_N3614_LOGIC_ZERO,
      IB => rx_output_fifo_N3614_LOGIC_ONE,
      SEL => rx_output_fifo_N3607,
      O => rx_output_fifo_N3615
    );
  rx_output_fifo_BU329 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => rx_output_fifo_N1577,
      ADR1 => rx_output_fifo_N1617,
      ADR2 => rx_output_fifo_N1569,
      ADR3 => rx_output_fifo_full_0,
      O => rx_output_fifo_N3607
    );
  rx_output_fifo_BU332 : X_LUT4
    generic map(
      INIT => X"D827"
    )
    port map (
      ADR0 => rx_output_fifo_full_0,
      ADR1 => rx_output_fifo_N1568,
      ADR2 => rx_output_fifo_N1576,
      ADR3 => rx_output_fifo_N1616,
      O => rx_output_fifo_N3606
    );
  rx_output_fifo_N3614_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N3614_CYMUXG,
      O => rx_output_fifo_N3614
    );
  rx_output_fifo_BU333 : X_MUX2
    port map (
      IA => rx_output_fifo_N3614_LOGIC_ZERO,
      IB => rx_output_fifo_N3615,
      SEL => rx_output_fifo_N3606,
      O => rx_output_fifo_N3614_CYMUXG
    );
  rx_output_fifo_N3612_LOGIC_ZERO_1606 : X_ZERO
    port map (
      O => rx_output_fifo_N3612_LOGIC_ZERO
    );
  rx_output_fifo_BU336 : X_MUX2
    port map (
      IA => rx_output_fifo_N3612_LOGIC_ZERO,
      IB => rx_output_fifo_N3612_CYINIT,
      SEL => rx_output_fifo_N3605,
      O => rx_output_fifo_N3613
    );
  rx_output_fifo_BU335 : X_LUT4
    generic map(
      INIT => X"E12D"
    )
    port map (
      ADR0 => rx_output_fifo_N1575,
      ADR1 => rx_output_fifo_full_0,
      ADR2 => rx_output_fifo_N1615,
      ADR3 => rx_output_fifo_N1567,
      O => rx_output_fifo_N3605
    );
  rx_output_fifo_BU338 : X_LUT4
    generic map(
      INIT => X"CA35"
    )
    port map (
      ADR0 => rx_output_fifo_N1574,
      ADR1 => rx_output_fifo_N1566,
      ADR2 => rx_output_fifo_full_0,
      ADR3 => rx_output_fifo_N1614,
      O => rx_output_fifo_N3604
    );
  rx_output_fifo_N3612_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N3612_CYMUXG,
      O => rx_output_fifo_N3612
    );
  rx_output_fifo_BU339 : X_MUX2
    port map (
      IA => rx_output_fifo_N3612_LOGIC_ZERO,
      IB => rx_output_fifo_N3613,
      SEL => rx_output_fifo_N3604,
      O => rx_output_fifo_N3612_CYMUXG
    );
  rx_output_fifo_N3612_CYINIT_1607 : X_BUF
    port map (
      I => rx_output_fifo_N3614,
      O => rx_output_fifo_N3612_CYINIT
    );
  rx_output_fifo_N3610_LOGIC_ZERO_1608 : X_ZERO
    port map (
      O => rx_output_fifo_N3610_LOGIC_ZERO
    );
  rx_output_fifo_BU342 : X_MUX2
    port map (
      IA => rx_output_fifo_N3610_LOGIC_ZERO,
      IB => rx_output_fifo_N3610_CYINIT,
      SEL => rx_output_fifo_N3603,
      O => rx_output_fifo_N3611
    );
  rx_output_fifo_BU341 : X_LUT4
    generic map(
      INIT => X"E21D"
    )
    port map (
      ADR0 => rx_output_fifo_N1573,
      ADR1 => rx_output_fifo_full_0,
      ADR2 => rx_output_fifo_N1565,
      ADR3 => rx_output_fifo_N1613,
      O => rx_output_fifo_N3603
    );
  rx_output_fifo_BU344 : X_LUT4
    generic map(
      INIT => X"A695"
    )
    port map (
      ADR0 => rx_output_fifo_N1612,
      ADR1 => rx_output_fifo_full_0,
      ADR2 => rx_output_fifo_N1564,
      ADR3 => rx_output_fifo_N1572,
      O => rx_output_fifo_N3602
    );
  rx_output_fifo_N3610_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N3610_CYMUXG,
      O => rx_output_fifo_N3610
    );
  rx_output_fifo_BU345 : X_MUX2
    port map (
      IA => rx_output_fifo_N3610_LOGIC_ZERO,
      IB => rx_output_fifo_N3611,
      SEL => rx_output_fifo_N3602,
      O => rx_output_fifo_N3610_CYMUXG
    );
  rx_output_fifo_N3610_CYINIT_1609 : X_BUF
    port map (
      I => rx_output_fifo_N3612,
      O => rx_output_fifo_N3610_CYINIT
    );
  rx_output_fifo_BU351_O_LOGIC_ZERO_1610 : X_ZERO
    port map (
      O => rx_output_fifo_BU351_O_LOGIC_ZERO
    );
  rx_output_fifo_BU348 : X_MUX2
    port map (
      IA => rx_output_fifo_BU351_O_LOGIC_ZERO,
      IB => rx_output_fifo_BU351_O_CYINIT,
      SEL => rx_output_fifo_N3601,
      O => rx_output_fifo_N3609
    );
  rx_output_fifo_BU347 : X_LUT4
    generic map(
      INIT => X"E21D"
    )
    port map (
      ADR0 => rx_output_fifo_N1571,
      ADR1 => rx_output_fifo_full_0,
      ADR2 => rx_output_fifo_N1563,
      ADR3 => rx_output_fifo_N1611,
      O => rx_output_fifo_N3601
    );
  rx_output_fifo_BU350 : X_LUT4
    generic map(
      INIT => X"E21D"
    )
    port map (
      ADR0 => rx_output_fifo_N1570,
      ADR1 => rx_output_fifo_full_0,
      ADR2 => rx_output_fifo_N1562,
      ADR3 => rx_output_fifo_N1610,
      O => rx_output_fifo_N3600
    );
  rx_output_fifo_BU351_O_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_BU351_O_CYMUXG,
      O => rx_output_fifo_BU351_O
    );
  rx_output_fifo_BU351 : X_MUX2
    port map (
      IA => rx_output_fifo_BU351_O_LOGIC_ZERO,
      IB => rx_output_fifo_N3609,
      SEL => rx_output_fifo_N3600,
      O => rx_output_fifo_BU351_O_CYMUXG
    );
  rx_output_fifo_BU351_O_CYINIT_1611 : X_BUF
    port map (
      I => rx_output_fifo_N3610,
      O => rx_output_fifo_BU351_O_CYINIT
    );
  tx_input_dl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(14),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_15_FFY_RST,
      O => tx_input_dl(14)
    );
  tx_input_dl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_15_FFY_RST
    );
  rx_output_fifo_BU354 : X_XOR2
    port map (
      I0 => rx_output_fifo_full_CYINIT,
      I1 => rx_output_fifo_full_FROM,
      O => rx_output_fifo_N3618
    );
  rx_output_fifo_full_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_full_FROM
    );
  rx_output_fifo_full_CYINIT_1612 : X_BUF
    port map (
      I => rx_output_fifo_BU351_O,
      O => rx_output_fifo_full_CYINIT
    );
  rx_output_fifo_N4763_LOGIC_ONE_1613 : X_ONE
    port map (
      O => rx_output_fifo_N4763_LOGIC_ONE
    );
  rx_output_fifo_BU477 : X_MUX2
    port map (
      IA => rx_output_fifo_N1609,
      IB => rx_output_fifo_N4763_LOGIC_ONE,
      SEL => rx_output_fifo_N4756,
      O => rx_output_fifo_N4759
    );
  rx_output_fifo_BU476 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1609,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N1593,
      ADR3 => VCC,
      O => rx_output_fifo_N4756
    );
  rx_output_fifo_BU479 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_output_fifo_N1608,
      ADR1 => rx_output_fifo_N1592,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N4760
    );
  rx_output_fifo_N4763_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N4763_CYMUXG,
      O => rx_output_fifo_N4763
    );
  rx_output_fifo_BU480 : X_MUX2
    port map (
      IA => rx_output_fifo_N1608,
      IB => rx_output_fifo_N4759,
      SEL => rx_output_fifo_N4760,
      O => rx_output_fifo_N4763_CYMUXG
    );
  rx_output_fifo_BU483 : X_MUX2
    port map (
      IA => rx_output_fifo_N1607,
      IB => rx_output_fifo_N4771_CYINIT,
      SEL => rx_output_fifo_N4764,
      O => rx_output_fifo_N4767
    );
  rx_output_fifo_BU482 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_output_fifo_N1607,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N1591,
      O => rx_output_fifo_N4764
    );
  rx_output_fifo_BU485 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_output_fifo_N1606,
      ADR1 => rx_output_fifo_N1590,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N4768
    );
  rx_output_fifo_N4771_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N4771_CYMUXG,
      O => rx_output_fifo_N4771
    );
  rx_output_fifo_BU486 : X_MUX2
    port map (
      IA => rx_output_fifo_N1606,
      IB => rx_output_fifo_N4767,
      SEL => rx_output_fifo_N4768,
      O => rx_output_fifo_N4771_CYMUXG
    );
  rx_output_fifo_N4771_CYINIT_1614 : X_BUF
    port map (
      I => rx_output_fifo_N4763,
      O => rx_output_fifo_N4771_CYINIT
    );
  rx_output_fifo_BU489 : X_MUX2
    port map (
      IA => rx_output_fifo_N1605,
      IB => rx_output_fifo_N4779_CYINIT,
      SEL => rx_output_fifo_N4772,
      O => rx_output_fifo_N4775
    );
  rx_output_fifo_BU488 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_output_fifo_N1605,
      ADR1 => rx_output_fifo_N1589,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N4772
    );
  rx_output_fifo_BU491 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_output_fifo_N1604,
      ADR1 => rx_output_fifo_N1588,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N4776
    );
  rx_output_fifo_N4779_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N4779_CYMUXG,
      O => rx_output_fifo_N4779
    );
  rx_output_fifo_BU492 : X_MUX2
    port map (
      IA => rx_output_fifo_N1604,
      IB => rx_output_fifo_N4775,
      SEL => rx_output_fifo_N4776,
      O => rx_output_fifo_N4779_CYMUXG
    );
  rx_output_fifo_N4779_CYINIT_1615 : X_BUF
    port map (
      I => rx_output_fifo_N4771,
      O => rx_output_fifo_N4779_CYINIT
    );
  tx_input_bp_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_29,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_13_FFX_RST,
      O => txbp(13)
    );
  txbp_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_13_FFX_RST
    );
  rx_output_fifo_BU495 : X_MUX2
    port map (
      IA => rx_output_fifo_N1603,
      IB => rx_output_fifo_wrcount_0_CYINIT,
      SEL => rx_output_fifo_N4780,
      O => rx_output_fifo_N4783
    );
  rx_output_fifo_BU496 : X_XOR2
    port map (
      I0 => rx_output_fifo_wrcount_0_CYINIT,
      I1 => rx_output_fifo_N4780,
      O => rx_output_fifo_N4754
    );
  rx_output_fifo_BU494 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_output_fifo_N1603,
      ADR1 => rx_output_fifo_N1587,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N4780
    );
  rx_output_fifo_BU500 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_output_fifo_N1602,
      ADR1 => rx_output_fifo_N1586,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N4786
    );
  rx_output_fifo_BU502 : X_XOR2
    port map (
      I0 => rx_output_fifo_N4783,
      I1 => rx_output_fifo_N4786,
      O => rx_output_fifo_N4755
    );
  rx_output_fifo_wrcount_0_CYINIT_1616 : X_BUF
    port map (
      I => rx_output_fifo_N4779,
      O => rx_output_fifo_wrcount_0_CYINIT
    );
  mac_control_bitcnt_104_LOGIC_ZERO_1617 : X_ZERO
    port map (
      O => mac_control_bitcnt_104_LOGIC_ZERO
    );
  mac_control_bitcnt_inst_cy_287_1618 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_20,
      IB => mac_control_bitcnt_104_LOGIC_ZERO,
      SEL => mac_control_Mshreg_scslll_103_rt,
      O => mac_control_bitcnt_inst_cy_287
    );
  mac_control_Mshreg_scslll_103_rt_1619 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_20,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_Mshreg_scslll_103,
      O => mac_control_Mshreg_scslll_103_rt
    );
  mac_control_bitcnt_inst_lut3_1861 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_4,
      ADR1 => VCC,
      ADR2 => mac_control_Mshreg_scslll_103,
      ADR3 => mac_control_bitcnt_104,
      O => mac_control_bitcnt_inst_lut3_186
    );
  mac_control_bitcnt_104_COUTUSED : X_BUF
    port map (
      I => mac_control_bitcnt_104_CYMUXG,
      O => mac_control_bitcnt_inst_cy_288
    );
  mac_control_bitcnt_inst_cy_288_1620 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_4,
      IB => mac_control_bitcnt_inst_cy_287,
      SEL => mac_control_bitcnt_inst_lut3_186,
      O => mac_control_bitcnt_104_CYMUXG
    );
  mac_control_bitcnt_inst_sum_251_1621 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_inst_cy_287,
      I1 => mac_control_bitcnt_inst_lut3_186,
      O => mac_control_bitcnt_inst_sum_251
    );
  mac_control_bitcnt_105_LOGIC_ZERO_1622 : X_ZERO
    port map (
      O => mac_control_bitcnt_105_LOGIC_ZERO
    );
  mac_control_bitcnt_inst_cy_289_1623 : X_MUX2
    port map (
      IA => mac_control_bitcnt_105_LOGIC_ZERO,
      IB => mac_control_bitcnt_105_CYINIT,
      SEL => mac_control_bitcnt_inst_lut3_187,
      O => mac_control_bitcnt_inst_cy_289
    );
  mac_control_bitcnt_inst_sum_252_1624 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_105_CYINIT,
      I1 => mac_control_bitcnt_inst_lut3_187,
      O => mac_control_bitcnt_inst_sum_252
    );
  mac_control_bitcnt_inst_lut3_1871 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_bitcnt_105,
      ADR2 => mac_control_Mshreg_scslll_103,
      ADR3 => VCC,
      O => mac_control_bitcnt_inst_lut3_187
    );
  mac_control_bitcnt_inst_lut3_1881 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_Mshreg_scslll_103,
      ADR2 => VCC,
      ADR3 => mac_control_bitcnt_106,
      O => mac_control_bitcnt_inst_lut3_188
    );
  mac_control_bitcnt_105_COUTUSED : X_BUF
    port map (
      I => mac_control_bitcnt_105_CYMUXG,
      O => mac_control_bitcnt_inst_cy_290
    );
  mac_control_bitcnt_inst_cy_290_1625 : X_MUX2
    port map (
      IA => mac_control_bitcnt_105_LOGIC_ZERO,
      IB => mac_control_bitcnt_inst_cy_289,
      SEL => mac_control_bitcnt_inst_lut3_188,
      O => mac_control_bitcnt_105_CYMUXG
    );
  mac_control_bitcnt_inst_sum_253_1626 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_inst_cy_289,
      I1 => mac_control_bitcnt_inst_lut3_188,
      O => mac_control_bitcnt_inst_sum_253
    );
  mac_control_bitcnt_105_CYINIT_1627 : X_BUF
    port map (
      I => mac_control_bitcnt_inst_cy_288,
      O => mac_control_bitcnt_105_CYINIT
    );
  mac_control_bitcnt_107_LOGIC_ZERO_1628 : X_ZERO
    port map (
      O => mac_control_bitcnt_107_LOGIC_ZERO
    );
  mac_control_bitcnt_inst_cy_291_1629 : X_MUX2
    port map (
      IA => mac_control_bitcnt_107_LOGIC_ZERO,
      IB => mac_control_bitcnt_107_CYINIT,
      SEL => mac_control_bitcnt_inst_lut3_189,
      O => mac_control_bitcnt_inst_cy_291
    );
  mac_control_bitcnt_inst_sum_254_1630 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_107_CYINIT,
      I1 => mac_control_bitcnt_inst_lut3_189,
      O => mac_control_bitcnt_inst_sum_254
    );
  mac_control_bitcnt_inst_lut3_1891 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_Mshreg_scslll_103,
      ADR3 => mac_control_bitcnt_107,
      O => mac_control_bitcnt_inst_lut3_189
    );
  mac_control_bitcnt_inst_lut3_1901 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_Mshreg_scslll_103,
      ADR2 => mac_control_bitcnt_108,
      ADR3 => VCC,
      O => mac_control_bitcnt_inst_lut3_190
    );
  mac_control_bitcnt_107_COUTUSED : X_BUF
    port map (
      I => mac_control_bitcnt_107_CYMUXG,
      O => mac_control_bitcnt_inst_cy_292
    );
  mac_control_bitcnt_inst_cy_292_1631 : X_MUX2
    port map (
      IA => mac_control_bitcnt_107_LOGIC_ZERO,
      IB => mac_control_bitcnt_inst_cy_291,
      SEL => mac_control_bitcnt_inst_lut3_190,
      O => mac_control_bitcnt_107_CYMUXG
    );
  mac_control_bitcnt_inst_sum_255_1632 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_inst_cy_291,
      I1 => mac_control_bitcnt_inst_lut3_190,
      O => mac_control_bitcnt_inst_sum_255
    );
  mac_control_bitcnt_107_CYINIT_1633 : X_BUF
    port map (
      I => mac_control_bitcnt_inst_cy_290,
      O => mac_control_bitcnt_107_CYINIT
    );
  tx_output_cs_Out101 : X_LUT4
    generic map(
      INIT => X"0003"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd2,
      ADR2 => tx_output_cs_FFd7,
      ADR3 => tx_output_cs_FFd3,
      O => tx_output_crcsel(0)
    );
  tx_output_crcsell_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_crcsell_1_CEMUXNOT
    );
  mac_control_n00631 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_din(1),
      ADR1 => mac_control_newcmd,
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_N52236,
      O => mac_control_n0063
    );
  mac_control_n00641 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_newcmd,
      ADR1 => mac_control_din(2),
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_N52236,
      O => mac_control_n0064
    );
  rx_input_memio_addrchk_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"3210"
    )
    port map (
      ADR0 => rx_input_memio_brdy,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => rx_input_memio_addrchk_cs_FFd4,
      ADR3 => rx_input_memio_addrchk_cs_FFd5,
      O => rx_input_memio_addrchk_cs_FFd4_In
    );
  rx_input_memio_addrchk_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"0E04"
    )
    port map (
      ADR0 => rx_input_memio_brdy,
      ADR1 => rx_input_memio_addrchk_cs_FFd3,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => rx_input_memio_addrchk_cs_FFd4,
      O => rx_input_memio_addrchk_cs_FFd3_In
    );
  rx_input_memio_cs_FFd10_In1 : X_LUT4
    generic map(
      INIT => X"AE04"
    )
    port map (
      ADR0 => rx_input_invalid,
      ADR1 => rx_input_memio_cs_FFd12,
      ADR2 => rx_input_endf,
      ADR3 => rx_input_memio_cs_FFd10,
      O => rx_input_memio_cs_FFd10_In
    );
  rx_input_memio_cs_FFd9_In1 : X_LUT4
    generic map(
      INIT => X"DCCC"
    )
    port map (
      ADR0 => rx_input_invalid,
      ADR1 => rx_input_memio_cs_FFd11,
      ADR2 => rx_input_memio_cs_FFd12,
      ADR3 => rx_input_endf,
      O => rx_input_memio_cs_FFd9_In
    );
  mac_control_PHY_status_MII_Interface_n0014_3_1 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_n0079,
      ADR1 => mac_control_PHY_status_MII_Interface_n0078(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_n0014(3)
    );
  mac_control_PHY_status_MII_Interface_n0014_2_1 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_n0078(2),
      ADR1 => mac_control_PHY_status_MII_Interface_n0079,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_n0014(2)
    );
  mac_control_PHY_status_MII_Interface_n0014_5_1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_n0079,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_n0078(5),
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_n0014(5)
    );
  mac_control_PHY_status_MII_Interface_n0014_4_1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_n0079,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_n0078(4),
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_n0014(4)
    );
  rx_input_memio_Mmux_lma_Result_1_1 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => rx_input_memio_macnt_71,
      ADR1 => rx_input_memio_wbpl,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bpl(1),
      O => rx_input_memio_lma(1)
    );
  rx_input_memio_Mmux_lma_Result_0_1 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bpl(0),
      ADR3 => rx_input_memio_macnt_70,
      O => rx_input_memio_lma(0)
    );
  tx_input_dl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(15),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_15_FFX_RST,
      O => tx_input_dl(15)
    );
  tx_input_dl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_15_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd3_In_1634 : X_LUT4
    generic map(
      INIT => X"5073"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_n0004,
      ADR1 => mac_control_PHY_status_MII_Interface_N69539,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd3,
      ADR3 => mac_control_PHY_status_MII_Interface_mdccnt_37,
      O => mac_control_PHY_status_MII_Interface_cs_FFd3_In
    );
  rx_input_memio_Mmux_lma_Result_3_1 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_macnt_73,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bpl(3),
      O => rx_input_memio_lma(3)
    );
  rx_input_memio_Mmux_lma_Result_2_1 : X_LUT4
    generic map(
      INIT => X"F3C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_wbpl,
      ADR2 => rx_input_memio_bpl(2),
      ADR3 => rx_input_memio_macnt_72,
      O => rx_input_memio_lma(2)
    );
  mac_control_PHY_status_MII_Interface_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"AAA8"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd6,
      ADR1 => mac_control_PHY_status_cs_FFd3,
      ADR2 => mac_control_PHY_status_cs_FFd6,
      ADR3 => mac_control_PHY_status_cs_FFd8,
      O => mac_control_PHY_status_MII_Interface_cs_FFd5_In
    );
  mac_control_PHY_status_MII_Interface_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"FABA"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => MDC_OBUF,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd4,
      ADR3 => mac_control_PHY_status_MII_Interface_mdccnt_37,
      O => mac_control_PHY_status_MII_Interface_cs_FFd4_In
    );
  rx_input_memio_Mmux_lma_Result_5_1 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bpl(5),
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_75,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(5)
    );
  rx_input_memio_Mmux_lma_Result_4_1 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bpl(4),
      ADR3 => rx_input_memio_macnt_74,
      O => rx_input_memio_lma(4)
    );
  rx_input_memio_Mmux_lma_Result_7_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_bpl(7),
      ADR2 => VCC,
      ADR3 => rx_input_memio_macnt_77,
      O => rx_input_memio_lma(7)
    );
  rx_input_memio_Mmux_lma_Result_6_1 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_macnt_76,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bpl(6),
      O => rx_input_memio_lma(6)
    );
  rx_input_memio_Mmux_lma_Result_9_1 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => rx_input_memio_bpl(9),
      ADR1 => rx_input_memio_macnt_79,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lma(9)
    );
  rx_input_memio_Mmux_lma_Result_8_1 : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => rx_input_memio_macnt_78,
      ADR1 => rx_input_memio_bpl(8),
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lma(8)
    );
  rx_input_memio_Mmux_lmd_Result_1_1 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(1),
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(1),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(1)
    );
  rx_input_memio_Mmux_lmd_Result_0_1 : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => rx_input_memio_doutl(0),
      ADR1 => rx_input_memio_bcntl(0),
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lmd(0)
    );
  rx_input_memio_Mmux_lmd_Result_3_1 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_wbpl,
      ADR2 => rx_input_memio_doutl(3),
      ADR3 => rx_input_memio_bcntl(3),
      O => rx_input_memio_lmd(3)
    );
  rx_input_memio_Mmux_lmd_Result_2_1 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcntl(2),
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_doutl(2),
      O => rx_input_memio_lmd(2)
    );
  rx_input_memio_Mmux_lmd_Result_5_1 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => rx_input_memio_doutl(5),
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcntl(5),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(5)
    );
  rx_input_memio_Mmux_lmd_Result_4_1 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(4),
      ADR1 => rx_input_memio_wbpl,
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(4),
      O => rx_input_memio_lmd(4)
    );
  rx_input_memio_Mmux_lmd_Result_7_1 : X_LUT4
    generic map(
      INIT => X"B8B8"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(7),
      ADR1 => rx_input_memio_wbpl,
      ADR2 => rx_input_memio_doutl(7),
      ADR3 => VCC,
      O => rx_input_memio_lmd(7)
    );
  rx_input_memio_Mmux_lmd_Result_6_1 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcntl(6),
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_doutl(6),
      O => rx_input_memio_lmd(6)
    );
  rx_input_memio_Mmux_lmd_Result_9_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_bcntl(9),
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(9),
      O => rx_input_memio_lmd(9)
    );
  rx_input_memio_Mmux_lmd_Result_8_1 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => rx_input_memio_doutl(8),
      ADR1 => rx_input_memio_wbpl,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bcntl(8),
      O => rx_input_memio_lmd(8)
    );
  tx_input_bp_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_31,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_15_FFX_RST,
      O => txbp(15)
    );
  txbp_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_15_FFX_RST
    );
  rx_input_memio_n0048_21_1 : X_LUT4
    generic map(
      INIT => X"F9F6"
    )
    port map (
      ADR0 => rx_input_memio_crcl(29),
      ADR1 => rx_input_memio_datal(2),
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crcl(13),
      O => rx_input_memio_n0048(21)
    );
  rx_input_memio_n0048_20_1 : X_LUT4
    generic map(
      INIT => X"F9F6"
    )
    port map (
      ADR0 => rx_input_memio_crcl(12),
      ADR1 => rx_input_memio_crcl(28),
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_datal(3),
      O => rx_input_memio_n0048(20)
    );
  rx_input_memio_addrchk_cs_FFd1_1635 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd1_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd1_FFY_RST,
      O => rx_input_memio_addrchk_cs_FFd1
    );
  rx_input_memio_addrchk_cs_FFd1_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd1_FFY_RST
    );
  rx_input_memio_crcl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_31_FFY_RST
    );
  rx_input_memio_crcl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(22),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_31_FFY_RST,
      O => rx_input_memio_crcl(22)
    );
  rx_input_memio_n0048_31_1 : X_LUT4
    generic map(
      INIT => X"FF96"
    )
    port map (
      ADR0 => rx_input_memio_crcl(23),
      ADR1 => rx_input_memio_crcl(29),
      ADR2 => rx_input_memio_datal(2),
      ADR3 => rx_input_memio_crcrst,
      O => rx_input_memio_n0048(31)
    );
  rx_input_memio_n0048_22_1 : X_LUT4
    generic map(
      INIT => X"EDDE"
    )
    port map (
      ADR0 => rx_input_memio_crcl(24),
      ADR1 => rx_input_memio_crcrst,
      ADR2 => rx_input_memio_crcl(14),
      ADR3 => rx_input_memio_datal(7),
      O => rx_input_memio_n0048(22)
    );
  rx_input_memio_cs_FFd12_In1 : X_LUT4
    generic map(
      INIT => X"DC10"
    )
    port map (
      ADR0 => rx_input_endf,
      ADR1 => rx_input_invalid,
      ADR2 => rx_input_memio_cs_FFd14,
      ADR3 => rx_input_memio_cs_FFd12,
      O => rx_input_memio_cs_FFd12_In
    );
  rx_input_memio_cs_FFd11_In1 : X_LUT4
    generic map(
      INIT => X"5000"
    )
    port map (
      ADR0 => rx_input_invalid,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd14,
      ADR3 => rx_input_endf,
      O => rx_input_memio_cs_FFd11_In
    );
  rx_input_memio_cs_FFd14_In1 : X_LUT4
    generic map(
      INIT => X"F022"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd15,
      ADR1 => rx_input_endf,
      ADR2 => rx_input_memio_cs_FFd14,
      ADR3 => rx_input_invalid,
      O => rx_input_memio_cs_FFd14_In
    );
  rx_input_memio_cs_FFd13_In1 : X_LUT4
    generic map(
      INIT => X"CCEC"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd15,
      ADR1 => rx_input_memio_cs_FFd8,
      ADR2 => rx_input_endf,
      ADR3 => rx_input_invalid,
      O => rx_input_memio_cs_FFd13_In
    );
  mac_control_n00651 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_din(3),
      ADR1 => mac_control_N52236,
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_newcmd,
      O => mac_control_n0065
    );
  mac_control_n00671 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_N52236,
      ADR1 => mac_control_N52118,
      ADR2 => mac_control_din(5),
      ADR3 => mac_control_newcmd,
      O => mac_control_n0067
    );
  rx_input_memio_cs_Out916 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_Out916_SW0_2,
      ADR2 => rx_input_memio_cs_Out916_2,
      ADR3 => rx_input_memio_CHOICE1570,
      O => rx_input_memio_menl_FROM
    );
  rx_input_memio_n01011 : X_LUT4
    generic map(
      INIT => X"F5F0"
    )
    port map (
      ADR0 => rx_input_memio_menl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => rx_input_memio_men,
      O => rx_input_memio_menl_GROM
    );
  rx_input_memio_menl_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_menl_CEMUXNOT
    );
  rx_input_memio_menl_XUSED : X_BUF
    port map (
      I => rx_input_memio_menl_FROM,
      O => rx_input_memio_men
    );
  rx_input_memio_menl_YUSED : X_BUF
    port map (
      I => rx_input_memio_menl_GROM,
      O => rx_input_memio_n0101
    );
  rx_input_memio_Mmux_lma_Result_11_1 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => rx_input_memio_macnt_81,
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_bpl(11),
      O => rx_input_memio_lma(11)
    );
  rx_input_memio_Mmux_lma_Result_10_1 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => rx_input_memio_macnt_80,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bpl(10),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(10)
    );
  rx_input_memio_Mmux_lma_Result_13_1 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bpl(13),
      ADR2 => rx_input_memio_macnt_83,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(13)
    );
  rx_input_memio_Mmux_lma_Result_12_1 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bpl(12),
      ADR2 => rx_input_memio_macnt_82,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(12)
    );
  rx_input_memio_addrchk_rxucastl_1636 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxucast,
      CE => rx_input_memio_addrchk_rxucastl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_rxucastl_FFY_RST,
      O => rx_input_memio_addrchk_rxucastl
    );
  rx_input_memio_addrchk_rxucastl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_rxucastl_FFY_RST
    );
  rx_input_memio_Mmux_lma_Result_15_1 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_macnt_85,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bpl(15),
      O => rx_input_memio_lma(15)
    );
  rx_input_memio_Mmux_lma_Result_14_1 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => rx_input_memio_bpl(14),
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_macnt_84,
      O => rx_input_memio_lma(14)
    );
  rx_input_memio_Mmux_lmd_Result_11_1 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_doutl(11),
      ADR2 => VCC,
      ADR3 => rx_input_memio_bcntl(11),
      O => rx_input_memio_lmd(11)
    );
  rx_input_memio_Mmux_lmd_Result_10_1 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(10),
      ADR1 => rx_input_memio_wbpl,
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(10),
      O => rx_input_memio_lmd(10)
    );
  rx_input_memio_Mmux_lmd_Result_21_1 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(21),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(21)
    );
  rx_input_memio_Mmux_lmd_Result_20_1 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_doutl(20),
      O => rx_input_memio_lmd(20)
    );
  rx_input_memio_Mmux_lmd_Result_13_1 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(13),
      ADR3 => rx_input_memio_bcntl(13),
      O => rx_input_memio_lmd(13)
    );
  rx_input_memio_Mmux_lmd_Result_12_1 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcntl(12),
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_doutl(12),
      O => rx_input_memio_lmd(12)
    );
  rx_input_memio_Mmux_lmd_Result_31_1 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(31),
      O => rx_input_memio_lmd(31)
    );
  rx_input_memio_Mmux_lmd_Result_30_1 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_doutl(30),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_lmd(30)
    );
  rx_input_memio_Mmux_lmd_Result_23_1 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(23),
      O => rx_input_memio_lmd(23)
    );
  rx_input_memio_Mmux_lmd_Result_22_1 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(22),
      ADR3 => VCC,
      O => rx_input_memio_lmd(22)
    );
  rx_input_memio_Mmux_lmd_Result_15_1 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(15),
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_doutl(15),
      O => rx_input_memio_lmd(15)
    );
  rx_input_memio_Mmux_lmd_Result_14_1 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_doutl(14),
      ADR2 => rx_input_memio_bcntl(14),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(14)
    );
  rx_input_memio_Mmux_lmd_Result_25_1 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_doutl(25),
      O => rx_input_memio_lmd(25)
    );
  rx_input_memio_Mmux_lmd_Result_24_1 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(24),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(24)
    );
  rx_input_memio_Mmux_lmd_Result_17_1 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => rx_input_memio_doutl(17),
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lmd(17)
    );
  rx_input_memio_Mmux_lmd_Result_16_1 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(16),
      ADR3 => VCC,
      O => rx_input_memio_lmd(16)
    );
  rx_input_memio_Mmux_lmd_Result_27_1 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_wbpl,
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(27),
      O => rx_input_memio_lmd(27)
    );
  rx_input_memio_Mmux_lmd_Result_26_1 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_doutl(26),
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lmd(26)
    );
  rx_input_memio_Mmux_lmd_Result_19_1 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => rx_input_memio_doutl(19),
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lmd(19)
    );
  rx_input_memio_Mmux_lmd_Result_18_1 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_doutl(18),
      ADR2 => VCC,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(18)
    );
  rx_input_memio_Mmux_lmd_Result_29_1 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => rx_input_memio_doutl(29),
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lmd(29)
    );
  rx_input_memio_Mmux_lmd_Result_28_1 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_doutl(28),
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lmd(28)
    );
  rx_output_Mmux_lma_Result_11_1 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => VCC,
      ADR2 => rx_output_mdl(11),
      ADR3 => rx_output_mdl(27),
      O => rx_output_lma(11)
    );
  rx_output_Mmux_lma_Result_10_1 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => rx_output_mdl(10),
      ADR1 => rx_output_lmasell,
      ADR2 => rx_output_mdl(26),
      ADR3 => VCC,
      O => rx_output_lma(10)
    );
  rx_output_fifodin_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_11_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_13_1 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => rx_output_mdl(13),
      ADR2 => rx_output_mdl(29),
      ADR3 => VCC,
      O => rx_output_lma(13)
    );
  rx_output_Mmux_lma_Result_12_1 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => rx_output_mdl(12),
      ADR2 => rx_output_mdl(28),
      ADR3 => VCC,
      O => rx_output_lma(12)
    );
  rx_output_fifodin_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_13_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_15_1 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => VCC,
      ADR2 => rx_output_mdl(31),
      ADR3 => rx_output_mdl(15),
      O => rx_output_lma(15)
    );
  rx_output_Mmux_lma_Result_14_1 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_mdl(30),
      ADR2 => rx_output_mdl(14),
      ADR3 => rx_output_lmasell,
      O => rx_output_lma(14)
    );
  rx_output_fifodin_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_15_CEMUXNOT
    );
  tx_input_enableintl_LOGIC_ONE_1637 : X_ONE
    port map (
      O => tx_input_enableintl_LOGIC_ONE
    );
  tx_input_srl16_enable_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_27,
      A1 => GLOBAL_LOGIC0_27,
      A2 => GLOBAL_LOGIC1_21,
      A3 => GLOBAL_LOGIC0_30,
      D => tx_input_enable,
      CE => tx_input_enableintl_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_enableintl_GSHIFT
    );
  tx_input_enableintl_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_enableintl_CEMUXNOT
    );
  tx_input_enableintl_YUSED : X_BUF
    port map (
      I => tx_input_enableintl_GSHIFT,
      O => tx_input_enableint
    );
  mac_control_PHY_status_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"BBAA"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd3,
      ADR1 => mac_control_PHY_status_done,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_cs_FFd2,
      O => mac_control_PHY_status_cs_FFd2_In
    );
  mac_control_PHY_status_cs_FFd1_In1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_done,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_cs_FFd2,
      O => mac_control_PHY_status_cs_FFd1_In
    );
  mac_control_PHY_status_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd5,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_done,
      ADR3 => VCC,
      O => mac_control_PHY_status_cs_FFd4_In
    );
  mac_control_PHY_status_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_phyaddrws,
      ADR3 => mac_control_PHY_status_cs_FFd4,
      O => mac_control_PHY_status_cs_FFd3_In
    );
  mac_control_PHY_status_cs_FFd6_In1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd7,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_done,
      ADR3 => VCC,
      O => mac_control_PHY_status_cs_FFd6_In
    );
  mac_control_PHY_status_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"FF0A"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd5,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_done,
      ADR3 => mac_control_PHY_status_cs_FFd6,
      O => mac_control_PHY_status_cs_FFd5_In
    );
  mac_control_PHY_status_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"AAEE"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd1,
      ADR1 => mac_control_PHY_status_cs_FFd4,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_phyaddrws,
      O => mac_control_PHY_status_cs_FFd8_In
    );
  mac_control_PHY_status_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"BABA"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd8,
      ADR1 => mac_control_PHY_status_done,
      ADR2 => mac_control_PHY_status_cs_FFd7,
      ADR3 => VCC,
      O => mac_control_PHY_status_cs_FFd7_In
    );
  slowclock_clkcnt_Madd_n0000_Mxor_Result_2_Result1 : X_LUT4
    generic map(
      INIT => X"5AAA"
    )
    port map (
      ADR0 => slowclock_clkcnt(2),
      ADR1 => VCC,
      ADR2 => slowclock_clkcnt(0),
      ADR3 => slowclock_clkcnt(1),
      O => slowclock_clkcnt_n0000(2)
    );
  tx_input_Mxor_lden_Result1 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_enableint,
      ADR2 => tx_input_enableintl,
      ADR3 => VCC,
      O => tx_input_lden
    );
  tx_input_den_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_den_CEMUXNOT
    );
  tx_input_Mmux_n0032_Result_1_1 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_n0074(1),
      ADR2 => tx_input_dinint(1),
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(1)
    );
  tx_input_Mmux_n0032_Result_0_1 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => tx_input_n0074(0),
      ADR1 => tx_input_dinint(0),
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(0)
    );
  tx_input_Mmux_n0032_Result_3_1 : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => tx_input_n0074(3),
      ADR1 => tx_input_dinint(3),
      ADR2 => tx_input_cs_FFd12,
      ADR3 => VCC,
      O => tx_input_n0032(3)
    );
  tx_input_Mmux_n0032_Result_2_1 : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => tx_input_dinint(2),
      ADR1 => tx_input_n0074(2),
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(2)
    );
  tx_input_Mmux_n0032_Result_5_1 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => tx_input_n0074(5),
      ADR1 => VCC,
      ADR2 => tx_input_dinint(5),
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(5)
    );
  tx_input_Mmux_n0032_Result_4_1 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_dinint(4),
      ADR2 => tx_input_cs_FFd12,
      ADR3 => tx_input_n0074(4),
      O => tx_input_n0032(4)
    );
  tx_input_Mmux_n0032_Result_7_1 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => tx_input_n0074(7),
      ADR1 => tx_input_dinint(7),
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(7)
    );
  tx_input_Mmux_n0032_Result_6_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => tx_input_dinint(6),
      ADR2 => VCC,
      ADR3 => tx_input_n0074(6),
      O => tx_input_n0032(6)
    );
  tx_input_Mmux_n0032_Result_9_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => tx_input_dinint(9),
      ADR2 => VCC,
      ADR3 => tx_input_n0074(9),
      O => tx_input_n0032(9)
    );
  tx_input_Mmux_n0032_Result_8_1 : X_LUT4
    generic map(
      INIT => X"B8B8"
    )
    port map (
      ADR0 => tx_input_dinint(8),
      ADR1 => tx_input_cs_FFd12,
      ADR2 => tx_input_n0074(8),
      ADR3 => VCC,
      O => tx_input_n0032(8)
    );
  rx_input_GMII_endf1 : X_LUT4
    generic map(
      INIT => X"FFBB"
    )
    port map (
      ADR0 => rx_input_GMII_rx_of,
      ADR1 => rx_input_GMII_rx_dvl,
      ADR2 => VCC,
      ADR3 => rx_input_GMII_rx_erl,
      O => rx_input_endfin_GROM
    );
  rx_input_endfin_YUSED : X_BUF
    port map (
      I => rx_input_endfin_GROM,
      O => rx_input_GMII_endf
    );
  rx_output_fifo_BU90 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N17,
      ADR2 => rx_output_fifo_N16,
      ADR3 => VCC,
      O => rx_output_fifo_N2259
    );
  rx_output_fifo_BU97 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N16,
      ADR3 => rx_output_fifo_N15,
      O => rx_output_fifo_N2299
    );
  tx_output_n0034_31_1 : X_LUT4
    generic map(
      INIT => X"F9F6"
    )
    port map (
      ADR0 => tx_output_data(2),
      ADR1 => tx_output_crcl(23),
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crcl(29),
      O => tx_output_n0034(31)
    );
  tx_output_n0034_2_1 : X_LUT4
    generic map(
      INIT => X"FF96"
    )
    port map (
      ADR0 => tx_output_crc_1_Q,
      ADR1 => tx_output_data(5),
      ADR2 => tx_output_crcl(26),
      ADR3 => tx_output_cs_FFd16,
      O => tx_output_n0034(2)
    );
  tx_output_cs_Out151 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd4,
      ADR1 => tx_output_cs_FFd5,
      ADR2 => tx_output_cs_FFd6,
      ADR3 => tx_output_cs_FFd8,
      O => tx_output_crcenl_FROM
    );
  tx_output_n00331 : X_LUT4
    generic map(
      INIT => X"0F0A"
    )
    port map (
      ADR0 => tx_output_cs_FFd12,
      ADR1 => VCC,
      ADR2 => RESET_IBUF,
      ADR3 => tx_output_decbcnt,
      O => tx_output_crcenl_GROM
    );
  tx_output_crcenl_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_crcenl_CEMUXNOT
    );
  tx_output_crcenl_XUSED : X_BUF
    port map (
      I => tx_output_crcenl_FROM,
      O => tx_output_decbcnt
    );
  tx_output_crcenl_YUSED : X_BUF
    port map (
      I => tx_output_crcenl_GROM,
      O => tx_output_n0033
    );
  mac_control_lsclkdelta1 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => mac_control_sclkl,
      ADR1 => mac_control_sclkll,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_lsclkdelta
    );
  mac_control_lmacaddr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_11_FFX_RST,
      O => mac_control_lmacaddr(11)
    );
  mac_control_lmacaddr_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_11_FFX_RST
    );
  rx_input_memio_crccomb_Mxor_CO_25_Xo_1_1_2_1638 : X_LUT4
    generic map(
      INIT => X"9696"
    )
    port map (
      ADR0 => rx_input_memio_crcl(26),
      ADR1 => rx_input_memio_crcl(17),
      ADR2 => rx_input_memio_datal(5),
      ADR3 => VCC,
      O => rx_input_memio_crcl_2_FROM
    );
  rx_input_memio_n0048_2_1 : X_LUT4
    generic map(
      INIT => X"F9F6"
    )
    port map (
      ADR0 => rx_input_memio_crc_1_Q,
      ADR1 => rx_input_memio_crcl(26),
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_datal(5),
      O => rx_input_memio_n0048(2)
    );
  rx_input_memio_crcl_2_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_2_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_25_Xo_1_1_2
    );
  mac_control_n00681 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_N52118,
      ADR1 => mac_control_din(6),
      ADR2 => mac_control_N52236,
      ADR3 => mac_control_newcmd,
      O => mac_control_n0068
    );
  mac_control_n00661 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_N52236,
      ADR1 => mac_control_N52118,
      ADR2 => mac_control_din(4),
      ADR3 => mac_control_newcmd,
      O => mac_control_n0066
    );
  rx_output_Mmux_lma_Result_1_1 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => rx_output_mdl(17),
      ADR1 => rx_output_lmasell,
      ADR2 => VCC,
      ADR3 => rx_output_mdl(1),
      O => rx_output_lma(1)
    );
  rx_output_Mmux_lma_Result_0_1 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => rx_output_mdl(0),
      ADR2 => rx_output_mdl(16),
      ADR3 => VCC,
      O => rx_output_lma(0)
    );
  rx_output_fifodin_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_1_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_3_1 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => VCC,
      ADR2 => rx_output_mdl(19),
      ADR3 => rx_output_mdl(3),
      O => rx_output_lma(3)
    );
  rx_output_Mmux_lma_Result_2_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => rx_output_mdl(18),
      ADR2 => VCC,
      ADR3 => rx_output_mdl(2),
      O => rx_output_lma(2)
    );
  rx_output_fifodin_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_3_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_5_1 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_mdl(21),
      ADR2 => rx_output_lmasell,
      ADR3 => rx_output_mdl(5),
      O => rx_output_lma(5)
    );
  rx_output_Mmux_lma_Result_4_1 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => rx_output_mdl(4),
      ADR1 => rx_output_lmasell,
      ADR2 => VCC,
      ADR3 => rx_output_mdl(20),
      O => rx_output_lma(4)
    );
  rx_output_fifodin_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_5_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_7_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => rx_output_mdl(23),
      ADR2 => VCC,
      ADR3 => rx_output_mdl(7),
      O => rx_output_lma(7)
    );
  rx_output_Mmux_lma_Result_6_1 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => rx_output_mdl(6),
      ADR2 => rx_output_mdl(22),
      ADR3 => VCC,
      O => rx_output_lma(6)
    );
  rx_output_fifodin_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_7_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_9_1 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => VCC,
      ADR2 => rx_output_mdl(9),
      ADR3 => rx_output_mdl(25),
      O => rx_output_lma(9)
    );
  rx_output_Mmux_lma_Result_8_1 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => VCC,
      ADR2 => rx_output_mdl(8),
      ADR3 => rx_output_mdl(24),
      O => rx_output_lma(8)
    );
  rx_output_fifodin_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_9_CEMUXNOT
    );
  rx_output_n00511 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => rx_output_fifo_wrcount(0),
      ADR1 => rx_output_fifo_wrcount(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0051
    );
  rx_output_fifo_full_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifo_full_CEMUXNOT
    );
  rx_input_GMII_lfifoin_0_11 : X_LUT4
    generic map(
      INIT => X"5000"
    )
    port map (
      ADR0 => rx_input_GMII_rx_of,
      ADR1 => VCC,
      ADR2 => rx_input_GMII_rx_dvl,
      ADR3 => rx_input_GMII_rxdl(0),
      O => rx_input_GMII_N80573
    );
  rx_input_GMII_lfifoin_1_11 : X_LUT4
    generic map(
      INIT => X"5000"
    )
    port map (
      ADR0 => rx_input_GMII_rx_erl,
      ADR1 => VCC,
      ADR2 => rx_input_GMII_rxdl(1),
      ADR3 => rx_input_GMII_rx_dvl,
      O => rx_input_GMII_N80576
    );
  rx_input_GMII_lfifoin_3_11 : X_LUT4
    generic map(
      INIT => X"2200"
    )
    port map (
      ADR0 => rx_input_GMII_rx_dvl,
      ADR1 => rx_input_GMII_rx_erl,
      ADR2 => VCC,
      ADR3 => rx_input_GMII_rxdl(3),
      O => rx_input_GMII_N80582
    );
  rx_input_GMII_lfifoin_2_11 : X_LUT4
    generic map(
      INIT => X"EECC"
    )
    port map (
      ADR0 => rx_input_GMII_rx_dvl,
      ADR1 => rx_input_GMII_rx_erl,
      ADR2 => VCC,
      ADR3 => rx_input_GMII_rxdl(2),
      O => rx_input_GMII_N80579
    );
  mac_control_lmacaddr_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_21_FFX_RST,
      O => mac_control_lmacaddr(21)
    );
  mac_control_lmacaddr_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_21_FFX_RST
    );
  rx_input_GMII_lfifoin_5_11 : X_LUT4
    generic map(
      INIT => X"0808"
    )
    port map (
      ADR0 => rx_input_GMII_rx_dvl,
      ADR1 => rx_input_GMII_rxdl(5),
      ADR2 => rx_input_GMII_rx_erl,
      ADR3 => VCC,
      O => rx_input_GMII_N80561
    );
  rx_input_GMII_lfifoin_4_11 : X_LUT4
    generic map(
      INIT => X"0C00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_GMII_rxdl(4),
      ADR2 => rx_input_GMII_rx_erl,
      ADR3 => rx_input_GMII_rx_dvl,
      O => rx_input_GMII_N80570
    );
  rx_input_GMII_lfifoin_7_11 : X_LUT4
    generic map(
      INIT => X"2200"
    )
    port map (
      ADR0 => rx_input_GMII_rxdl(7),
      ADR1 => rx_input_GMII_rx_erl,
      ADR2 => VCC,
      ADR3 => rx_input_GMII_rx_dvl,
      O => rx_input_GMII_N80567
    );
  rx_input_GMII_lfifoin_6_11 : X_LUT4
    generic map(
      INIT => X"00A0"
    )
    port map (
      ADR0 => rx_input_GMII_rx_dvl,
      ADR1 => VCC,
      ADR2 => rx_input_GMII_rxdl(6),
      ADR3 => rx_input_GMII_rx_erl,
      O => rx_input_GMII_N80564
    );
  tx_input_dinint_11_LOGIC_ONE_1639 : X_ONE
    port map (
      O => tx_input_dinint_11_LOGIC_ONE
    );
  tx_input_srl16_din_bit11_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_29,
      A1 => GLOBAL_LOGIC0_29,
      A2 => GLOBAL_LOGIC1_22,
      A3 => GLOBAL_LOGIC0_24,
      D => tx_input_dinl(11),
      CE => tx_input_dinint_11_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(11)
    );
  tx_input_srl16_din_bit10_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_29,
      A1 => GLOBAL_LOGIC0_29,
      A2 => GLOBAL_LOGIC1_22,
      A3 => GLOBAL_LOGIC0_24,
      D => tx_input_dinl(10),
      CE => tx_input_dinint_11_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(10)
    );
  tx_input_dinint_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_11_CEMUXNOT
    );
  tx_input_dinint_13_LOGIC_ONE_1640 : X_ONE
    port map (
      O => tx_input_dinint_13_LOGIC_ONE
    );
  tx_input_srl16_din_bit13_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_20,
      A1 => GLOBAL_LOGIC0_20,
      A2 => GLOBAL_LOGIC1_25,
      A3 => GLOBAL_LOGIC0_25,
      D => tx_input_dinl(13),
      CE => tx_input_dinint_13_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(13)
    );
  tx_input_srl16_din_bit12_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_20,
      A1 => GLOBAL_LOGIC0_20,
      A2 => GLOBAL_LOGIC1_25,
      A3 => GLOBAL_LOGIC0_25,
      D => tx_input_dinl(12),
      CE => tx_input_dinint_13_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(12)
    );
  tx_input_dinint_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_13_CEMUXNOT
    );
  tx_input_dinint_15_LOGIC_ONE_1641 : X_ONE
    port map (
      O => tx_input_dinint_15_LOGIC_ONE
    );
  tx_input_srl16_din_bit15_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_18,
      A1 => GLOBAL_LOGIC0_18,
      A2 => GLOBAL_LOGIC1_30,
      A3 => GLOBAL_LOGIC0_18,
      D => tx_input_dinl(15),
      CE => tx_input_dinint_15_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(15)
    );
  tx_input_srl16_din_bit14_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_18,
      A1 => GLOBAL_LOGIC0_19,
      A2 => GLOBAL_LOGIC1_30,
      A3 => GLOBAL_LOGIC0_18,
      D => tx_input_dinl(14),
      CE => tx_input_dinint_15_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(14)
    );
  tx_input_dinint_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_15_CEMUXNOT
    );
  rx_input_memio_n00611 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => rx_input_memio_crcequal,
      ADR1 => rx_input_memio_endbyte(2),
      ADR2 => rx_input_memio_cs_FFd5,
      ADR3 => rxfifofull,
      O => rx_input_memio_n0061
    );
  rx_input_memio_n00601 : X_LUT4
    generic map(
      INIT => X"0202"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd5,
      ADR1 => rx_input_memio_crcequal,
      ADR2 => rx_input_memio_endbyte(2),
      ADR3 => VCC,
      O => rx_input_memio_n0060
    );
  rxfifowerr_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxfifowerr_CEMUXNOT
    );
  rx_output_cs_FFd17_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd17_FFY_RST
    );
  rx_output_cs_FFd17_1642 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd17_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd17_FFY_RST,
      O => rx_output_cs_FFd17
    );
  rx_output_cs_FFd17_In1 : X_LUT4
    generic map(
      INIT => X"0200"
    )
    port map (
      ADR0 => rx_output_cs_FFd18,
      ADR1 => rx_output_n0017,
      ADR2 => memcontroller_clknum(0),
      ADR3 => memcontroller_clknum(1),
      O => rx_output_cs_FFd17_In
    );
  rx_output_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"0808"
    )
    port map (
      ADR0 => rx_output_nf,
      ADR1 => rx_output_cs_FFd7,
      ADR2 => rx_output_fifo_full,
      ADR3 => VCC,
      O => rx_output_cs_FFd5_In
    );
  rx_output_cs_FFd19_In1 : X_LUT4
    generic map(
      INIT => X"FCDC"
    )
    port map (
      ADR0 => rx_output_nf,
      ADR1 => rx_output_cs_FFd10,
      ADR2 => rx_output_cs_FFd19,
      ADR3 => rx_output_nfl,
      O => rx_output_cs_FFd19_In
    );
  rx_input_memio_n00581 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => rx_input_memio_endbyte(0),
      ADR1 => rx_input_memio_cs_FFd5,
      ADR2 => rx_input_memio_endbyte(1),
      ADR3 => rx_input_memio_endbyte(2),
      O => rx_input_memio_n0058
    );
  rx_input_memio_n00571 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => rx_input_memio_endbyte(1),
      ADR1 => rx_input_memio_endbyte(0),
      ADR2 => rx_input_memio_cs_FFd5,
      ADR3 => rx_input_memio_endbyte(2),
      O => rx_input_memio_n0057
    );
  rxoferr_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rxoferr_CEMUXNOT
    );
  tx_input_cs_FFd10_In_SW0 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_den,
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd10,
      O => tx_input_cs_FFd11_FROM
    );
  tx_input_cs_FFd11_In1 : X_LUT4
    generic map(
      INIT => X"8800"
    )
    port map (
      ADR0 => tx_input_newfint,
      ADR1 => tx_input_den,
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_cs_FFd11_In
    );
  tx_input_cs_FFd11_XUSED : X_BUF
    port map (
      I => tx_input_cs_FFd11_FROM,
      O => tx_input_N69350
    );
  tx_input_Mmux_n0032_Result_11_1 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => tx_input_n0074(11),
      ADR1 => tx_input_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_input_dinint(11),
      O => tx_input_n0032(11)
    );
  tx_input_Mmux_n0032_Result_10_1 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => tx_input_dinint(10),
      ADR1 => tx_input_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_input_n0074(10),
      O => tx_input_n0032(10)
    );
  mac_control_lmacaddr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_13_FFX_RST,
      O => mac_control_lmacaddr(13)
    );
  mac_control_lmacaddr_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_13_FFX_RST
    );
  tx_input_Mmux_n0032_Result_13_1 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => tx_input_n0074(13),
      ADR1 => VCC,
      ADR2 => tx_input_cs_FFd12,
      ADR3 => tx_input_dinint(13),
      O => tx_input_n0032(13)
    );
  tx_input_Mmux_n0032_Result_12_1 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => VCC,
      ADR2 => tx_input_n0074(12),
      ADR3 => tx_input_dinint(12),
      O => tx_input_n0032(12)
    );
  tx_input_Mmux_n0032_Result_15_1 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => tx_input_dinint(15),
      ADR1 => tx_input_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_input_n0074(15),
      O => tx_input_n0032(15)
    );
  tx_input_Mmux_n0032_Result_14_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => tx_input_dinint(14),
      ADR2 => VCC,
      ADR3 => tx_input_n0074(14),
      O => tx_input_n0032(14)
    );
  tx_input_dinint_1_LOGIC_ONE_1643 : X_ONE
    port map (
      O => tx_input_dinint_1_LOGIC_ONE
    );
  tx_input_srl16_din_bit1_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_33,
      A1 => GLOBAL_LOGIC0_2,
      A2 => GLOBAL_LOGIC1_36,
      A3 => GLOBAL_LOGIC0_2,
      D => tx_input_dinl(1),
      CE => tx_input_dinint_1_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(1)
    );
  tx_input_srl16_din_bit0_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_33,
      A1 => GLOBAL_LOGIC0_2,
      A2 => GLOBAL_LOGIC1_36,
      A3 => GLOBAL_LOGIC0_2,
      D => tx_input_dinl(0),
      CE => tx_input_dinint_1_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(0)
    );
  tx_input_dinint_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_1_CEMUXNOT
    );
  tx_input_dinint_3_LOGIC_ONE_1644 : X_ONE
    port map (
      O => tx_input_dinint_3_LOGIC_ONE
    );
  tx_input_srl16_din_bit3_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_28,
      A1 => GLOBAL_LOGIC0_28,
      A2 => GLOBAL_LOGIC1_23,
      A3 => GLOBAL_LOGIC0_26,
      D => tx_input_dinl(3),
      CE => tx_input_dinint_3_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(3)
    );
  tx_input_srl16_din_bit2_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_28,
      A1 => GLOBAL_LOGIC0_28,
      A2 => GLOBAL_LOGIC1_23,
      A3 => GLOBAL_LOGIC0_26,
      D => tx_input_dinl(2),
      CE => tx_input_dinint_3_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(2)
    );
  tx_input_dinint_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_3_CEMUXNOT
    );
  tx_input_dinint_5_LOGIC_ONE_1645 : X_ONE
    port map (
      O => tx_input_dinint_5_LOGIC_ONE
    );
  tx_input_srl16_din_bit5_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_26,
      A1 => GLOBAL_LOGIC0_28,
      A2 => GLOBAL_LOGIC1_23,
      A3 => GLOBAL_LOGIC0_28,
      D => tx_input_dinl(5),
      CE => tx_input_dinint_5_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(5)
    );
  tx_input_srl16_din_bit4_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_26,
      A1 => GLOBAL_LOGIC0_28,
      A2 => GLOBAL_LOGIC1_23,
      A3 => GLOBAL_LOGIC0_28,
      D => tx_input_dinl(4),
      CE => tx_input_dinint_5_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(4)
    );
  tx_input_dinint_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_5_CEMUXNOT
    );
  tx_input_dinint_7_LOGIC_ONE_1646 : X_ONE
    port map (
      O => tx_input_dinint_7_LOGIC_ONE
    );
  tx_input_srl16_din_bit7_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_23,
      A1 => GLOBAL_LOGIC0_23,
      A2 => GLOBAL_LOGIC1_26,
      A3 => GLOBAL_LOGIC0_22,
      D => tx_input_dinl(7),
      CE => tx_input_dinint_7_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(7)
    );
  tx_input_srl16_din_bit6_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_23,
      A1 => GLOBAL_LOGIC0_23,
      A2 => GLOBAL_LOGIC1_26,
      A3 => GLOBAL_LOGIC0_20,
      D => tx_input_dinl(6),
      CE => tx_input_dinint_7_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(6)
    );
  tx_input_dinint_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_7_CEMUXNOT
    );
  tx_input_dinint_9_LOGIC_ONE_1647 : X_ONE
    port map (
      O => tx_input_dinint_9_LOGIC_ONE
    );
  tx_input_srl16_din_bit9_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_24,
      A1 => GLOBAL_LOGIC0_24,
      A2 => GLOBAL_LOGIC1_29,
      A3 => GLOBAL_LOGIC0_20,
      D => tx_input_dinl(9),
      CE => tx_input_dinint_9_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(9)
    );
  tx_input_srl16_din_bit8_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_24,
      A1 => GLOBAL_LOGIC0_24,
      A2 => GLOBAL_LOGIC1_29,
      A3 => GLOBAL_LOGIC0_20,
      D => tx_input_dinl(8),
      CE => tx_input_dinint_9_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(8)
    );
  tx_input_dinint_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_9_CEMUXNOT
    );
  mac_control_Mshreg_scslll_srl_17 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_24,
      A1 => GLOBAL_LOGIC0_8,
      A2 => GLOBAL_LOGIC0_8,
      A3 => GLOBAL_LOGIC0_8,
      D => SCS_IBUF,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      Q => mac_control_Mshreg_scslll_net187
    );
  rx_input_memio_Mshreg_lbpout4_5_srl_10 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_49,
      A1 => GLOBAL_LOGIC1_9,
      A2 => GLOBAL_LOGIC0_49,
      A3 => GLOBAL_LOGIC0_45,
      D => rx_input_memio_bp(5),
      CE => rx_input_memio_Mshreg_lbpout4_5_64_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_5_net24
    );
  rx_input_memio_Mshreg_lbpout4_5_64_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_5_64_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_5_64_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_5_64_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_6_srl_9 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_44,
      A1 => GLOBAL_LOGIC1_12,
      A2 => GLOBAL_LOGIC0_44,
      A3 => GLOBAL_LOGIC0_42,
      D => rx_input_memio_bp(6),
      CE => rx_input_memio_Mshreg_lbpout4_6_63_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_6_net22
    );
  rx_input_memio_Mshreg_lbpout4_6_63_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_6_63_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_6_63_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_6_63_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_7_srl_8 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_48,
      A1 => GLOBAL_LOGIC1_10,
      A2 => GLOBAL_LOGIC0_44,
      A3 => GLOBAL_LOGIC0_44,
      D => rx_input_memio_bp(7),
      CE => rx_input_memio_Mshreg_lbpout4_7_62_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_7_net20
    );
  rx_input_memio_Mshreg_lbpout4_7_62_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_7_62_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_7_62_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_7_62_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_8_srl_7 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_36,
      A1 => GLOBAL_LOGIC1_16,
      A2 => GLOBAL_LOGIC0_36,
      A3 => GLOBAL_LOGIC0_37,
      D => rx_input_memio_bp(8),
      CE => rx_input_memio_Mshreg_lbpout4_8_61_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_8_net18
    );
  rx_input_memio_Mshreg_lbpout4_8_61_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_8_61_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_8_61_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_8_61_SRMUX_OUTPUTNOT
    );
  mac_control_lmacaddr_33 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_33_FFX_RST,
      O => mac_control_lmacaddr(33)
    );
  mac_control_lmacaddr_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_33_FFX_RST
    );
  rx_input_memio_Mshreg_lbpout4_9_srl_6 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_38,
      A1 => GLOBAL_LOGIC1_13,
      A2 => GLOBAL_LOGIC0_41,
      A3 => GLOBAL_LOGIC0_41,
      D => rx_input_memio_bp(9),
      CE => rx_input_memio_Mshreg_lbpout4_9_60_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_9_net16
    );
  rx_input_memio_Mshreg_lbpout4_9_60_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_9_60_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_9_60_SRMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_9_60_SRMUX_OUTPUTNOT
    );
  tx_input_newfint_LOGIC_ONE_1648 : X_ONE
    port map (
      O => tx_input_newfint_LOGIC_ONE
    );
  tx_input_srl16_newframe_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_31,
      A1 => GLOBAL_LOGIC0_27,
      A2 => GLOBAL_LOGIC1_18,
      A3 => GLOBAL_LOGIC0_31,
      D => tx_input_newframel,
      CE => tx_input_newfint_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_lnewfint
    );
  tx_input_newfint_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_newfint_CEMUXNOT
    );
  tx_output_n0034_21_1 : X_LUT4
    generic map(
      INIT => X"EBBE"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => tx_output_data(2),
      ADR2 => tx_output_crcl(29),
      ADR3 => tx_output_crcl(13),
      O => tx_output_n0034(21)
    );
  tx_output_n0034_20_1 : X_LUT4
    generic map(
      INIT => X"F9F6"
    )
    port map (
      ADR0 => tx_output_data(3),
      ADR1 => tx_output_crcl(12),
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crcl(28),
      O => tx_output_n0034(20)
    );
  tx_output_crc_loigc_Mxor_CO_26_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(28),
      ADR1 => tx_output_data(3),
      ADR2 => tx_output_crcl(24),
      ADR3 => tx_output_data(7),
      O => tx_output_crcl_22_FROM
    );
  tx_output_n0034_22_1 : X_LUT4
    generic map(
      INIT => X"EDDE"
    )
    port map (
      ADR0 => tx_output_crcl(24),
      ADR1 => tx_output_cs_FFd16,
      ADR2 => tx_output_crcl(14),
      ADR3 => tx_output_data(7),
      O => tx_output_n0034(22)
    );
  tx_output_crcl_22_XUSED : X_BUF
    port map (
      I => tx_output_crcl_22_FROM,
      O => tx_output_crc_loigc_Mxor_CO_26_Xo(1)
    );
  mac_control_Mmux_n0017_Result_0_9 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_N52118,
      ADR1 => mac_control_rxoferr_cnt(0),
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_rxf_cnt(0),
      O => mac_control_CHOICE2197_FROM
    );
  mac_control_Mmux_n0017_Result_10_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(10),
      ADR1 => mac_control_rxoferr_cnt(10),
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_N52111,
      O => mac_control_CHOICE2197_GROM
    );
  mac_control_CHOICE2197_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2197_FROM,
      O => mac_control_CHOICE2197
    );
  mac_control_CHOICE2197_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2197_GROM,
      O => mac_control_CHOICE2423
    );
  mac_control_Mmux_n0017_Result_2_31 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_txf_cnt(2),
      ADR1 => mac_control_phydi(2),
      ADR2 => mac_control_N52132,
      ADR3 => mac_control_N52118,
      O => mac_control_CHOICE2277_FROM
    );
  mac_control_Mmux_n0017_Result_10_31 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_txf_cnt(10),
      ADR1 => mac_control_phydi(10),
      ADR2 => mac_control_N52132,
      ADR3 => mac_control_N52118,
      O => mac_control_CHOICE2277_GROM
    );
  mac_control_CHOICE2277_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2277_FROM,
      O => mac_control_CHOICE2277
    );
  mac_control_CHOICE2277_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2277_GROM,
      O => mac_control_CHOICE2429
    );
  mac_control_Mmux_n0017_Result_26_34 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0078,
      ADR1 => mac_control_n0079,
      ADR2 => mac_control_txf_cnt(26),
      ADR3 => mac_control_rxf_cnt(26),
      O => mac_control_CHOICE2021_FROM
    );
  mac_control_Mmux_n0017_Result_11_20 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0078,
      ADR1 => mac_control_rxf_cnt(11),
      ADR2 => mac_control_n0079,
      ADR3 => mac_control_txf_cnt(11),
      O => mac_control_CHOICE2021_GROM
    );
  mac_control_CHOICE2021_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2021_FROM,
      O => mac_control_CHOICE2021
    );
  mac_control_CHOICE2021_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2021_GROM,
      O => mac_control_CHOICE2857
    );
  mac_control_Mmux_n0017_Result_11_30 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_n0073,
      ADR1 => mac_control_phystat(11),
      ADR2 => mac_control_n0074,
      ADR3 => mac_control_N81785,
      O => mac_control_dout_11_FROM
    );
  mac_control_Mmux_n0017_Result_11_108 : X_LUT4
    generic map(
      INIT => X"FAEA"
    )
    port map (
      ADR0 => mac_control_N82013,
      ADR1 => mac_control_CHOICE2874,
      ADR2 => mac_control_N52163,
      ADR3 => mac_control_CHOICE2859,
      O => mac_control_N79864
    );
  mac_control_dout_11_XUSED : X_BUF
    port map (
      I => mac_control_dout_11_FROM,
      O => mac_control_CHOICE2859
    );
  mac_control_Mmux_n0017_Result_10_39 : X_LUT4
    generic map(
      INIT => X"A888"
    )
    port map (
      ADR0 => mac_control_N52220,
      ADR1 => mac_control_CHOICE2429,
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_rxphyerr_cnt(10),
      O => mac_control_CHOICE2431_FROM
    );
  mac_control_Mmux_n0017_Result_10_45 : X_LUT4
    generic map(
      INIT => X"FFA8"
    )
    port map (
      ADR0 => mac_control_N52228,
      ADR1 => mac_control_CHOICE2420,
      ADR2 => mac_control_CHOICE2423,
      ADR3 => mac_control_CHOICE2431,
      O => mac_control_CHOICE2431_GROM
    );
  mac_control_CHOICE2431_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2431_FROM,
      O => mac_control_CHOICE2431
    );
  mac_control_CHOICE2431_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2431_GROM,
      O => mac_control_CHOICE2432
    );
  mac_control_Mmux_n0017_Result_7_15 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0077,
      ADR1 => mac_control_phydi(7),
      ADR2 => mac_control_n0076,
      ADR3 => mac_control_phydo(7),
      O => mac_control_CHOICE2822_FROM
    );
  mac_control_Mmux_n0017_Result_11_15 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0077,
      ADR1 => mac_control_phydo(11),
      ADR2 => mac_control_n0076,
      ADR3 => mac_control_phydi(11),
      O => mac_control_CHOICE2822_GROM
    );
  mac_control_CHOICE2822_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2822_FROM,
      O => mac_control_CHOICE2822
    );
  mac_control_CHOICE2822_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2822_GROM,
      O => mac_control_CHOICE2854
    );
  mac_control_Mmux_n0017_Result_12_12 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_phydi(12),
      ADR1 => mac_control_n0073,
      ADR2 => mac_control_n0076,
      ADR3 => mac_control_phystat(12),
      O => mac_control_CHOICE2665_FROM
    );
  mac_control_Mmux_n0017_Result_12_94_1_1649 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE2662,
      ADR3 => mac_control_CHOICE2665,
      O => mac_control_CHOICE2665_GROM
    );
  mac_control_CHOICE2665_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2665_FROM,
      O => mac_control_CHOICE2665
    );
  mac_control_CHOICE2665_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2665_GROM,
      O => mac_control_Mmux_n0017_Result_12_94_1
    );
  mac_control_lmacaddr_41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_41_FFX_RST,
      O => mac_control_lmacaddr(41)
    );
  mac_control_lmacaddr_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_41_FFX_RST
    );
  mac_control_Mmux_n0017_Result_11_60 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_lmacaddr(11),
      ADR1 => mac_control_n0085,
      ADR2 => mac_control_rxcrcerr_cnt(11),
      ADR3 => mac_control_n0084,
      O => mac_control_CHOICE2869_FROM
    );
  mac_control_Mmux_n0017_Result_11_74_SW0 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(11),
      ADR1 => mac_control_CHOICE2872,
      ADR2 => mac_control_n0081,
      ADR3 => mac_control_CHOICE2869,
      O => mac_control_CHOICE2869_GROM
    );
  mac_control_CHOICE2869_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2869_FROM,
      O => mac_control_CHOICE2869
    );
  mac_control_CHOICE2869_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2869_GROM,
      O => mac_control_N81769
    );
  mac_control_Mmux_n0017_Result_20_12 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0082,
      ADR1 => mac_control_rxoferr_cnt(20),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_rxphyerr_cnt(20),
      O => mac_control_CHOICE1942_FROM
    );
  mac_control_Mmux_n0017_Result_20_66_1_1650 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_CHOICE1939,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE1942,
      O => mac_control_CHOICE1942_GROM
    );
  mac_control_CHOICE1942_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1942_FROM,
      O => mac_control_CHOICE1942
    );
  mac_control_CHOICE1942_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1942_GROM,
      O => mac_control_Mmux_n0017_Result_20_66_1
    );
  mac_control_Mmux_n0017_Result_6_69 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cnt(6),
      ADR1 => mac_control_txfifowerr_cnt(6),
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_N52118,
      O => mac_control_CHOICE2322_FROM
    );
  mac_control_Mmux_n0017_Result_10_69 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_N52111,
      ADR1 => mac_control_N52118,
      ADR2 => mac_control_txfifowerr_cnt(10),
      ADR3 => mac_control_rxcrcerr_cnt(10),
      O => mac_control_CHOICE2322_GROM
    );
  mac_control_CHOICE2322_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2322_FROM,
      O => mac_control_CHOICE2322
    );
  mac_control_CHOICE2322_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2322_GROM,
      O => mac_control_CHOICE2436
    );
  mac_control_Mmux_n0017_Result_5_86 : X_LUT4
    generic map(
      INIT => X"8A80"
    )
    port map (
      ADR0 => mac_control_N52143,
      ADR1 => mac_control_lmacaddr(37),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_lmacaddr(21),
      O => mac_control_CHOICE2366_FROM
    );
  mac_control_Mmux_n0017_Result_10_86 : X_LUT4
    generic map(
      INIT => X"E040"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => mac_control_lmacaddr(26),
      ADR2 => mac_control_N52143,
      ADR3 => mac_control_lmacaddr(42),
      O => mac_control_CHOICE2366_GROM
    );
  mac_control_CHOICE2366_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2366_FROM,
      O => mac_control_CHOICE2366
    );
  mac_control_CHOICE2366_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2366_GROM,
      O => mac_control_CHOICE2442
    );
  mac_control_Mmux_n0017_Result_12_40 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(12),
      ADR1 => mac_control_txfifowerr_cnt(12),
      ADR2 => mac_control_n0080,
      ADR3 => mac_control_n0079,
      O => mac_control_CHOICE2673_FROM
    );
  mac_control_Mmux_n0017_Result_12_94_SW0_2_1651 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => mac_control_CHOICE2676,
      ADR1 => mac_control_CHOICE2668,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2673,
      O => mac_control_CHOICE2673_GROM
    );
  mac_control_CHOICE2673_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2673_FROM,
      O => mac_control_CHOICE2673
    );
  mac_control_CHOICE2673_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2673_GROM,
      O => mac_control_Mmux_n0017_Result_12_94_SW0_2
    );
  mac_control_Mmux_n0017_Result_7_48 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxoferr_cnt(7),
      ADR1 => mac_control_rxphyerr_cnt(7),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_n0082,
      O => mac_control_CHOICE2833_FROM
    );
  mac_control_Mmux_n0017_Result_11_48 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(11),
      ADR1 => mac_control_rxoferr_cnt(11),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_n0082,
      O => mac_control_CHOICE2833_GROM
    );
  mac_control_CHOICE2833_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2833_FROM,
      O => mac_control_CHOICE2833
    );
  mac_control_CHOICE2833_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2833_GROM,
      O => mac_control_CHOICE2865
    );
  mac_control_Mmux_n0017_Result_4_17 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cnt(4),
      ADR1 => mac_control_n0078,
      ADR2 => mac_control_phydo(4),
      ADR3 => mac_control_n0077,
      O => mac_control_CHOICE2606_FROM
    );
  mac_control_Mmux_n0017_Result_12_17 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phydo(12),
      ADR1 => mac_control_n0078,
      ADR2 => mac_control_txf_cnt(12),
      ADR3 => mac_control_n0077,
      O => mac_control_CHOICE2606_GROM
    );
  mac_control_CHOICE2606_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2606_FROM,
      O => mac_control_CHOICE2606
    );
  mac_control_CHOICE2606_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2606_GROM,
      O => mac_control_CHOICE2668
    );
  mac_control_Mmux_n0017_Result_2_86 : X_LUT4
    generic map(
      INIT => X"CA00"
    )
    port map (
      ADR0 => mac_control_lmacaddr(18),
      ADR1 => mac_control_lmacaddr(34),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_N52143,
      O => mac_control_CHOICE2290_FROM
    );
  mac_control_Mmux_n0017_Result_11_65 : X_LUT4
    generic map(
      INIT => X"A0C0"
    )
    port map (
      ADR0 => mac_control_lmacaddr(43),
      ADR1 => mac_control_lmacaddr(27),
      ADR2 => mac_control_N52143,
      ADR3 => mac_control_addr(0),
      O => mac_control_CHOICE2290_GROM
    );
  mac_control_CHOICE2290_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2290_FROM,
      O => mac_control_CHOICE2290
    );
  mac_control_CHOICE2290_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2290_GROM,
      O => mac_control_CHOICE2872
    );
  mac_control_Mmux_n0017_Result_20_7 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(20),
      ADR1 => mac_control_rxfifowerr_cnt(20),
      ADR2 => mac_control_n0081,
      ADR3 => mac_control_n0080,
      O => mac_control_CHOICE1939_FROM
    );
  mac_control_Mmux_n0017_Result_11_74 : X_LUT4
    generic map(
      INIT => X"FEEE"
    )
    port map (
      ADR0 => mac_control_CHOICE2865,
      ADR1 => mac_control_N81769,
      ADR2 => mac_control_n0080,
      ADR3 => mac_control_txfifowerr_cnt(11),
      O => mac_control_CHOICE1939_GROM
    );
  mac_control_CHOICE1939_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1939_FROM,
      O => mac_control_CHOICE1939
    );
  mac_control_CHOICE1939_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1939_GROM,
      O => mac_control_CHOICE2874
    );
  mac_control_lmacaddr_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_17_FFX_RST,
      O => mac_control_lmacaddr(17)
    );
  mac_control_lmacaddr_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_17_FFX_RST
    );
  mac_control_Mmux_n0017_Result_20_42 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_20_42_1,
      ADR1 => mac_control_CHOICE1952,
      ADR2 => mac_control_CHOICE1949,
      ADR3 => mac_control_Mmux_n0017_Result_20_42_SW0_1,
      O => mac_control_dout_20_FROM
    );
  mac_control_Mmux_n0017_Result_20_77 : X_LUT4
    generic map(
      INIT => X"BBB3"
    )
    port map (
      ADR0 => mac_control_N52163,
      ADR1 => mac_control_Mmux_n0017_Result_20_77_1,
      ADR2 => mac_control_Mmux_n0017_Result_20_66_1,
      ADR3 => mac_control_CHOICE1954,
      O => mac_control_N74952
    );
  mac_control_dout_20_XUSED : X_BUF
    port map (
      I => mac_control_dout_20_FROM,
      O => mac_control_CHOICE1954
    );
  mac_control_Mmux_n0017_Result_7_20 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(7),
      ADR1 => mac_control_n0079,
      ADR2 => mac_control_n0078,
      ADR3 => mac_control_txf_cnt(7),
      O => mac_control_CHOICE2825_FROM
    );
  mac_control_Mmux_n0017_Result_20_34 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0078,
      ADR1 => mac_control_n0079,
      ADR2 => mac_control_rxf_cnt(20),
      ADR3 => mac_control_txf_cnt(20),
      O => mac_control_CHOICE2825_GROM
    );
  mac_control_CHOICE2825_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2825_FROM,
      O => mac_control_CHOICE2825
    );
  mac_control_CHOICE2825_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2825_GROM,
      O => mac_control_CHOICE1952
    );
  mac_control_Mmux_n0017_Result_21_12 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0083,
      ADR1 => mac_control_rxcrcerr_cnt(21),
      ADR2 => mac_control_n0084,
      ADR3 => mac_control_rxoferr_cnt(21),
      O => mac_control_CHOICE2151_FROM
    );
  mac_control_Mmux_n0017_Result_21_69_1_1652 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => mac_control_CHOICE2148,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2151,
      O => mac_control_CHOICE2151_GROM
    );
  mac_control_CHOICE2151_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2151_FROM,
      O => mac_control_CHOICE2151
    );
  mac_control_CHOICE2151_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2151_GROM,
      O => mac_control_Mmux_n0017_Result_21_69_1
    );
  mac_control_Mmux_n0017_Result_13_12 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phystat(13),
      ADR1 => mac_control_phydi(13),
      ADR2 => mac_control_n0076,
      ADR3 => mac_control_n0073,
      O => mac_control_CHOICE2696_FROM
    );
  mac_control_Mmux_n0017_Result_13_94_1_1653 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => mac_control_CHOICE2693,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2696,
      O => mac_control_CHOICE2696_GROM
    );
  mac_control_CHOICE2696_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2696_FROM,
      O => mac_control_CHOICE2696
    );
  mac_control_CHOICE2696_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2696_GROM,
      O => mac_control_Mmux_n0017_Result_13_94_1
    );
  mac_control_Mmux_n0017_Result_17_7 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0081,
      ADR1 => mac_control_rxphyerr_cnt(17),
      ADR2 => mac_control_rxfifowerr_cnt(17),
      ADR3 => mac_control_n0082,
      O => mac_control_CHOICE2124_FROM
    );
  mac_control_Mmux_n0017_Result_12_45 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(12),
      ADR1 => mac_control_rxphyerr_cnt(12),
      ADR2 => mac_control_n0081,
      ADR3 => mac_control_n0082,
      O => mac_control_CHOICE2124_GROM
    );
  mac_control_CHOICE2124_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2124_FROM,
      O => mac_control_CHOICE2124
    );
  mac_control_CHOICE2124_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2124_GROM,
      O => mac_control_CHOICE2676
    );
  mac_control_Mmux_n0017_Result_26_29 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phystat(26),
      ADR1 => mac_control_n0073,
      ADR2 => mac_control_n0076,
      ADR3 => mac_control_phydi(26),
      O => mac_control_CHOICE2018_FROM
    );
  mac_control_Mmux_n0017_Result_20_29 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0073,
      ADR1 => mac_control_n0076,
      ADR2 => mac_control_phydi(20),
      ADR3 => mac_control_phystat(20),
      O => mac_control_CHOICE2018_GROM
    );
  mac_control_CHOICE2018_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2018_FROM,
      O => mac_control_CHOICE2018
    );
  mac_control_CHOICE2018_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2018_GROM,
      O => mac_control_CHOICE1949
    );
  mac_control_Mmux_n0017_Result_12_62 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_lmacaddr(28),
      ADR1 => mac_control_n0085,
      ADR2 => mac_control_n0086,
      ADR3 => mac_control_lmacaddr(12),
      O => mac_control_CHOICE2683_FROM
    );
  mac_control_Mmux_n0017_Result_12_63 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => mac_control_CHOICE2680,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2683,
      O => mac_control_CHOICE2683_GROM
    );
  mac_control_CHOICE2683_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2683_FROM,
      O => mac_control_CHOICE2683
    );
  mac_control_CHOICE2683_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2683_GROM,
      O => mac_control_CHOICE2684
    );
  mac_control_Mmux_n0017_Result_16_32 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0076,
      ADR1 => mac_control_txf_cnt(16),
      ADR2 => mac_control_n0078,
      ADR3 => mac_control_phydi(16),
      O => mac_control_CHOICE2111_FROM
    );
  mac_control_Mmux_n0017_Result_21_32 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0076,
      ADR1 => mac_control_txf_cnt(21),
      ADR2 => mac_control_phydi(21),
      ADR3 => mac_control_n0078,
      O => mac_control_CHOICE2111_GROM
    );
  mac_control_CHOICE2111_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2111_FROM,
      O => mac_control_CHOICE2111
    );
  mac_control_CHOICE2111_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2111_GROM,
      O => mac_control_CHOICE2159
    );
  mac_control_lmacaddr_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_25_FFX_RST,
      O => mac_control_lmacaddr(25)
    );
  mac_control_lmacaddr_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_25_FFX_RST
    );
  mac_control_Mmux_n0017_Result_13_40 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(13),
      ADR1 => mac_control_n0080,
      ADR2 => mac_control_txfifowerr_cnt(13),
      ADR3 => mac_control_n0079,
      O => mac_control_CHOICE2704_FROM
    );
  mac_control_Mmux_n0017_Result_13_94_SW0_2_1654 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_CHOICE2707,
      ADR2 => mac_control_CHOICE2699,
      ADR3 => mac_control_CHOICE2704,
      O => mac_control_CHOICE2704_GROM
    );
  mac_control_CHOICE2704_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2704_FROM,
      O => mac_control_CHOICE2704
    );
  mac_control_CHOICE2704_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2704_GROM,
      O => mac_control_Mmux_n0017_Result_13_94_SW0_2
    );
  mac_control_Mmux_n0017_Result_4_57 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0083,
      ADR1 => mac_control_rxoferr_cnt(4),
      ADR2 => mac_control_n0084,
      ADR3 => mac_control_rxcrcerr_cnt(4),
      O => mac_control_CHOICE2618_FROM
    );
  mac_control_Mmux_n0017_Result_12_57 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cnt(12),
      ADR1 => mac_control_n0083,
      ADR2 => mac_control_n0084,
      ADR3 => mac_control_rxoferr_cnt(12),
      O => mac_control_CHOICE2618_GROM
    );
  mac_control_CHOICE2618_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2618_FROM,
      O => mac_control_CHOICE2618
    );
  mac_control_CHOICE2618_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2618_GROM,
      O => mac_control_CHOICE2680
    );
  mac_control_Mmux_n0017_Result_9_17 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0078,
      ADR1 => mac_control_txf_cnt(9),
      ADR2 => mac_control_n0077,
      ADR3 => mac_control_phydo(9),
      O => mac_control_CHOICE2637_FROM
    );
  mac_control_Mmux_n0017_Result_13_17 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cnt(13),
      ADR1 => mac_control_n0078,
      ADR2 => mac_control_n0077,
      ADR3 => mac_control_phydo(13),
      O => mac_control_CHOICE2637_GROM
    );
  mac_control_CHOICE2637_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2637_FROM,
      O => mac_control_CHOICE2637
    );
  mac_control_CHOICE2637_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2637_GROM,
      O => mac_control_CHOICE2699
    );
  mac_control_Mmux_n0017_Result_8_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_N52118,
      ADR1 => mac_control_rxoferr_cnt(8),
      ADR2 => mac_control_rxf_cnt(8),
      ADR3 => mac_control_N52111,
      O => mac_control_CHOICE2385_FROM
    );
  mac_control_Mmux_n0017_Result_14_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxoferr_cnt(14),
      ADR1 => mac_control_rxf_cnt(14),
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_N52118,
      O => mac_control_CHOICE2385_GROM
    );
  mac_control_CHOICE2385_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2385_FROM,
      O => mac_control_CHOICE2385
    );
  mac_control_CHOICE2385_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2385_GROM,
      O => mac_control_CHOICE2461
    );
  mac_control_Mmux_n0017_Result_30_12 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxoferr_cnt(30),
      ADR1 => mac_control_n0083,
      ADR2 => mac_control_rxphyerr_cnt(30),
      ADR3 => mac_control_n0082,
      O => mac_control_CHOICE2057_FROM
    );
  mac_control_Mmux_n0017_Result_30_66_1_1655 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => mac_control_CHOICE2054,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2057,
      O => mac_control_CHOICE2057_GROM
    );
  mac_control_CHOICE2057_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2057_FROM,
      O => mac_control_CHOICE2057
    );
  mac_control_CHOICE2057_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2057_GROM,
      O => mac_control_Mmux_n0017_Result_30_66_1
    );
  mac_control_Mmux_n0017_Result_22_12 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0083,
      ADR1 => mac_control_rxoferr_cnt(22),
      ADR2 => mac_control_rxphyerr_cnt(22),
      ADR3 => mac_control_n0082,
      O => mac_control_CHOICE1965_FROM
    );
  mac_control_Mmux_n0017_Result_22_66_1_1656 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => mac_control_CHOICE1962,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE1965,
      O => mac_control_CHOICE1965_GROM
    );
  mac_control_CHOICE1965_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1965_FROM,
      O => mac_control_CHOICE1965
    );
  mac_control_CHOICE1965_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1965_GROM,
      O => mac_control_Mmux_n0017_Result_22_66_1
    );
  mac_control_Mmux_n0017_Result_16_37 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(16),
      ADR1 => mac_control_n0080,
      ADR2 => mac_control_txfifowerr_cnt(16),
      ADR3 => mac_control_n0079,
      O => mac_control_CHOICE2114_FROM
    );
  mac_control_Mmux_n0017_Result_21_37 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0079,
      ADR1 => mac_control_n0080,
      ADR2 => mac_control_txfifowerr_cnt(21),
      ADR3 => mac_control_rxf_cnt(21),
      O => mac_control_CHOICE2114_GROM
    );
  mac_control_CHOICE2114_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2114_FROM,
      O => mac_control_CHOICE2114
    );
  mac_control_CHOICE2114_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2114_GROM,
      O => mac_control_CHOICE2162
    );
  mac_control_Mmux_n0017_Result_4_45 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0082,
      ADR1 => mac_control_n0081,
      ADR2 => mac_control_rxfifowerr_cnt(4),
      ADR3 => mac_control_rxphyerr_cnt(4),
      O => mac_control_CHOICE2614_FROM
    );
  mac_control_Mmux_n0017_Result_13_45 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(13),
      ADR1 => mac_control_rxfifowerr_cnt(13),
      ADR2 => mac_control_n0082,
      ADR3 => mac_control_n0081,
      O => mac_control_CHOICE2614_GROM
    );
  mac_control_CHOICE2614_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2614_FROM,
      O => mac_control_CHOICE2614
    );
  mac_control_CHOICE2614_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2614_GROM,
      O => mac_control_CHOICE2707
    );
  mac_control_Mmux_n0017_Result_12_94 : X_LUT4
    generic map(
      INIT => X"F0E0"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_12_94_1,
      ADR1 => mac_control_CHOICE2684,
      ADR2 => mac_control_N52163,
      ADR3 => mac_control_Mmux_n0017_Result_12_94_SW0_2,
      O => mac_control_dout_12_FROM
    );
  mac_control_Mmux_n0017_Result_12_105 : X_LUT4
    generic map(
      INIT => X"FF0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_dout(11),
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_CHOICE2687,
      O => mac_control_N78899
    );
  mac_control_dout_12_XUSED : X_BUF
    port map (
      I => mac_control_dout_12_FROM,
      O => mac_control_CHOICE2687
    );
  mac_control_Mmux_n0017_Result_13_62 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0085,
      ADR1 => mac_control_n0086,
      ADR2 => mac_control_lmacaddr(29),
      ADR3 => mac_control_lmacaddr(13),
      O => mac_control_CHOICE2714_FROM
    );
  mac_control_Mmux_n0017_Result_13_63 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_CHOICE2711,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2714,
      O => mac_control_CHOICE2714_GROM
    );
  mac_control_CHOICE2714_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2714_FROM,
      O => mac_control_CHOICE2714
    );
  mac_control_CHOICE2714_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2714_GROM,
      O => mac_control_CHOICE2715
    );
  mac_control_Mmux_n0017_Result_21_47 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => mac_control_n0073,
      ADR1 => mac_control_N52081,
      ADR2 => mac_control_phystat(21),
      ADR3 => mac_control_N81813,
      O => mac_control_dout_21_FROM
    );
  mac_control_Mmux_n0017_Result_21_80 : X_LUT4
    generic map(
      INIT => X"DDD5"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_21_80_1,
      ADR1 => mac_control_N52163,
      ADR2 => mac_control_Mmux_n0017_Result_21_69_1,
      ADR3 => mac_control_CHOICE2164,
      O => mac_control_N76020
    );
  mac_control_dout_21_XUSED : X_BUF
    port map (
      I => mac_control_dout_21_FROM,
      O => mac_control_CHOICE2164
    );
  mac_control_lmacaddr_35 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_35_FFX_RST,
      O => mac_control_lmacaddr(35)
    );
  mac_control_lmacaddr_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_35_FFX_RST
    );
  mac_control_Mmux_n0017_Result_8_31 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cnt(8),
      ADR1 => mac_control_N52118,
      ADR2 => mac_control_phydi(8),
      ADR3 => mac_control_N52132,
      O => mac_control_CHOICE2391_FROM
    );
  mac_control_Mmux_n0017_Result_14_31 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_N52118,
      ADR1 => mac_control_phydi(14),
      ADR2 => mac_control_N52132,
      ADR3 => mac_control_txf_cnt(14),
      O => mac_control_CHOICE2391_GROM
    );
  mac_control_CHOICE2391_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2391_FROM,
      O => mac_control_CHOICE2391
    );
  mac_control_CHOICE2391_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2391_GROM,
      O => mac_control_CHOICE2467
    );
  mac_control_Mmux_n0017_Result_30_42 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2067,
      ADR1 => mac_control_Mmux_n0017_Result_30_42_1,
      ADR2 => mac_control_Mmux_n0017_Result_30_42_SW0_1,
      ADR3 => mac_control_CHOICE2064,
      O => mac_control_dout_30_FROM
    );
  mac_control_Mmux_n0017_Result_30_77 : X_LUT4
    generic map(
      INIT => X"F5D5"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_30_77_1,
      ADR1 => mac_control_Mmux_n0017_Result_30_66_1,
      ADR2 => mac_control_N52163,
      ADR3 => mac_control_CHOICE2069,
      O => mac_control_N75537
    );
  mac_control_dout_30_XUSED : X_BUF
    port map (
      I => mac_control_dout_30_FROM,
      O => mac_control_CHOICE2069
    );
  mac_control_Mmux_n0017_Result_18_34 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0078,
      ADR1 => mac_control_rxf_cnt(18),
      ADR2 => mac_control_n0079,
      ADR3 => mac_control_txf_cnt(18),
      O => mac_control_CHOICE1929_FROM
    );
  mac_control_Mmux_n0017_Result_30_34 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cnt(30),
      ADR1 => mac_control_n0078,
      ADR2 => mac_control_n0079,
      ADR3 => mac_control_rxf_cnt(30),
      O => mac_control_CHOICE1929_GROM
    );
  mac_control_CHOICE1929_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1929_FROM,
      O => mac_control_CHOICE1929
    );
  mac_control_CHOICE1929_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1929_GROM,
      O => mac_control_CHOICE2067
    );
  mac_control_Mmux_n0017_Result_22_42 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_22_42_1,
      ADR1 => mac_control_CHOICE1972,
      ADR2 => mac_control_CHOICE1975,
      ADR3 => mac_control_Mmux_n0017_Result_22_42_SW0_1,
      O => mac_control_dout_22_FROM
    );
  mac_control_Mmux_n0017_Result_22_77 : X_LUT4
    generic map(
      INIT => X"F5D5"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_22_77_1,
      ADR1 => mac_control_Mmux_n0017_Result_22_66_1,
      ADR2 => mac_control_N52163,
      ADR3 => mac_control_CHOICE1977,
      O => mac_control_N75069
    );
  mac_control_dout_22_XUSED : X_BUF
    port map (
      I => mac_control_dout_22_FROM,
      O => mac_control_CHOICE1977
    );
  mac_control_Mmux_n0017_Result_25_34 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cnt(25),
      ADR1 => mac_control_n0078,
      ADR2 => mac_control_n0079,
      ADR3 => mac_control_rxf_cnt(25),
      O => mac_control_CHOICE1998_FROM
    );
  mac_control_Mmux_n0017_Result_22_34 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0078,
      ADR1 => mac_control_rxf_cnt(22),
      ADR2 => mac_control_txf_cnt(22),
      ADR3 => mac_control_n0079,
      O => mac_control_CHOICE1998_GROM
    );
  mac_control_CHOICE1998_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1998_FROM,
      O => mac_control_CHOICE1998
    );
  mac_control_CHOICE1998_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1998_GROM,
      O => mac_control_CHOICE1975
    );
  mac_control_Mmux_n0017_Result_28_34 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(28),
      ADR1 => mac_control_n0078,
      ADR2 => mac_control_n0079,
      ADR3 => mac_control_txf_cnt(28),
      O => mac_control_CHOICE2044_FROM
    );
  mac_control_Mmux_n0017_Result_15_20 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0079,
      ADR1 => mac_control_rxf_cnt(15),
      ADR2 => mac_control_n0078,
      ADR3 => mac_control_txf_cnt(15),
      O => mac_control_CHOICE2044_GROM
    );
  mac_control_CHOICE2044_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2044_FROM,
      O => mac_control_CHOICE2044
    );
  mac_control_CHOICE2044_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2044_GROM,
      O => mac_control_CHOICE2889
    );
  mac_control_Mmux_n0017_Result_18_29 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_phystat(18),
      ADR1 => mac_control_n0076,
      ADR2 => mac_control_n0073,
      ADR3 => mac_control_phydi(18),
      O => mac_control_CHOICE1926_FROM
    );
  mac_control_Mmux_n0017_Result_22_29 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phydi(22),
      ADR1 => mac_control_n0076,
      ADR2 => mac_control_n0073,
      ADR3 => mac_control_phystat(22),
      O => mac_control_CHOICE1926_GROM
    );
  mac_control_CHOICE1926_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1926_FROM,
      O => mac_control_CHOICE1926
    );
  mac_control_CHOICE1926_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1926_GROM,
      O => mac_control_CHOICE1972
    );
  mac_control_Mmux_n0017_Result_15_30 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_N81757,
      ADR1 => mac_control_phystat(15),
      ADR2 => mac_control_n0073,
      ADR3 => mac_control_n0074,
      O => mac_control_dout_15_FROM
    );
  mac_control_Mmux_n0017_Result_15_108 : X_LUT4
    generic map(
      INIT => X"FCF8"
    )
    port map (
      ADR0 => mac_control_CHOICE2906,
      ADR1 => mac_control_N52163,
      ADR2 => mac_control_N82001,
      ADR3 => mac_control_CHOICE2891,
      O => mac_control_N80026
    );
  mac_control_dout_15_XUSED : X_BUF
    port map (
      I => mac_control_dout_15_FROM,
      O => mac_control_CHOICE2891
    );
  mac_control_Mmux_n0017_Result_13_94 : X_LUT4
    generic map(
      INIT => X"CCC8"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_13_94_1,
      ADR1 => mac_control_N52163,
      ADR2 => mac_control_Mmux_n0017_Result_13_94_SW0_2,
      ADR3 => mac_control_CHOICE2715,
      O => mac_control_dout_13_FROM
    );
  mac_control_Mmux_n0017_Result_13_105 : X_LUT4
    generic map(
      INIT => X"FF44"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_dout(12),
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2718,
      O => mac_control_N79056
    );
  mac_control_dout_13_XUSED : X_BUF
    port map (
      I => mac_control_dout_13_FROM,
      O => mac_control_CHOICE2718
    );
  mac_control_Mmux_n0017_Result_14_39 : X_LUT4
    generic map(
      INIT => X"EC00"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(14),
      ADR1 => mac_control_CHOICE2467,
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_N52220,
      O => mac_control_CHOICE2469_FROM
    );
  mac_control_Mmux_n0017_Result_14_45 : X_LUT4
    generic map(
      INIT => X"FFE0"
    )
    port map (
      ADR0 => mac_control_CHOICE2461,
      ADR1 => mac_control_CHOICE2458,
      ADR2 => mac_control_N52228,
      ADR3 => mac_control_CHOICE2469,
      O => mac_control_CHOICE2469_GROM
    );
  mac_control_CHOICE2469_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2469_FROM,
      O => mac_control_CHOICE2469
    );
  mac_control_CHOICE2469_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2469_GROM,
      O => mac_control_CHOICE2470
    );
  mac_control_Mmux_n0017_Result_25_29 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phydi(25),
      ADR1 => mac_control_n0076,
      ADR2 => mac_control_phystat(25),
      ADR3 => mac_control_n0073,
      O => mac_control_CHOICE1995_FROM
    );
  mac_control_Mmux_n0017_Result_15_15 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phydi(15),
      ADR1 => mac_control_phydo(15),
      ADR2 => mac_control_n0077,
      ADR3 => mac_control_n0076,
      O => mac_control_CHOICE1995_GROM
    );
  mac_control_CHOICE1995_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1995_FROM,
      O => mac_control_CHOICE1995
    );
  mac_control_CHOICE1995_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1995_GROM,
      O => mac_control_CHOICE2886
    );
  mac_control_lmacaddr_43 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_43_FFX_RST,
      O => mac_control_lmacaddr(43)
    );
  mac_control_lmacaddr_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_43_FFX_RST
    );
  tx_output_crc_loigc_Mxor_CO_13_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(0),
      ADR1 => tx_output_data(4),
      ADR2 => tx_output_crcl(31),
      ADR3 => tx_output_crcl(27),
      O => tx_output_crcl_19_FROM
    );
  tx_output_n0034_19_1 : X_LUT4
    generic map(
      INIT => X"AFFA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => VCC,
      ADR2 => tx_output_crcl(11),
      ADR3 => tx_output_crc_loigc_Mxor_CO_13_Xo(2),
      O => tx_output_n0034(19)
    );
  tx_output_crcl_19_XUSED : X_BUF
    port map (
      I => tx_output_crcl_19_FROM,
      O => tx_output_crc_loigc_Mxor_CO_13_Xo(2)
    );
  mac_control_Mmux_n0017_Result_0_114 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => mac_control_N52244,
      ADR1 => mac_control_CHOICE2223,
      ADR2 => mac_control_CHOICE2210,
      ADR3 => mac_control_CHOICE2216,
      O => mac_control_dout_0_FROM
    );
  mac_control_Mmux_n0017_Result_0_137 : X_LUT4
    generic map(
      INIT => X"CCC8"
    )
    port map (
      ADR0 => mac_control_N52081,
      ADR1 => mac_control_N52163,
      ADR2 => mac_control_CHOICE2206,
      ADR3 => mac_control_CHOICE2224,
      O => mac_control_N76337
    );
  mac_control_dout_0_XUSED : X_BUF
    port map (
      I => mac_control_dout_0_FROM,
      O => mac_control_CHOICE2224
    );
  mac_control_Mmux_n0017_Result_6_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_N52118,
      ADR1 => mac_control_rxf_cnt(6),
      ADR2 => mac_control_rxoferr_cnt(6),
      ADR3 => mac_control_N52111,
      O => mac_control_CHOICE2309_FROM
    );
  mac_control_Mmux_n0017_Result_31_44 : X_LUT4
    generic map(
      INIT => X"FAF8"
    )
    port map (
      ADR0 => mac_control_N52111,
      ADR1 => mac_control_CHOICE1805,
      ADR2 => mac_control_CHOICE1813,
      ADR3 => mac_control_CHOICE1802,
      O => mac_control_CHOICE2309_GROM
    );
  mac_control_CHOICE2309_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2309_FROM,
      O => mac_control_CHOICE2309
    );
  mac_control_CHOICE2309_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2309_GROM,
      O => mac_control_CHOICE1814
    );
  mac_control_Mmux_n0017_Result_16_12 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxoferr_cnt(16),
      ADR1 => mac_control_rxcrcerr_cnt(16),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_n0084,
      O => mac_control_CHOICE2103_FROM
    );
  mac_control_Mmux_n0017_Result_16_69_1_1657 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => mac_control_CHOICE2100,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2103,
      O => mac_control_CHOICE2103_GROM
    );
  mac_control_CHOICE2103_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2103_FROM,
      O => mac_control_CHOICE2103
    );
  mac_control_CHOICE2103_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2103_GROM,
      O => mac_control_Mmux_n0017_Result_16_69_1
    );
  mac_control_Mmux_n0017_Result_1_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_N52118,
      ADR1 => mac_control_rxf_cnt(1),
      ADR2 => mac_control_rxoferr_cnt(1),
      ADR3 => mac_control_N52111,
      O => mac_control_CHOICE2233_FROM
    );
  mac_control_Mmux_n0017_Result_23_44 : X_LUT4
    generic map(
      INIT => X"FAEA"
    )
    port map (
      ADR0 => mac_control_CHOICE1869,
      ADR1 => mac_control_CHOICE1861,
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_CHOICE1858,
      O => mac_control_CHOICE2233_GROM
    );
  mac_control_CHOICE2233_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2233_FROM,
      O => mac_control_CHOICE2233
    );
  mac_control_CHOICE2233_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2233_GROM,
      O => mac_control_CHOICE1870
    );
  mac_control_Mmux_n0017_Result_15_60 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0084,
      ADR1 => mac_control_rxcrcerr_cnt(15),
      ADR2 => mac_control_n0085,
      ADR3 => mac_control_lmacaddr(15),
      O => mac_control_CHOICE2901_FROM
    );
  mac_control_Mmux_n0017_Result_15_74_SW0 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(15),
      ADR1 => mac_control_n0081,
      ADR2 => mac_control_CHOICE2904,
      ADR3 => mac_control_CHOICE2901,
      O => mac_control_CHOICE2901_GROM
    );
  mac_control_CHOICE2901_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2901_FROM,
      O => mac_control_CHOICE2901
    );
  mac_control_CHOICE2901_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2901_GROM,
      O => mac_control_N81745
    );
  mac_control_Mmux_n0017_Result_24_12 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0084,
      ADR1 => mac_control_rxcrcerr_cnt(24),
      ADR2 => mac_control_rxoferr_cnt(24),
      ADR3 => mac_control_n0083,
      O => mac_control_CHOICE2175_FROM
    );
  mac_control_Mmux_n0017_Result_24_69_1_1658 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_CHOICE2172,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2175,
      O => mac_control_CHOICE2175_GROM
    );
  mac_control_CHOICE2175_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2175_FROM,
      O => mac_control_CHOICE2175
    );
  mac_control_CHOICE2175_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2175_GROM,
      O => mac_control_Mmux_n0017_Result_24_69_1
    );
  mac_control_Mmux_n0017_Result_5_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_N52111,
      ADR1 => mac_control_rxoferr_cnt(5),
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_rxf_cnt(5),
      O => mac_control_CHOICE2347_FROM
    );
  mac_control_Mmux_n0017_Result_14_69 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cnt(14),
      ADR1 => mac_control_N52118,
      ADR2 => mac_control_txfifowerr_cnt(14),
      ADR3 => mac_control_N52111,
      O => mac_control_CHOICE2347_GROM
    );
  mac_control_CHOICE2347_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2347_FROM,
      O => mac_control_CHOICE2347
    );
  mac_control_CHOICE2347_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2347_GROM,
      O => mac_control_CHOICE2474
    );
  mac_control_Mmux_n0017_Result_0_85 : X_LUT4
    generic map(
      INIT => X"E040"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => mac_control_lmacaddr(16),
      ADR2 => mac_control_N52143,
      ADR3 => mac_control_lmacaddr(32),
      O => mac_control_CHOICE2216_FROM
    );
  mac_control_Mmux_n0017_Result_14_86 : X_LUT4
    generic map(
      INIT => X"88C0"
    )
    port map (
      ADR0 => mac_control_lmacaddr(46),
      ADR1 => mac_control_N52143,
      ADR2 => mac_control_lmacaddr(30),
      ADR3 => mac_control_addr(0),
      O => mac_control_CHOICE2216_GROM
    );
  mac_control_CHOICE2216_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2216_FROM,
      O => mac_control_CHOICE2216
    );
  mac_control_CHOICE2216_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2216_GROM,
      O => mac_control_CHOICE2480
    );
  mac_control_Mmux_n0017_Result_17_32 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0078,
      ADR1 => mac_control_phydi(17),
      ADR2 => mac_control_txf_cnt(17),
      ADR3 => mac_control_n0076,
      O => mac_control_CHOICE2135_FROM
    );
  mac_control_Mmux_n0017_Result_24_32 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0076,
      ADR1 => mac_control_n0078,
      ADR2 => mac_control_phydi(24),
      ADR3 => mac_control_txf_cnt(24),
      O => mac_control_CHOICE2135_GROM
    );
  mac_control_CHOICE2135_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2135_FROM,
      O => mac_control_CHOICE2135
    );
  mac_control_CHOICE2135_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2135_GROM,
      O => mac_control_CHOICE2183
    );
  mac_control_Mmux_n0017_Result_9_57 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0084,
      ADR1 => mac_control_rxoferr_cnt(9),
      ADR2 => mac_control_rxcrcerr_cnt(9),
      ADR3 => mac_control_n0083,
      O => mac_control_CHOICE2649_FROM
    );
  mac_control_Mmux_n0017_Result_15_48 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0082,
      ADR1 => mac_control_rxoferr_cnt(15),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_rxphyerr_cnt(15),
      O => mac_control_CHOICE2649_GROM
    );
  mac_control_CHOICE2649_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2649_FROM,
      O => mac_control_CHOICE2649
    );
  mac_control_CHOICE2649_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2649_GROM,
      O => mac_control_CHOICE2897
    );
  mac_control_lmacaddr_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_19_FFX_RST,
      O => mac_control_lmacaddr(19)
    );
  mac_control_lmacaddr_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_19_FFX_RST
    );
  mac_control_Mmux_n0017_Result_19_9 : X_LUT4
    generic map(
      INIT => X"A280"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_rxcrcerr_cnt(19),
      ADR3 => mac_control_rxoferr_cnt(19),
      O => mac_control_CHOICE1833_FROM
    );
  mac_control_Mmux_n0017_Result_31_57 : X_LUT4
    generic map(
      INIT => X"0D08"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => mac_control_phydi(31),
      ADR2 => mac_control_addr(1),
      ADR3 => mac_control_phyaddr(31),
      O => mac_control_CHOICE1833_GROM
    );
  mac_control_CHOICE1833_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1833_FROM,
      O => mac_control_CHOICE1833
    );
  mac_control_CHOICE1833_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1833_GROM,
      O => mac_control_CHOICE1817
    );
  mac_control_Mmux_n0017_Result_19_4 : X_LUT4
    generic map(
      INIT => X"4450"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_rxphyerr_cnt(19),
      ADR2 => mac_control_rxfifowerr_cnt(19),
      ADR3 => mac_control_addr(0),
      O => mac_control_CHOICE1830_FROM
    );
  mac_control_Mmux_n0017_Result_23_57 : X_LUT4
    generic map(
      INIT => X"5044"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_phyaddr(23),
      ADR2 => mac_control_phydi(23),
      ADR3 => mac_control_addr(0),
      O => mac_control_CHOICE1830_GROM
    );
  mac_control_CHOICE1830_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1830_FROM,
      O => mac_control_CHOICE1830
    );
  mac_control_CHOICE1830_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1830_GROM,
      O => mac_control_CHOICE1873
    );
  mac_control_Mmux_n0017_Result_8_86 : X_LUT4
    generic map(
      INIT => X"B080"
    )
    port map (
      ADR0 => mac_control_lmacaddr(40),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_N52143,
      ADR3 => mac_control_lmacaddr(24),
      O => mac_control_CHOICE2404_FROM
    );
  mac_control_Mmux_n0017_Result_15_65 : X_LUT4
    generic map(
      INIT => X"B080"
    )
    port map (
      ADR0 => mac_control_lmacaddr(47),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_N52143,
      ADR3 => mac_control_lmacaddr(31),
      O => mac_control_CHOICE2404_GROM
    );
  mac_control_CHOICE2404_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2404_FROM,
      O => mac_control_CHOICE2404
    );
  mac_control_CHOICE2404_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2404_GROM,
      O => mac_control_CHOICE2904
    );
  mac_control_Mmux_n0017_Result_29_7 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(29),
      ADR1 => mac_control_rxfifowerr_cnt(29),
      ADR2 => mac_control_n0081,
      ADR3 => mac_control_n0080,
      O => mac_control_CHOICE2077_FROM
    );
  mac_control_Mmux_n0017_Result_15_74 : X_LUT4
    generic map(
      INIT => X"FEFC"
    )
    port map (
      ADR0 => mac_control_n0080,
      ADR1 => mac_control_N81745,
      ADR2 => mac_control_CHOICE2897,
      ADR3 => mac_control_txfifowerr_cnt(15),
      O => mac_control_CHOICE2077_GROM
    );
  mac_control_CHOICE2077_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2077_FROM,
      O => mac_control_CHOICE2077
    );
  mac_control_CHOICE2077_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2077_GROM,
      O => mac_control_CHOICE2906
    );
  mac_control_Mmux_n0017_Result_27_67 : X_LUT4
    generic map(
      INIT => X"8880"
    )
    port map (
      ADR0 => mac_control_N52125,
      ADR1 => mac_control_addr(1),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_phystat(27),
      O => mac_control_CHOICE1905_FROM
    );
  mac_control_Mmux_n0017_Result_23_67 : X_LUT4
    generic map(
      INIT => X"C080"
    )
    port map (
      ADR0 => mac_control_phystat(23),
      ADR1 => mac_control_N52125,
      ADR2 => mac_control_addr(1),
      ADR3 => mac_control_addr(0),
      O => mac_control_CHOICE1905_GROM
    );
  mac_control_CHOICE1905_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1905_FROM,
      O => mac_control_CHOICE1905
    );
  mac_control_CHOICE1905_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1905_GROM,
      O => mac_control_CHOICE1877
    );
  tx_output_crc_loigc_Mxor_CO_13_Xo_5_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_Mxor_CO_18_Xo(0),
      ADR1 => tx_output_crc_loigc_Mxor_n0007_Xo(0),
      ADR2 => tx_output_crc_loigc_Mxor_CO_13_Xo(2),
      ADR3 => tx_output_crcl(5),
      O => tx_output_crcl_13_FROM
    );
  tx_output_n0034_13_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crc_13_Q,
      O => tx_output_n0034(13)
    );
  tx_output_crcl_13_XUSED : X_BUF
    port map (
      I => tx_output_crcl_13_FROM,
      O => tx_output_crc_13_Q
    );
  mac_control_Mmux_n0017_Result_17_12 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0083,
      ADR1 => mac_control_rxcrcerr_cnt(17),
      ADR2 => mac_control_rxoferr_cnt(17),
      ADR3 => mac_control_n0084,
      O => mac_control_CHOICE2127_FROM
    );
  mac_control_Mmux_n0017_Result_17_69_1_1659 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_CHOICE2124,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2127,
      O => mac_control_CHOICE2127_GROM
    );
  mac_control_CHOICE2127_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2127_FROM,
      O => mac_control_CHOICE2127
    );
  mac_control_CHOICE2127_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2127_GROM,
      O => mac_control_Mmux_n0017_Result_17_69_1
    );
  mac_control_Mmux_n0017_Result_25_12 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0082,
      ADR1 => mac_control_rxoferr_cnt(25),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_rxphyerr_cnt(25),
      O => mac_control_CHOICE1988_FROM
    );
  mac_control_Mmux_n0017_Result_25_66_1_1660 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => mac_control_CHOICE1985,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE1988,
      O => mac_control_CHOICE1988_GROM
    );
  mac_control_CHOICE1988_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1988_FROM,
      O => mac_control_CHOICE1988
    );
  mac_control_CHOICE1988_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1988_GROM,
      O => mac_control_Mmux_n0017_Result_25_66_1
    );
  mac_control_Mmux_n0017_Result_17_37 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(17),
      ADR1 => mac_control_n0079,
      ADR2 => mac_control_n0080,
      ADR3 => mac_control_rxf_cnt(17),
      O => mac_control_CHOICE2138_FROM
    );
  mac_control_Mmux_n0017_Result_24_37 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0080,
      ADR1 => mac_control_n0079,
      ADR2 => mac_control_rxf_cnt(24),
      ADR3 => mac_control_txfifowerr_cnt(24),
      O => mac_control_CHOICE2138_GROM
    );
  mac_control_CHOICE2138_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2138_FROM,
      O => mac_control_CHOICE2138
    );
  mac_control_CHOICE2138_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2138_GROM,
      O => mac_control_CHOICE2186
    );
  mac_control_Mmux_n0017_Result_16_47 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_phystat(16),
      ADR1 => mac_control_n0073,
      ADR2 => mac_control_N81793,
      ADR3 => mac_control_N52081,
      O => mac_control_dout_16_FROM
    );
  mac_control_Mmux_n0017_Result_16_80 : X_LUT4
    generic map(
      INIT => X"DDD5"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_16_80_1,
      ADR1 => mac_control_N52163,
      ADR2 => mac_control_Mmux_n0017_Result_16_69_1,
      ADR3 => mac_control_CHOICE2116,
      O => mac_control_N75776
    );
  mac_control_dout_16_XUSED : X_BUF
    port map (
      I => mac_control_dout_16_FROM,
      O => mac_control_CHOICE2116
    );
  mac_control_Mmux_n0017_Result_24_47 : X_LUT4
    generic map(
      INIT => X"FEEE"
    )
    port map (
      ADR0 => mac_control_N52081,
      ADR1 => mac_control_N81789,
      ADR2 => mac_control_n0073,
      ADR3 => mac_control_phystat(24),
      O => mac_control_dout_24_FROM
    );
  mac_control_Mmux_n0017_Result_24_80 : X_LUT4
    generic map(
      INIT => X"DDD5"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_24_80_1,
      ADR1 => mac_control_N52163,
      ADR2 => mac_control_Mmux_n0017_Result_24_69_1,
      ADR3 => mac_control_CHOICE2188,
      O => mac_control_N76142
    );
  mac_control_dout_24_XUSED : X_BUF
    port map (
      I => mac_control_dout_24_FROM,
      O => mac_control_CHOICE2188
    );
  mac_control_lmacaddr_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_27_FFX_RST,
      O => mac_control_lmacaddr(27)
    );
  mac_control_lmacaddr_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_27_FFX_RST
    );
  mac_control_Mmux_n0017_Result_25_42 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE1995,
      ADR1 => mac_control_CHOICE1998,
      ADR2 => mac_control_Mmux_n0017_Result_25_42_1,
      ADR3 => mac_control_Mmux_n0017_Result_25_42_SW0_1,
      O => mac_control_dout_25_FROM
    );
  mac_control_Mmux_n0017_Result_25_77 : X_LUT4
    generic map(
      INIT => X"DDD5"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_25_77_1,
      ADR1 => mac_control_N52163,
      ADR2 => mac_control_Mmux_n0017_Result_25_66_1,
      ADR3 => mac_control_CHOICE2000,
      O => mac_control_N75186
    );
  mac_control_dout_25_XUSED : X_BUF
    port map (
      I => mac_control_dout_25_FROM,
      O => mac_control_CHOICE2000
    );
  mac_control_Mmux_n0017_Result_1_107 : X_LUT4
    generic map(
      INIT => X"8854"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => mac_control_N52125,
      ADR2 => mac_control_N82137,
      ADR3 => mac_control_addr(1),
      O => mac_control_CHOICE2258_FROM
    );
  mac_control_Mmux_n0017_Result_1_113 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_N52244,
      ADR1 => mac_control_CHOICE2246,
      ADR2 => mac_control_CHOICE2252,
      ADR3 => mac_control_CHOICE2258,
      O => mac_control_CHOICE2258_GROM
    );
  mac_control_CHOICE2258_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2258_FROM,
      O => mac_control_CHOICE2258
    );
  mac_control_CHOICE2258_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2258_GROM,
      O => mac_control_CHOICE2259
    );
  mac_control_Mmux_n0017_Result_26_12 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0082,
      ADR1 => mac_control_rxoferr_cnt(26),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_rxphyerr_cnt(26),
      O => mac_control_CHOICE2011_FROM
    );
  mac_control_Mmux_n0017_Result_26_66_1_1661 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE2008,
      ADR3 => mac_control_CHOICE2011,
      O => mac_control_CHOICE2011_GROM
    );
  mac_control_CHOICE2011_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2011_FROM,
      O => mac_control_CHOICE2011
    );
  mac_control_CHOICE2011_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2011_GROM,
      O => mac_control_Mmux_n0017_Result_26_66_1
    );
  mac_control_Mmux_n0017_Result_18_12 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(18),
      ADR1 => mac_control_rxoferr_cnt(18),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_n0082,
      O => mac_control_CHOICE1919_FROM
    );
  mac_control_Mmux_n0017_Result_18_66_1_1662 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_CHOICE1916,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE1919,
      O => mac_control_CHOICE1919_GROM
    );
  mac_control_CHOICE1919_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1919_FROM,
      O => mac_control_CHOICE1919
    );
  mac_control_CHOICE1919_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1919_GROM,
      O => mac_control_Mmux_n0017_Result_18_66_1
    );
  mac_control_Mmux_n0017_Result_17_47 : X_LUT4
    generic map(
      INIT => X"FEEE"
    )
    port map (
      ADR0 => mac_control_N81749,
      ADR1 => mac_control_N52081,
      ADR2 => mac_control_phystat(17),
      ADR3 => mac_control_n0073,
      O => mac_control_dout_17_FROM
    );
  mac_control_Mmux_n0017_Result_17_80 : X_LUT4
    generic map(
      INIT => X"CF8F"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_17_69_1,
      ADR1 => mac_control_N52163,
      ADR2 => mac_control_Mmux_n0017_Result_17_80_1,
      ADR3 => mac_control_CHOICE2140,
      O => mac_control_N75898
    );
  mac_control_dout_17_XUSED : X_BUF
    port map (
      I => mac_control_dout_17_FROM,
      O => mac_control_CHOICE2140
    );
  mac_control_Mmux_n0017_Result_18_42 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE1929,
      ADR1 => mac_control_Mmux_n0017_Result_18_42_1,
      ADR2 => mac_control_CHOICE1926,
      ADR3 => mac_control_Mmux_n0017_Result_18_42_SW0_1,
      O => mac_control_dout_18_FROM
    );
  mac_control_Mmux_n0017_Result_18_77 : X_LUT4
    generic map(
      INIT => X"F3B3"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_18_66_1,
      ADR1 => mac_control_Mmux_n0017_Result_18_77_1,
      ADR2 => mac_control_N52163,
      ADR3 => mac_control_CHOICE1931,
      O => mac_control_N74835
    );
  mac_control_dout_18_XUSED : X_BUF
    port map (
      I => mac_control_dout_18_FROM,
      O => mac_control_CHOICE1931
    );
  mac_control_Mmux_n0017_Result_26_42 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2018,
      ADR1 => mac_control_CHOICE2021,
      ADR2 => mac_control_Mmux_n0017_Result_26_42_SW0_1,
      ADR3 => mac_control_Mmux_n0017_Result_26_42_1,
      O => mac_control_dout_26_FROM
    );
  mac_control_Mmux_n0017_Result_26_77 : X_LUT4
    generic map(
      INIT => X"CF8F"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_26_66_1,
      ADR1 => mac_control_N52163,
      ADR2 => mac_control_Mmux_n0017_Result_26_77_1,
      ADR3 => mac_control_CHOICE2023,
      O => mac_control_N75303
    );
  mac_control_dout_26_XUSED : X_BUF
    port map (
      I => mac_control_dout_26_FROM,
      O => mac_control_CHOICE2023
    );
  mac_control_Mmux_n0017_Result_2_107 : X_LUT4
    generic map(
      INIT => X"8584"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_N52125,
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_N82113,
      O => mac_control_CHOICE2296_FROM
    );
  mac_control_Mmux_n0017_Result_2_113 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => mac_control_N52244,
      ADR1 => mac_control_CHOICE2290,
      ADR2 => mac_control_CHOICE2284,
      ADR3 => mac_control_CHOICE2296,
      O => mac_control_CHOICE2296_GROM
    );
  mac_control_CHOICE2296_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2296_FROM,
      O => mac_control_CHOICE2296
    );
  mac_control_CHOICE2296_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2296_GROM,
      O => mac_control_CHOICE2297
    );
  mac_control_Mmux_n0017_Result_1_69 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_N52111,
      ADR1 => mac_control_rxcrcerr_cnt(1),
      ADR2 => mac_control_txfifowerr_cnt(1),
      ADR3 => mac_control_N52118,
      O => mac_control_CHOICE2246_FROM
    );
  mac_control_Mmux_n0017_Result_27_44 : X_LUT4
    generic map(
      INIT => X"FFE0"
    )
    port map (
      ADR0 => mac_control_CHOICE1889,
      ADR1 => mac_control_CHOICE1886,
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_CHOICE1897,
      O => mac_control_CHOICE2246_GROM
    );
  mac_control_CHOICE2246_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2246_FROM,
      O => mac_control_CHOICE2246
    );
  mac_control_CHOICE2246_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2246_GROM,
      O => mac_control_CHOICE1898
    );
  mac_control_Mmux_n0017_Result_28_12 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxoferr_cnt(28),
      ADR1 => mac_control_rxphyerr_cnt(28),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_n0082,
      O => mac_control_CHOICE2034_FROM
    );
  mac_control_Mmux_n0017_Result_28_66_1_1663 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE2031,
      ADR3 => mac_control_CHOICE2034,
      O => mac_control_CHOICE2034_GROM
    );
  mac_control_CHOICE2034_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2034_FROM,
      O => mac_control_CHOICE2034
    );
  mac_control_CHOICE2034_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2034_GROM,
      O => mac_control_Mmux_n0017_Result_28_66_1
    );
  mac_control_Mmux_n0017_Result_5_69 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(5),
      ADR1 => mac_control_rxcrcerr_cnt(5),
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_N52118,
      O => mac_control_CHOICE2360_FROM
    );
  mac_control_Mmux_n0017_Result_19_44 : X_LUT4
    generic map(
      INIT => X"FAF8"
    )
    port map (
      ADR0 => mac_control_N52111,
      ADR1 => mac_control_CHOICE1830,
      ADR2 => mac_control_CHOICE1841,
      ADR3 => mac_control_CHOICE1833,
      O => mac_control_CHOICE2360_GROM
    );
  mac_control_CHOICE2360_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2360_FROM,
      O => mac_control_CHOICE2360
    );
  mac_control_CHOICE2360_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2360_GROM,
      O => mac_control_CHOICE1842
    );
  mac_control_lmacaddr_37 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_37_FFX_RST,
      O => mac_control_lmacaddr(37)
    );
  mac_control_lmacaddr_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_37_FFX_RST
    );
  mac_control_Mmux_n0017_Result_31_9 : X_LUT4
    generic map(
      INIT => X"C480"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => mac_control_addr(1),
      ADR2 => mac_control_rxcrcerr_cnt(31),
      ADR3 => mac_control_rxoferr_cnt(31),
      O => mac_control_CHOICE1805_FROM
    );
  mac_control_Mmux_n0017_Result_27_57 : X_LUT4
    generic map(
      INIT => X"00CA"
    )
    port map (
      ADR0 => mac_control_phyaddr(27),
      ADR1 => mac_control_phydi(27),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_addr(1),
      O => mac_control_CHOICE1805_GROM
    );
  mac_control_CHOICE1805_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1805_FROM,
      O => mac_control_CHOICE1805
    );
  mac_control_CHOICE1805_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1805_GROM,
      O => mac_control_CHOICE1901
    );
  mac_control_Mmux_n0017_Result_31_4 : X_LUT4
    generic map(
      INIT => X"0D08"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => mac_control_rxphyerr_cnt(31),
      ADR2 => mac_control_addr(1),
      ADR3 => mac_control_rxfifowerr_cnt(31),
      O => mac_control_CHOICE1802_FROM
    );
  mac_control_Mmux_n0017_Result_19_57 : X_LUT4
    generic map(
      INIT => X"0E02"
    )
    port map (
      ADR0 => mac_control_phyaddr(19),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_addr(1),
      ADR3 => mac_control_phydi(19),
      O => mac_control_CHOICE1802_GROM
    );
  mac_control_CHOICE1802_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1802_FROM,
      O => mac_control_CHOICE1802
    );
  mac_control_CHOICE1802_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1802_GROM,
      O => mac_control_CHOICE1845
    );
  mac_control_Mmux_n0017_Result_28_42 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2044,
      ADR1 => mac_control_Mmux_n0017_Result_28_42_SW0_1,
      ADR2 => mac_control_CHOICE2041,
      ADR3 => mac_control_Mmux_n0017_Result_28_42_1,
      O => mac_control_dout_28_FROM
    );
  mac_control_Mmux_n0017_Result_28_77 : X_LUT4
    generic map(
      INIT => X"F3B3"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_28_66_1,
      ADR1 => mac_control_Mmux_n0017_Result_28_77_1,
      ADR2 => mac_control_N52163,
      ADR3 => mac_control_CHOICE2046,
      O => mac_control_N75420
    );
  mac_control_dout_28_XUSED : X_BUF
    port map (
      I => mac_control_dout_28_FROM,
      O => mac_control_CHOICE2046
    );
  mac_control_Mmux_n0017_Result_27_9 : X_LUT4
    generic map(
      INIT => X"A808"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_rxoferr_cnt(27),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_rxcrcerr_cnt(27),
      O => mac_control_CHOICE1889_FROM
    );
  mac_control_Mmux_n0017_Result_19_67 : X_LUT4
    generic map(
      INIT => X"E000"
    )
    port map (
      ADR0 => mac_control_phystat(19),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_N52125,
      ADR3 => mac_control_addr(1),
      O => mac_control_CHOICE1889_GROM
    );
  mac_control_CHOICE1889_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1889_FROM,
      O => mac_control_CHOICE1889
    );
  mac_control_CHOICE1889_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1889_GROM,
      O => mac_control_CHOICE1849
    );
  mac_control_Mmux_n0017_Result_29_12 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0082,
      ADR1 => mac_control_rxoferr_cnt(29),
      ADR2 => mac_control_n0083,
      ADR3 => mac_control_rxphyerr_cnt(29),
      O => mac_control_CHOICE2080_FROM
    );
  mac_control_Mmux_n0017_Result_29_66_1_1664 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_CHOICE2077,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2080,
      O => mac_control_CHOICE2080_GROM
    );
  mac_control_CHOICE2080_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2080_FROM,
      O => mac_control_CHOICE2080
    );
  mac_control_CHOICE2080_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2080_GROM,
      O => mac_control_Mmux_n0017_Result_29_66_1
    );
  mac_control_Mmux_n0017_Result_29_29 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0073,
      ADR1 => mac_control_phydi(29),
      ADR2 => mac_control_n0076,
      ADR3 => mac_control_phystat(29),
      O => mac_control_CHOICE2087_FROM
    );
  mac_control_Mmux_n0017_Result_28_29 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phydi(28),
      ADR1 => mac_control_n0076,
      ADR2 => mac_control_phystat(28),
      ADR3 => mac_control_n0073,
      O => mac_control_CHOICE2087_GROM
    );
  mac_control_CHOICE2087_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2087_FROM,
      O => mac_control_CHOICE2087
    );
  mac_control_CHOICE2087_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2087_GROM,
      O => mac_control_CHOICE2041
    );
  mac_control_Mmux_n0017_Result_29_42 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2087,
      ADR1 => mac_control_CHOICE2090,
      ADR2 => mac_control_Mmux_n0017_Result_29_42_SW0_1,
      ADR3 => mac_control_Mmux_n0017_Result_29_42_1,
      O => mac_control_dout_29_FROM
    );
  mac_control_Mmux_n0017_Result_29_77 : X_LUT4
    generic map(
      INIT => X"F5D5"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_29_77_1,
      ADR1 => mac_control_Mmux_n0017_Result_29_66_1,
      ADR2 => mac_control_N52163,
      ADR3 => mac_control_CHOICE2092,
      O => mac_control_N75654
    );
  mac_control_dout_29_XUSED : X_BUF
    port map (
      I => mac_control_dout_29_FROM,
      O => mac_control_CHOICE2092
    );
  mac_control_Mmux_n0017_Result_29_34 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(29),
      ADR1 => mac_control_n0079,
      ADR2 => mac_control_txf_cnt(29),
      ADR3 => mac_control_n0078,
      O => mac_control_CHOICE2090_GROM
    );
  mac_control_CHOICE2090_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2090_GROM,
      O => mac_control_CHOICE2090
    );
  mac_control_Mmux_n0017_Result_5_107 : X_LUT4
    generic map(
      INIT => X"C032"
    )
    port map (
      ADR0 => mac_control_N82133,
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_N52125,
      ADR3 => mac_control_addr(1),
      O => mac_control_CHOICE2372_FROM
    );
  mac_control_Mmux_n0017_Result_5_113 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_CHOICE2360,
      ADR1 => mac_control_N52244,
      ADR2 => mac_control_CHOICE2366,
      ADR3 => mac_control_CHOICE2372,
      O => mac_control_CHOICE2372_GROM
    );
  mac_control_CHOICE2372_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2372_FROM,
      O => mac_control_CHOICE2372
    );
  mac_control_CHOICE2372_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2372_GROM,
      O => mac_control_CHOICE2373
    );
  rx_input_memio_crccomb_Mxor_CO_6_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0124(0),
      ADR1 => rx_input_memio_crccomb_Mxor_n0007_Xo(0),
      ADR2 => rx_input_memio_crccomb_Mxor_CO_18_Xo(0),
      ADR3 => rx_input_memio_crccomb_n0115(0),
      O => rx_input_memio_crcl_6_FROM
    );
  rx_input_memio_n0048_6_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_6_Q,
      O => rx_input_memio_n0048(6)
    );
  rx_input_memio_crcl_6_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_6_FROM,
      O => rx_input_memio_crc_6_Q
    );
  mac_control_Mmux_n0017_Result_6_107 : X_LUT4
    generic map(
      INIT => X"8382"
    )
    port map (
      ADR0 => mac_control_N52125,
      ADR1 => mac_control_addr(1),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_N82125,
      O => mac_control_CHOICE2334_FROM
    );
  mac_control_Mmux_n0017_Result_6_113 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => mac_control_CHOICE2322,
      ADR1 => mac_control_CHOICE2328,
      ADR2 => mac_control_N52244,
      ADR3 => mac_control_CHOICE2334,
      O => mac_control_CHOICE2334_GROM
    );
  mac_control_CHOICE2334_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2334_FROM,
      O => mac_control_CHOICE2334
    );
  mac_control_CHOICE2334_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2334_GROM,
      O => mac_control_CHOICE2335
    );
  mac_control_lmacaddr_45 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_45_FFX_RST,
      O => mac_control_lmacaddr(45)
    );
  mac_control_lmacaddr_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_45_FFX_RST
    );
  tx_output_crcsell_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_crcsell_3_CEMUXNOT
    );
  mac_control_Mmux_n0017_Result_8_107 : X_LUT4
    generic map(
      INIT => X"C00E"
    )
    port map (
      ADR0 => mac_control_N82129,
      ADR1 => mac_control_N52125,
      ADR2 => mac_control_addr(1),
      ADR3 => mac_control_addr(0),
      O => mac_control_CHOICE2410_FROM
    );
  mac_control_Mmux_n0017_Result_8_113 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => mac_control_N52244,
      ADR1 => mac_control_CHOICE2404,
      ADR2 => mac_control_CHOICE2398,
      ADR3 => mac_control_CHOICE2410,
      O => mac_control_CHOICE2410_GROM
    );
  mac_control_CHOICE2410_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2410_FROM,
      O => mac_control_CHOICE2410
    );
  mac_control_CHOICE2410_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2410_GROM,
      O => mac_control_CHOICE2411
    );
  tx_input_Ker34480137_SW0 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => tx_input_CHOICE1717,
      ADR1 => tx_input_CHOICE1702,
      ADR2 => tx_input_CHOICE1710,
      ADR3 => tx_input_CHOICE1695,
      O => tx_input_cs_FFd5_FROM
    );
  tx_input_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"EEEC"
    )
    port map (
      ADR0 => tx_input_cs_FFd6,
      ADR1 => tx_input_cs_FFd4,
      ADR2 => tx_input_Ker34480137_2,
      ADR3 => tx_input_N81681,
      O => tx_input_cs_FFd5_In
    );
  tx_input_cs_FFd5_XUSED : X_BUF
    port map (
      I => tx_input_cs_FFd5_FROM,
      O => tx_input_N81681
    );
  rx_input_RESET_1_1665 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => RESET_IBUF_2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_RESET_1_FROM
    );
  rx_input_memio_n00451 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd15,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_RESET_1,
      O => rx_input_RESET_1_GROM
    );
  rx_input_RESET_1_XUSED : X_BUF
    port map (
      I => rx_input_RESET_1_FROM,
      O => rx_input_RESET_1
    );
  rx_input_RESET_1_YUSED : X_BUF
    port map (
      I => rx_input_RESET_1_GROM,
      O => rx_input_memio_n0045
    );
  memcontroller_dnl2_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_1_CEMUXNOT
    );
  memcontroller_dnl2_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_3_CEMUXNOT
    );
  memcontroller_dnl2_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_5_CEMUXNOT
    );
  mac_control_lmacaddr_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_29_FFX_RST,
      O => mac_control_lmacaddr(29)
    );
  mac_control_lmacaddr_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_29_FFX_RST
    );
  memcontroller_dnl2_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_7_CEMUXNOT
    );
  memcontroller_dnl2_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_9_CEMUXNOT
    );
  rx_input_memio_crccomb_Mxor_CO_7_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0118(1),
      ADR1 => rx_input_memio_crccomb_n0118(0),
      ADR2 => rx_input_memio_crccomb_Mxor_CO_7_Xo(1),
      ADR3 => rx_input_memio_crccomb_n0124(0),
      O => rx_input_memio_crcl_7_FROM
    );
  rx_input_memio_n0048_7_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_7_Q,
      O => rx_input_memio_n0048(7)
    );
  rx_input_memio_crcl_7_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_7_FROM,
      O => rx_input_memio_crc_7_Q
    );
  slowclock_rxcrcerrl_LOGIC_ZERO_1666 : X_ZERO
    port map (
      O => slowclock_rxcrcerrl_LOGIC_ZERO
    );
  slowclock_rxcrcerrl_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => slowclock_rxcrcerrl_GROM
    );
  mac_control_lmacaddr_39 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lmacaddr_39_FFX_RST,
      O => mac_control_lmacaddr(39)
    );
  mac_control_lmacaddr_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_39_FFX_RST
    );
  tx_output_addr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(8),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_8_FFX_RST,
      O => addr2ext(8)
    );
  addr2ext_8_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_8_FFX_RST
    );
  tx_output_addr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(10),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_10_FFX_RST,
      O => addr2ext(10)
    );
  addr2ext_10_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_10_FFX_RST
    );
  tx_output_addr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(12),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_12_FFX_RST,
      O => addr2ext(12)
    );
  addr2ext_12_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_12_FFX_RST
    );
  tx_output_addr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(15),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_14_FFY_RST,
      O => addr2ext(15)
    );
  addr2ext_14_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_14_FFY_RST
    );
  rx_input_memio_bcnt_86_1667 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_235,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_86_FFY_RST,
      O => rx_input_memio_bcnt_86
    );
  rx_input_memio_bcnt_86_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_86_FFY_RST
    );
  tx_output_addr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(4),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_4_FFX_RST,
      O => addr2ext(4)
    );
  addr2ext_4_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_4_FFX_RST
    );
  tx_output_addr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(6),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_6_FFX_RST,
      O => addr2ext(6)
    );
  addr2ext_6_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_6_FFX_RST
    );
  tx_output_addr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(9),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_8_FFY_RST,
      O => addr2ext(9)
    );
  addr2ext_8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_8_FFY_RST
    );
  tx_output_addr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(11),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_10_FFY_RST,
      O => addr2ext(11)
    );
  addr2ext_10_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_10_FFY_RST
    );
  tx_output_addr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(13),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_12_FFY_RST,
      O => addr2ext(13)
    );
  addr2ext_12_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_12_FFY_RST
    );
  rx_input_memio_bcnt_95_1668 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_244,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_95_FFX_RST,
      O => rx_input_memio_bcnt_95
    );
  rx_input_memio_bcnt_95_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_95_FFX_RST
    );
  rx_input_memio_bcnt_97_1669 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_246,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_97_FFX_RST,
      O => rx_input_memio_bcnt_97
    );
  rx_input_memio_bcnt_97_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_97_FFX_RST
    );
  rx_input_memio_bcnt_100_1670 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_249,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_99_FFY_RST,
      O => rx_input_memio_bcnt_100
    );
  rx_input_memio_bcnt_99_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_99_FFY_RST
    );
  rx_input_memio_bcnt_101_1671 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_250,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_101_FFX_RST,
      O => rx_input_memio_bcnt_101
    );
  rx_input_memio_bcnt_101_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_101_FFX_RST
    );
  rx_input_memio_bcnt_99_1672 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_248,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_99_FFX_RST,
      O => rx_input_memio_bcnt_99
    );
  rx_input_memio_bcnt_99_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_99_FFX_RST
    );
  mac_control_rxcrcerr_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(1),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(1)
    );
  mac_control_rxcrcerr_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(3),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(3)
    );
  mac_control_rxcrcerr_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(8),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(8)
    );
  mac_control_rxcrcerr_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(10),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(10)
    );
  mac_control_rxcrcerr_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(13),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(13)
    );
  mac_control_rxcrcerr_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(17),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(17)
    );
  mac_control_rxcrcerr_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(12),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(12)
    );
  mac_control_rxcrcerr_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(15),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(15)
    );
  mac_control_rxoferr_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(12),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(12)
    );
  mac_control_rxoferr_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(14),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(14)
    );
  mac_control_rxoferr_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(21),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(21)
    );
  mac_control_rxoferr_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(16),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(16)
    );
  mac_control_rxoferr_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(19),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(19)
    );
  mac_control_rxoferr_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(23),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(23)
    );
  rx_input_memio_BPOUT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_15_54,
      CE => rxbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_15_FFX_RST,
      O => rxbp(15)
    );
  rxbp_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_15_FFX_RST
    );
  rx_output_cs_FFd10_In11_1_1673 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_cs_FFd7,
      ADR2 => rx_output_cs_FFd9,
      ADR3 => VCC,
      O => rx_output_cs_FFd10_In11_1_GROM
    );
  rx_output_cs_FFd10_In11_1_YUSED : X_BUF
    port map (
      I => rx_output_cs_FFd10_In11_1_GROM,
      O => rx_output_cs_FFd10_In11_1
    );
  rx_output_fifo_BU30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1835,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => rx_output_invalid_FFX_RST,
      O => rx_output_invalid
    );
  rx_output_invalid_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_invalid_FFX_RST
    );
  rx_input_memio_crcll_1_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_1_CEMUXNOT
    );
  rx_input_memio_crcll_3_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_3_CEMUXNOT
    );
  rx_input_memio_crcll_5_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_5_CEMUXNOT
    );
  rx_input_memio_crcll_7_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_7_CEMUXNOT
    );
  memcontroller_Q2_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(2),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_3_FFY_RST,
      O => q2(2)
    );
  q2_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_3_FFY_RST
    );
  rx_input_memio_crcll_9_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_9_CEMUXNOT
    );
  memcontroller_Q2_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(1),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_1_FFX_RST,
      O => q2(1)
    );
  q2_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_1_FFX_RST
    );
  tx_output_ltxd_3_1 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => tx_output_outselll(3),
      ADR1 => tx_output_datal(3),
      ADR2 => tx_output_outselll(0),
      ADR3 => tx_output_ncrcbytel(4),
      O => tx_output_ltxd_3_FROM
    );
  tx_output_ltxd_1_1 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => tx_output_outselll(0),
      ADR1 => tx_output_datal(1),
      ADR2 => tx_output_ncrcbytel(6),
      ADR3 => tx_output_outselll(3),
      O => tx_output_ltxd_3_GROM
    );
  tx_output_ltxd_3_XUSED : X_BUF
    port map (
      I => tx_output_ltxd_3_FROM,
      O => tx_output_ltxd(3)
    );
  tx_output_ltxd_3_YUSED : X_BUF
    port map (
      I => tx_output_ltxd_3_GROM,
      O => tx_output_ltxd(1)
    );
  tx_output_ltxd_5_1 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => tx_output_outselll(3),
      ADR1 => tx_output_outselll(0),
      ADR2 => tx_output_ncrcbytel(2),
      ADR3 => tx_output_datal(5),
      O => tx_output_ltxd_5_GROM
    );
  tx_output_ltxd_5_YUSED : X_BUF
    port map (
      I => tx_output_ltxd_5_GROM,
      O => tx_output_ltxd(5)
    );
  tx_output_crc_loigc_Mxor_CO_17_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0104(0),
      ADR1 => tx_output_crc_loigc_n0122(0),
      ADR2 => tx_output_crcl(9),
      ADR3 => tx_output_crc_loigc_n0118(0),
      O => tx_output_crcl_17_FROM
    );
  tx_output_n0034_17_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crc_17_Q,
      O => tx_output_n0034(17)
    );
  tx_output_crcl_17_XUSED : X_BUF
    port map (
      I => tx_output_crcl_17_FROM,
      O => tx_output_crc_17_Q
    );
  rx_input_memio_crccomb_Mxor_CO_12_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_datal(2),
      ADR1 => rx_input_memio_crccomb_Mxor_CO_23_Xo(0),
      ADR2 => rx_input_memio_crcl(29),
      ADR3 => rx_input_memio_crccomb_n0118(1),
      O => rx_input_memio_crcl_12_FROM
    );
  rx_input_memio_n0048_12_1 : X_LUT4
    generic map(
      INIT => X"BBEE"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_2,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crccomb_Mxor_CO_12_Xo(1),
      O => rx_input_memio_n0048(12)
    );
  rx_input_memio_crcl_12_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_12_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_12_Xo(1)
    );
  rx_input_memio_dout_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_21_FFY_RST
    );
  rx_input_memio_dout_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_21_FFY_RST,
      O => rx_input_memio_dout(20)
    );
  rx_input_memio_dout_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_13_FFY_RST
    );
  rx_input_memio_dout_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_13_FFY_RST,
      O => rx_input_memio_dout(12)
    );
  mac_control_PHY_status_MII_Interface_dreg_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_12_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(10),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_12_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(11)
    );
  memcontroller_Q2_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(3),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_3_FFX_RST,
      O => q2(3)
    );
  q2_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_3_FFX_RST
    );
  rx_input_memio_dout_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_23_FFY_RST
    );
  rx_input_memio_dout_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_23_FFY_RST,
      O => rx_input_memio_dout(22)
    );
  rx_input_memio_dout_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_15_FFY_RST
    );
  rx_input_memio_dout_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_15_FFY_RST,
      O => rx_input_memio_dout(14)
    );
  mac_control_PHY_status_MII_Interface_dreg_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_14_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(12),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_14_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(13)
    );
  rx_input_memio_dout_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_17_FFY_RST
    );
  rx_input_memio_dout_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_17_FFY_RST,
      O => rx_input_memio_dout(16)
    );
  mac_control_PHY_status_MII_Interface_dreg_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_15_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(14),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_15_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(15)
    );
  memcontroller_Q2_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(4),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_5_FFY_RST,
      O => q2(4)
    );
  q2_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_5_FFY_RST
    );
  rx_input_memio_dout_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_19_FFY_RST
    );
  rx_input_memio_dout_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_19_FFY_RST,
      O => rx_input_memio_dout(18)
    );
  rx_input_memio_dout_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_29_FFY_RST
    );
  rx_input_memio_dout_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_29_FFY_RST,
      O => rx_input_memio_dout(28)
    );
  mac_control_phydi_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_1_FFY_RST
    );
  mac_control_phydi_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_1_FFY_RST,
      O => mac_control_phydi(0)
    );
  rx_input_memio_bpen_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_bpen_CEMUXNOT
    );
  memcontroller_Q2_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(5),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_5_FFX_RST,
      O => q2(5)
    );
  q2_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_5_FFX_RST
    );
  rx_input_memio_addrchk_n0053_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_rxbcastl,
      ADR1 => rx_input_memio_addrchk_validbcast,
      ADR2 => rx_input_memio_addrchk_rxmcastl,
      ADR3 => rx_input_memio_addrchk_validmcast,
      O => rx_input_memio_destok_FROM
    );
  rx_input_memio_addrchk_n0053_1674 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_rxallfl,
      ADR1 => rx_input_memio_addrchk_rxucastl,
      ADR2 => rx_input_memio_addrchk_validucast,
      ADR3 => rx_input_memio_addrchk_N70965,
      O => rx_input_memio_addrchk_n0053
    );
  rx_input_memio_destok_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_destok_CEMUXNOT
    );
  rx_input_memio_destok_XUSED : X_BUF
    port map (
      I => rx_input_memio_destok_FROM,
      O => rx_input_memio_addrchk_N70965
    );
  mac_control_n0033102_SW0_2_1675 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => mac_control_CHOICE2974,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE2971,
      ADR3 => mac_control_CHOICE2966,
      O => mac_control_n0033102_SW0_2_FROM
    );
  mac_control_n0033102_SW0 : X_LUT4
    generic map(
      INIT => X"0005"
    )
    port map (
      ADR0 => mac_control_CHOICE2978,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE2981,
      ADR3 => mac_control_n0033102_SW0_2,
      O => mac_control_n0033102_SW0_2_GROM
    );
  mac_control_n0033102_SW0_2_XUSED : X_BUF
    port map (
      I => mac_control_n0033102_SW0_2_FROM,
      O => mac_control_n0033102_SW0_2
    );
  mac_control_n0033102_SW0_2_YUSED : X_BUF
    port map (
      I => mac_control_n0033102_SW0_2_GROM,
      O => mac_control_N81729
    );
  rx_output_cs_FFd10_In9 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_output_cs_FFd1,
      ADR1 => rx_output_cs_FFd3,
      ADR2 => rx_output_cs_FFd11,
      ADR3 => rx_output_cs_FFd2,
      O => rx_output_cs_FFd10_FROM
    );
  rx_output_cs_FFd10_In24 : X_LUT4
    generic map(
      INIT => X"0F0E"
    )
    port map (
      ADR0 => rx_output_cs_FFd10_In11_1,
      ADR1 => rx_output_CHOICE1557,
      ADR2 => rx_output_nf,
      ADR3 => rx_output_CHOICE1560,
      O => rx_output_cs_FFd10_In
    );
  rx_output_cs_FFd10_XUSED : X_BUF
    port map (
      I => rx_output_cs_FFd10_FROM,
      O => rx_output_CHOICE1560
    );
  tx_output_crc_loigc_Mxor_CO_18_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(26),
      ADR1 => tx_output_data(5),
      ADR2 => tx_output_data(1),
      ADR3 => tx_output_crcl(30),
      O => tx_output_crcl_18_FROM
    );
  tx_output_n0034_18_1 : X_LUT4
    generic map(
      INIT => X"AFFA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => VCC,
      ADR2 => tx_output_crc_loigc_Mxor_CO_18_Xo_2_1_2,
      ADR3 => tx_output_crc_loigc_Mxor_CO_18_Xo(0),
      O => tx_output_n0034(18)
    );
  tx_output_crcl_18_XUSED : X_BUF
    port map (
      I => tx_output_crcl_18_FROM,
      O => tx_output_crc_loigc_Mxor_CO_18_Xo(0)
    );
  tx_output_crc_loigc_Mxor_CO_26_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_Mxor_CO_26_Xo(1),
      ADR1 => tx_output_crc_loigc_n0124(1),
      ADR2 => tx_output_crc_loigc_n0104(0),
      ADR3 => tx_output_crcl(18),
      O => tx_output_crcl_26_FROM
    );
  tx_output_n0034_26_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16,
      ADR2 => VCC,
      ADR3 => tx_output_crc_26_Q,
      O => tx_output_n0034(26)
    );
  tx_output_crcl_26_XUSED : X_BUF
    port map (
      I => tx_output_crcl_26_FROM,
      O => tx_output_crc_26_Q
    );
  memcontroller_Q3_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(1),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_1_FFX_RST,
      O => q3(1)
    );
  q3_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_1_FFX_RST
    );
  mac_control_Mmux_n0017_Result_8_149_SW0 : X_LUT4
    generic map(
      INIT => X"0013"
    )
    port map (
      ADR0 => mac_control_lmacaddr(8),
      ADR1 => mac_control_CHOICE2394,
      ADR2 => mac_control_n0085,
      ADR3 => mac_control_CHOICE2411,
      O => mac_control_dout_8_FROM
    );
  mac_control_Mmux_n0017_Result_8_149 : X_LUT4
    generic map(
      INIT => X"3074"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_n0060,
      ADR2 => mac_control_dout(7),
      ADR3 => mac_control_N81653,
      O => mac_control_N77375
    );
  mac_control_dout_8_XUSED : X_BUF
    port map (
      I => mac_control_dout_8_FROM,
      O => mac_control_N81653
    );
  rx_input_memio_crccomb_Mxor_CO_13_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(27),
      ADR1 => rx_input_memio_crcl(31),
      ADR2 => rx_input_memio_datal(4),
      ADR3 => rx_input_memio_datal(0),
      O => rx_input_memio_crcl_19_FROM
    );
  rx_input_memio_n0048_19_1 : X_LUT4
    generic map(
      INIT => X"BBEE"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => rx_input_memio_crcl(11),
      ADR2 => VCC,
      ADR3 => rx_input_memio_crccomb_Mxor_CO_13_Xo(2),
      O => rx_input_memio_n0048(19)
    );
  rx_input_memio_crcl_19_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_19_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_13_Xo(2)
    );
  slowclock_rxphyerrl_LOGIC_ZERO_1676 : X_ZERO
    port map (
      O => slowclock_rxphyerrl_LOGIC_ZERO
    );
  slowclock_rxphyerrl_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => slowclock_rxphyerrl_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_13_Xo_5_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_Mxor_n0007_Xo(0),
      ADR1 => rx_input_memio_crccomb_Mxor_CO_13_Xo(2),
      ADR2 => rx_input_memio_crccomb_Mxor_CO_18_Xo(0),
      ADR3 => rx_input_memio_crcl(5),
      O => rx_input_memio_crcl_13_FROM
    );
  rx_input_memio_n0048_13_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_13_Q,
      O => rx_input_memio_n0048(13)
    );
  rx_input_memio_crcl_13_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_13_FROM,
      O => rx_input_memio_crc_13_Q
    );
  mac_control_Mmux_n0017_Result_16_7 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0082,
      ADR1 => mac_control_n0081,
      ADR2 => mac_control_rxfifowerr_cnt(16),
      ADR3 => mac_control_rxphyerr_cnt(16),
      O => mac_control_CHOICE2100_FROM
    );
  mac_control_Mmux_n0017_Result_21_7 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0081,
      ADR1 => mac_control_rxfifowerr_cnt(21),
      ADR2 => mac_control_rxphyerr_cnt(21),
      ADR3 => mac_control_n0082,
      O => mac_control_CHOICE2100_GROM
    );
  mac_control_CHOICE2100_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2100_FROM,
      O => mac_control_CHOICE2100
    );
  mac_control_CHOICE2100_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2100_GROM,
      O => mac_control_CHOICE2148
    );
  mac_control_Mmux_n0017_Result_26_7 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(26),
      ADR1 => mac_control_n0080,
      ADR2 => mac_control_n0081,
      ADR3 => mac_control_rxfifowerr_cnt(26),
      O => mac_control_CHOICE2008_FROM
    );
  mac_control_Mmux_n0017_Result_22_7 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0081,
      ADR1 => mac_control_n0080,
      ADR2 => mac_control_rxfifowerr_cnt(22),
      ADR3 => mac_control_txfifowerr_cnt(22),
      O => mac_control_CHOICE2008_GROM
    );
  mac_control_CHOICE2008_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2008_FROM,
      O => mac_control_CHOICE2008
    );
  mac_control_CHOICE2008_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2008_GROM,
      O => mac_control_CHOICE1962
    );
  mac_control_Mmux_n0017_Result_27_4 : X_LUT4
    generic map(
      INIT => X"3202"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(27),
      ADR1 => mac_control_addr(1),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_rxphyerr_cnt(27),
      O => mac_control_CHOICE1886_FROM
    );
  mac_control_Mmux_n0017_Result_23_4 : X_LUT4
    generic map(
      INIT => X"00AC"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(23),
      ADR1 => mac_control_rxfifowerr_cnt(23),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_addr(1),
      O => mac_control_CHOICE1886_GROM
    );
  mac_control_CHOICE1886_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1886_FROM,
      O => mac_control_CHOICE1886
    );
  mac_control_CHOICE1886_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1886_GROM,
      O => mac_control_CHOICE1858
    );
  mac_control_Mmux_n0017_Result_6_31 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phydi(6),
      ADR1 => mac_control_txf_cnt(6),
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_N52132,
      O => mac_control_CHOICE2315_FROM
    );
  mac_control_Mmux_n0017_Result_0_30 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phydi(0),
      ADR1 => mac_control_txf_cnt(0),
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_N52132,
      O => mac_control_CHOICE2315_GROM
    );
  mac_control_CHOICE2315_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2315_FROM,
      O => mac_control_CHOICE2315
    );
  mac_control_CHOICE2315_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2315_GROM,
      O => mac_control_CHOICE2203
    );
  mac_control_Mmux_n0017_Result_7_65 : X_LUT4
    generic map(
      INIT => X"B080"
    )
    port map (
      ADR0 => mac_control_lmacaddr(39),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_N52143,
      ADR3 => mac_control_lmacaddr(23),
      O => mac_control_CHOICE2840_FROM
    );
  mac_control_Mmux_n0017_Result_23_9 : X_LUT4
    generic map(
      INIT => X"A820"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_rxoferr_cnt(23),
      ADR3 => mac_control_rxcrcerr_cnt(23),
      O => mac_control_CHOICE2840_GROM
    );
  mac_control_CHOICE2840_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2840_FROM,
      O => mac_control_CHOICE2840
    );
  mac_control_CHOICE2840_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2840_GROM,
      O => mac_control_CHOICE1861
    );
  mac_control_Mmux_n0017_Result_18_7 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(18),
      ADR1 => mac_control_n0080,
      ADR2 => mac_control_n0081,
      ADR3 => mac_control_rxfifowerr_cnt(18),
      O => mac_control_CHOICE1916_FROM
    );
  mac_control_Mmux_n0017_Result_24_7 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0082,
      ADR1 => mac_control_rxfifowerr_cnt(24),
      ADR2 => mac_control_n0081,
      ADR3 => mac_control_rxphyerr_cnt(24),
      O => mac_control_CHOICE1916_GROM
    );
  mac_control_CHOICE1916_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1916_FROM,
      O => mac_control_CHOICE1916
    );
  mac_control_CHOICE1916_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1916_GROM,
      O => mac_control_CHOICE2172
    );
  memcontroller_Q2_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(7),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_7_FFX_RST,
      O => q2(7)
    );
  q2_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_7_FFX_RST
    );
  mac_control_Mmux_n0017_Result_0_38 : X_LUT4
    generic map(
      INIT => X"F080"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(0),
      ADR1 => mac_control_N52111,
      ADR2 => mac_control_N52220,
      ADR3 => mac_control_CHOICE2203,
      O => mac_control_CHOICE2205_FROM
    );
  mac_control_Mmux_n0017_Result_0_44 : X_LUT4
    generic map(
      INIT => X"FFE0"
    )
    port map (
      ADR0 => mac_control_CHOICE2197,
      ADR1 => mac_control_CHOICE2194,
      ADR2 => mac_control_N52228,
      ADR3 => mac_control_CHOICE2205,
      O => mac_control_CHOICE2205_GROM
    );
  mac_control_CHOICE2205_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2205_FROM,
      O => mac_control_CHOICE2205
    );
  mac_control_CHOICE2205_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2205_GROM,
      O => mac_control_CHOICE2206
    );
  mac_control_Mmux_n0017_Result_28_7 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0080,
      ADR1 => mac_control_txfifowerr_cnt(28),
      ADR2 => mac_control_n0081,
      ADR3 => mac_control_rxfifowerr_cnt(28),
      O => mac_control_CHOICE2031_FROM
    );
  mac_control_Mmux_n0017_Result_25_7 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0081,
      ADR1 => mac_control_txfifowerr_cnt(25),
      ADR2 => mac_control_rxfifowerr_cnt(25),
      ADR3 => mac_control_n0080,
      O => mac_control_CHOICE2031_GROM
    );
  mac_control_CHOICE2031_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2031_FROM,
      O => mac_control_CHOICE2031
    );
  mac_control_CHOICE2031_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2031_GROM,
      O => mac_control_CHOICE1985
    );
  mac_control_Mmux_n0017_Result_2_69 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_N52118,
      ADR1 => mac_control_txfifowerr_cnt(2),
      ADR2 => mac_control_rxcrcerr_cnt(2),
      ADR3 => mac_control_N52111,
      O => mac_control_CHOICE2284_FROM
    );
  mac_control_Mmux_n0017_Result_0_68 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_N52111,
      ADR1 => mac_control_N52118,
      ADR2 => mac_control_rxcrcerr_cnt(0),
      ADR3 => mac_control_txfifowerr_cnt(0),
      O => mac_control_CHOICE2284_GROM
    );
  mac_control_CHOICE2284_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2284_FROM,
      O => mac_control_CHOICE2284
    );
  mac_control_CHOICE2284_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2284_GROM,
      O => mac_control_CHOICE2210
    );
  mac_control_Mmux_n0017_Result_1_39 : X_LUT4
    generic map(
      INIT => X"EC00"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(1),
      ADR1 => mac_control_CHOICE2239,
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_N52220,
      O => mac_control_CHOICE2241_FROM
    );
  mac_control_Mmux_n0017_Result_1_45 : X_LUT4
    generic map(
      INIT => X"FFA8"
    )
    port map (
      ADR0 => mac_control_N52228,
      ADR1 => mac_control_CHOICE2233,
      ADR2 => mac_control_CHOICE2230,
      ADR3 => mac_control_CHOICE2241,
      O => mac_control_CHOICE2241_GROM
    );
  mac_control_CHOICE2241_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2241_FROM,
      O => mac_control_CHOICE2241
    );
  mac_control_CHOICE2241_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2241_GROM,
      O => mac_control_CHOICE2242
    );
  mac_control_Mmux_n0017_Result_6_86 : X_LUT4
    generic map(
      INIT => X"B800"
    )
    port map (
      ADR0 => mac_control_lmacaddr(38),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_lmacaddr(22),
      ADR3 => mac_control_N52143,
      O => mac_control_CHOICE2328_FROM
    );
  mac_control_Mmux_n0017_Result_1_86 : X_LUT4
    generic map(
      INIT => X"E020"
    )
    port map (
      ADR0 => mac_control_lmacaddr(17),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_N52143,
      ADR3 => mac_control_lmacaddr(33),
      O => mac_control_CHOICE2328_GROM
    );
  mac_control_CHOICE2328_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2328_FROM,
      O => mac_control_CHOICE2328
    );
  mac_control_CHOICE2328_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2328_GROM,
      O => mac_control_CHOICE2252
    );
  mac_control_Mmux_n0017_Result_3_30 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_n0073,
      ADR1 => mac_control_phystat(3),
      ADR2 => mac_control_n0074,
      ADR3 => mac_control_N81741,
      O => mac_control_dout_3_FROM
    );
  mac_control_Mmux_n0017_Result_3_108 : X_LUT4
    generic map(
      INIT => X"3F2F"
    )
    port map (
      ADR0 => mac_control_CHOICE2810,
      ADR1 => mac_control_Mmux_n0017_Result_3_96_1,
      ADR2 => mac_control_Mmux_n0017_Result_3_108_1,
      ADR3 => mac_control_CHOICE2795,
      O => mac_control_N79540
    );
  mac_control_dout_3_XUSED : X_BUF
    port map (
      I => mac_control_dout_3_FROM,
      O => mac_control_CHOICE2795
    );
  mac_control_Mmux_n0017_Result_2_39 : X_LUT4
    generic map(
      INIT => X"E0A0"
    )
    port map (
      ADR0 => mac_control_CHOICE2277,
      ADR1 => mac_control_N52111,
      ADR2 => mac_control_N52220,
      ADR3 => mac_control_rxphyerr_cnt(2),
      O => mac_control_CHOICE2279_FROM
    );
  mac_control_Mmux_n0017_Result_2_45 : X_LUT4
    generic map(
      INIT => X"FFC8"
    )
    port map (
      ADR0 => mac_control_CHOICE2271,
      ADR1 => mac_control_N52228,
      ADR2 => mac_control_CHOICE2268,
      ADR3 => mac_control_CHOICE2279,
      O => mac_control_CHOICE2279_GROM
    );
  mac_control_CHOICE2279_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2279_FROM,
      O => mac_control_CHOICE2279
    );
  mac_control_CHOICE2279_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2279_GROM,
      O => mac_control_CHOICE2280
    );
  mac_control_Mmux_n0017_Result_4_12 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phydi(4),
      ADR1 => mac_control_n0076,
      ADR2 => mac_control_phystat(4),
      ADR3 => mac_control_n0073,
      O => mac_control_CHOICE2603_FROM
    );
  mac_control_Mmux_n0017_Result_4_94_1_1677 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_CHOICE2600,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2603,
      O => mac_control_CHOICE2603_GROM
    );
  mac_control_CHOICE2603_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2603_FROM,
      O => mac_control_CHOICE2603
    );
  mac_control_CHOICE2603_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2603_GROM,
      O => mac_control_Mmux_n0017_Result_4_94_1
    );
  mac_control_Mmux_n0017_Result_3_60 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0085,
      ADR1 => mac_control_lmacaddr(3),
      ADR2 => mac_control_n0084,
      ADR3 => mac_control_rxcrcerr_cnt(3),
      O => mac_control_CHOICE2805_FROM
    );
  mac_control_Mmux_n0017_Result_3_74_SW0 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_CHOICE2808,
      ADR1 => mac_control_n0081,
      ADR2 => mac_control_rxfifowerr_cnt(3),
      ADR3 => mac_control_CHOICE2805,
      O => mac_control_CHOICE2805_GROM
    );
  mac_control_CHOICE2805_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2805_FROM,
      O => mac_control_CHOICE2805
    );
  mac_control_CHOICE2805_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2805_GROM,
      O => mac_control_N81693
    );
  mac_control_Mmux_n0017_Result_4_40 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(4),
      ADR1 => mac_control_n0079,
      ADR2 => mac_control_rxf_cnt(4),
      ADR3 => mac_control_n0080,
      O => mac_control_CHOICE2611_FROM
    );
  mac_control_Mmux_n0017_Result_4_94_SW0_2_1678 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => mac_control_CHOICE2614,
      ADR1 => mac_control_CHOICE2606,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2611,
      O => mac_control_CHOICE2611_GROM
    );
  mac_control_CHOICE2611_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2611_FROM,
      O => mac_control_CHOICE2611
    );
  mac_control_CHOICE2611_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2611_GROM,
      O => mac_control_Mmux_n0017_Result_4_94_SW0_2
    );
  mac_control_Mmux_n0017_Result_3_65 : X_LUT4
    generic map(
      INIT => X"A820"
    )
    port map (
      ADR0 => mac_control_N52143,
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_lmacaddr(19),
      ADR3 => mac_control_lmacaddr(35),
      O => mac_control_CHOICE2808_GROM
    );
  mac_control_CHOICE2808_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2808_GROM,
      O => mac_control_CHOICE2808
    );
  memcontroller_Q3_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(3),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_3_FFX_RST,
      O => q3(3)
    );
  q3_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_3_FFX_RST
    );
  mac_control_Mmux_n0017_Result_4_62 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_lmacaddr(20),
      ADR1 => mac_control_n0086,
      ADR2 => mac_control_n0085,
      ADR3 => mac_control_lmacaddr(4),
      O => mac_control_CHOICE2621_FROM
    );
  mac_control_Mmux_n0017_Result_4_63 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE2618,
      ADR3 => mac_control_CHOICE2621,
      O => mac_control_CHOICE2621_GROM
    );
  mac_control_CHOICE2621_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2621_FROM,
      O => mac_control_CHOICE2621
    );
  mac_control_CHOICE2621_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2621_GROM,
      O => mac_control_CHOICE2622
    );
  mac_control_Mmux_n0017_Result_8_69 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_N52111,
      ADR1 => mac_control_txfifowerr_cnt(8),
      ADR2 => mac_control_N52118,
      ADR3 => mac_control_rxcrcerr_cnt(8),
      O => mac_control_CHOICE2398_FROM
    );
  mac_control_Mmux_n0017_Result_5_31 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_N52118,
      ADR1 => mac_control_phydi(5),
      ADR2 => mac_control_txf_cnt(5),
      ADR3 => mac_control_N52132,
      O => mac_control_CHOICE2398_GROM
    );
  mac_control_CHOICE2398_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2398_FROM,
      O => mac_control_CHOICE2398
    );
  mac_control_CHOICE2398_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2398_GROM,
      O => mac_control_CHOICE2353
    );
  mac_control_Mmux_n0017_Result_4_94 : X_LUT4
    generic map(
      INIT => X"F0E0"
    )
    port map (
      ADR0 => mac_control_Mmux_n0017_Result_4_94_1,
      ADR1 => mac_control_Mmux_n0017_Result_4_94_SW0_2,
      ADR2 => mac_control_N52163,
      ADR3 => mac_control_CHOICE2622,
      O => mac_control_dout_4_FROM
    );
  mac_control_Mmux_n0017_Result_4_105 : X_LUT4
    generic map(
      INIT => X"FF44"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_dout(3),
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2625,
      O => mac_control_N78585
    );
  mac_control_dout_4_XUSED : X_BUF
    port map (
      I => mac_control_dout_4_FROM,
      O => mac_control_CHOICE2625
    );
  mac_control_Mmux_n0017_Result_5_39 : X_LUT4
    generic map(
      INIT => X"C8C0"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(5),
      ADR1 => mac_control_N52220,
      ADR2 => mac_control_CHOICE2353,
      ADR3 => mac_control_N52111,
      O => mac_control_CHOICE2355_FROM
    );
  mac_control_Mmux_n0017_Result_5_45 : X_LUT4
    generic map(
      INIT => X"FFC8"
    )
    port map (
      ADR0 => mac_control_CHOICE2344,
      ADR1 => mac_control_N52228,
      ADR2 => mac_control_CHOICE2347,
      ADR3 => mac_control_CHOICE2355,
      O => mac_control_CHOICE2355_GROM
    );
  mac_control_CHOICE2355_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2355_FROM,
      O => mac_control_CHOICE2355
    );
  mac_control_CHOICE2355_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2355_GROM,
      O => mac_control_CHOICE2356
    );
  mac_control_Mmux_n0017_Result_7_30 : X_LUT4
    generic map(
      INIT => X"FEEE"
    )
    port map (
      ADR0 => mac_control_N81817,
      ADR1 => mac_control_n0074,
      ADR2 => mac_control_phystat(7),
      ADR3 => mac_control_n0073,
      O => mac_control_dout_7_FROM
    );
  mac_control_Mmux_n0017_Result_7_108 : X_LUT4
    generic map(
      INIT => X"EEEA"
    )
    port map (
      ADR0 => mac_control_N82019,
      ADR1 => mac_control_N52163,
      ADR2 => mac_control_CHOICE2842,
      ADR3 => mac_control_CHOICE2827,
      O => mac_control_N79702
    );
  mac_control_dout_7_XUSED : X_BUF
    port map (
      I => mac_control_dout_7_FROM,
      O => mac_control_CHOICE2827
    );
  mac_control_Mmux_n0017_Result_6_39 : X_LUT4
    generic map(
      INIT => X"A8A0"
    )
    port map (
      ADR0 => mac_control_N52220,
      ADR1 => mac_control_N52111,
      ADR2 => mac_control_CHOICE2315,
      ADR3 => mac_control_rxphyerr_cnt(6),
      O => mac_control_CHOICE2317_FROM
    );
  mac_control_Mmux_n0017_Result_6_45 : X_LUT4
    generic map(
      INIT => X"FFA8"
    )
    port map (
      ADR0 => mac_control_N52228,
      ADR1 => mac_control_CHOICE2309,
      ADR2 => mac_control_CHOICE2306,
      ADR3 => mac_control_CHOICE2317,
      O => mac_control_CHOICE2317_GROM
    );
  mac_control_CHOICE2317_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2317_FROM,
      O => mac_control_CHOICE2317
    );
  mac_control_CHOICE2317_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2317_GROM,
      O => mac_control_CHOICE2318
    );
  mac_control_Mmux_n0017_Result_7_60 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_lmacaddr(7),
      ADR1 => mac_control_rxcrcerr_cnt(7),
      ADR2 => mac_control_n0085,
      ADR3 => mac_control_n0084,
      O => mac_control_CHOICE2837_FROM
    );
  mac_control_Mmux_n0017_Result_7_74_SW0 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_n0081,
      ADR1 => mac_control_rxfifowerr_cnt(7),
      ADR2 => mac_control_CHOICE2840,
      ADR3 => mac_control_CHOICE2837,
      O => mac_control_CHOICE2837_GROM
    );
  mac_control_CHOICE2837_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2837_FROM,
      O => mac_control_CHOICE2837
    );
  mac_control_CHOICE2837_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2837_GROM,
      O => mac_control_N81809
    );
  mac_control_Mmux_n0017_Result_7_74 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_n0080,
      ADR1 => mac_control_txfifowerr_cnt(7),
      ADR2 => mac_control_N81809,
      ADR3 => mac_control_CHOICE2833,
      O => mac_control_CHOICE2842_GROM
    );
  mac_control_CHOICE2842_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2842_GROM,
      O => mac_control_CHOICE2842
    );
  mac_control_Mmux_n0017_Result_9_12 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phydi(9),
      ADR1 => mac_control_n0076,
      ADR2 => mac_control_n0073,
      ADR3 => mac_control_phystat(9),
      O => mac_control_CHOICE2634_FROM
    );
  mac_control_Mmux_n0017_Result_9_94_1_1679 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE2631,
      ADR3 => mac_control_CHOICE2634,
      O => mac_control_CHOICE2634_GROM
    );
  mac_control_CHOICE2634_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2634_FROM,
      O => mac_control_CHOICE2634
    );
  mac_control_CHOICE2634_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2634_GROM,
      O => mac_control_Mmux_n0017_Result_9_94_1
    );
  mac_control_Mmux_n0017_Result_8_39 : X_LUT4
    generic map(
      INIT => X"AA80"
    )
    port map (
      ADR0 => mac_control_N52220,
      ADR1 => mac_control_rxphyerr_cnt(8),
      ADR2 => mac_control_N52111,
      ADR3 => mac_control_CHOICE2391,
      O => mac_control_CHOICE2393_FROM
    );
  mac_control_Mmux_n0017_Result_8_45 : X_LUT4
    generic map(
      INIT => X"FFA8"
    )
    port map (
      ADR0 => mac_control_N52228,
      ADR1 => mac_control_CHOICE2382,
      ADR2 => mac_control_CHOICE2385,
      ADR3 => mac_control_CHOICE2393,
      O => mac_control_CHOICE2393_GROM
    );
  mac_control_CHOICE2393_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2393_FROM,
      O => mac_control_CHOICE2393
    );
  mac_control_CHOICE2393_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2393_GROM,
      O => mac_control_CHOICE2394
    );
  mac_control_Mmux_n0017_Result_9_40 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxf_cnt(9),
      ADR1 => mac_control_txfifowerr_cnt(9),
      ADR2 => mac_control_n0079,
      ADR3 => mac_control_n0080,
      O => mac_control_CHOICE2642_FROM
    );
  mac_control_Mmux_n0017_Result_9_94_SW0_2_1680 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => mac_control_CHOICE2645,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE2637,
      ADR3 => mac_control_CHOICE2642,
      O => mac_control_CHOICE2642_GROM
    );
  mac_control_CHOICE2642_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2642_FROM,
      O => mac_control_CHOICE2642
    );
  mac_control_CHOICE2642_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2642_GROM,
      O => mac_control_Mmux_n0017_Result_9_94_SW0_2
    );
  memcontroller_Q2_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(9),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_9_FFX_RST,
      O => q2(9)
    );
  q2_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_9_FFX_RST
    );
  mac_control_Mmux_n0017_Result_9_62 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0085,
      ADR1 => mac_control_lmacaddr(25),
      ADR2 => mac_control_lmacaddr(9),
      ADR3 => mac_control_n0086,
      O => mac_control_CHOICE2652_FROM
    );
  mac_control_Mmux_n0017_Result_9_63 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => mac_control_CHOICE2649,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2652,
      O => mac_control_CHOICE2652_GROM
    );
  mac_control_CHOICE2652_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2652_FROM,
      O => mac_control_CHOICE2652
    );
  mac_control_CHOICE2652_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2652_GROM,
      O => mac_control_CHOICE2653
    );
  mac_control_Mmux_n0017_Result_9_94 : X_LUT4
    generic map(
      INIT => X"AAA8"
    )
    port map (
      ADR0 => mac_control_N52163,
      ADR1 => mac_control_Mmux_n0017_Result_9_94_SW0_2,
      ADR2 => mac_control_Mmux_n0017_Result_9_94_1,
      ADR3 => mac_control_CHOICE2653,
      O => mac_control_dout_9_FROM
    );
  mac_control_Mmux_n0017_Result_9_105 : X_LUT4
    generic map(
      INIT => X"FF22"
    )
    port map (
      ADR0 => mac_control_dout(8),
      ADR1 => mac_control_n0060,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2656,
      O => mac_control_N78742
    );
  mac_control_dout_9_XUSED : X_BUF
    port map (
      I => mac_control_dout_9_FROM,
      O => mac_control_CHOICE2656
    );
  tx_output_crc_loigc_Mxor_CO_27_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0124(0),
      ADR1 => tx_output_crc_loigc_n0118(0),
      ADR2 => tx_output_crc_loigc_Mxor_CO_9_Xo(0),
      ADR3 => tx_output_crcl(19),
      O => tx_output_crcl_27_FROM
    );
  tx_output_n0034_27_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crc_27_Q,
      O => tx_output_n0034(27)
    );
  tx_output_crcl_27_XUSED : X_BUF
    port map (
      I => tx_output_crcl_27_FROM,
      O => tx_output_crc_27_Q
    );
  tx_input_cs_FFd12_In_SW0 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => txfifowerr,
      ADR3 => tx_input_DONE,
      O => tx_input_cs_FFd12_FROM
    );
  tx_input_cs_FFd12_In_1681 : X_LUT4
    generic map(
      INIT => X"FF2A"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => tx_input_den,
      ADR2 => tx_input_newfint,
      ADR3 => tx_input_N69386,
      O => tx_input_cs_FFd12_In
    );
  tx_input_cs_FFd12_XUSED : X_BUF
    port map (
      I => tx_input_cs_FFd12_FROM,
      O => tx_input_N69386
    );
  mac_control_Mmux_n0017_Result_3_30_SW0 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_phyaddr(3),
      ADR1 => mac_control_n0103,
      ADR2 => mac_control_CHOICE2793,
      ADR3 => mac_control_CHOICE2790,
      O => mac_control_N81741_GROM
    );
  mac_control_N81741_YUSED : X_BUF
    port map (
      I => mac_control_N81741_GROM,
      O => mac_control_N81741
    );
  mac_control_Mmux_n0017_Result_18_42_1_1682 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0084,
      ADR2 => mac_control_rxcrcerr_cnt(18),
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_18_42_1_FROM
    );
  mac_control_Mmux_n0017_Result_20_42_1_1683 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => mac_control_n0084,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(20),
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_18_42_1_GROM
    );
  mac_control_Mmux_n0017_Result_18_42_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_18_42_1_FROM,
      O => mac_control_Mmux_n0017_Result_18_42_1
    );
  mac_control_Mmux_n0017_Result_18_42_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_18_42_1_GROM,
      O => mac_control_Mmux_n0017_Result_20_42_1
    );
  rx_input_memio_addrchk_macaddrl_11_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_11_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_21_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(20),
      CE => rx_input_memio_addrchk_macaddrl_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_21_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(20)
    );
  rx_input_memio_addrchk_macaddrl_21_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_21_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_13_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(12),
      CE => rx_input_memio_addrchk_macaddrl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_13_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(12)
    );
  rx_input_memio_addrchk_macaddrl_13_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_13_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_31_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(30),
      CE => rx_input_memio_addrchk_macaddrl_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_31_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(30)
    );
  rx_input_memio_addrchk_macaddrl_31_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_31_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_23_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_23_CEMUXNOT
    );
  memcontroller_Q3_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(5),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_5_FFX_RST,
      O => q3(5)
    );
  q3_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_5_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_15_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(14),
      CE => rx_input_memio_addrchk_macaddrl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_15_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(14)
    );
  rx_input_memio_addrchk_macaddrl_15_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_15_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_41_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_40 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(40),
      CE => rx_input_memio_addrchk_macaddrl_41_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_41_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(40)
    );
  rx_input_memio_addrchk_macaddrl_41_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_41_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_33_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_32 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(32),
      CE => rx_input_memio_addrchk_macaddrl_33_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_33_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(32)
    );
  rx_input_memio_addrchk_macaddrl_33_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_33_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_25_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(24),
      CE => rx_input_memio_addrchk_macaddrl_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_25_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(24)
    );
  rx_input_memio_addrchk_macaddrl_25_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_25_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_17_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(16),
      CE => rx_input_memio_addrchk_macaddrl_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_17_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(16)
    );
  rx_input_memio_addrchk_macaddrl_17_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_17_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_43_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_42 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(42),
      CE => rx_input_memio_addrchk_macaddrl_43_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_43_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(42)
    );
  rx_input_memio_addrchk_macaddrl_43_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_43_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_35_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_35_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_27_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(26),
      CE => rx_input_memio_addrchk_macaddrl_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_27_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(26)
    );
  rx_input_memio_addrchk_macaddrl_27_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_27_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_19_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(18),
      CE => rx_input_memio_addrchk_macaddrl_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_19_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(18)
    );
  rx_input_memio_addrchk_macaddrl_19_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_19_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_45_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_44 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(44),
      CE => rx_input_memio_addrchk_macaddrl_45_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_45_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(44)
    );
  rx_input_memio_addrchk_macaddrl_45_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_45_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_37_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_37_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_36 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(36),
      CE => rx_input_memio_addrchk_macaddrl_37_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_37_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(36)
    );
  rx_input_memio_addrchk_macaddrl_37_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_37_CEMUXNOT
    );
  rx_output_FBBP_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(11),
      CE => rxfbbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_11_FFX_RST,
      O => rxfbbp(11)
    );
  rxfbbp_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_11_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_29_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(28),
      CE => rx_input_memio_addrchk_macaddrl_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_29_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(28)
    );
  rx_input_memio_addrchk_macaddrl_29_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_29_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_47_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_46 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(46),
      CE => rx_input_memio_addrchk_macaddrl_47_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_47_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(46)
    );
  rx_input_memio_addrchk_macaddrl_47_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_47_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_39_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_39_CEMUXNOT
    );
  mac_control_Mmux_n0017_Result_18_77_1_1684 : X_LUT4
    generic map(
      INIT => X"F5F5"
    )
    port map (
      ADR0 => mac_control_dout(17),
      ADR1 => VCC,
      ADR2 => mac_control_n0060,
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_18_77_1_FROM
    );
  mac_control_Mmux_n0017_Result_20_77_1_1685 : X_LUT4
    generic map(
      INIT => X"FF55"
    )
    port map (
      ADR0 => mac_control_dout(19),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_n0060,
      O => mac_control_Mmux_n0017_Result_18_77_1_GROM
    );
  mac_control_Mmux_n0017_Result_18_77_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_18_77_1_FROM,
      O => mac_control_Mmux_n0017_Result_18_77_1
    );
  mac_control_Mmux_n0017_Result_18_77_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_18_77_1_GROM,
      O => mac_control_Mmux_n0017_Result_20_77_1
    );
  mac_control_Mmux_n0017_Result_30_77_1_1686 : X_LUT4
    generic map(
      INIT => X"DDDD"
    )
    port map (
      ADR0 => mac_control_dout(29),
      ADR1 => mac_control_n0060,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_30_77_1_FROM
    );
  mac_control_Mmux_n0017_Result_21_80_1_1687 : X_LUT4
    generic map(
      INIT => X"DDDD"
    )
    port map (
      ADR0 => mac_control_dout(20),
      ADR1 => mac_control_n0060,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_30_77_1_GROM
    );
  mac_control_Mmux_n0017_Result_30_77_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_30_77_1_FROM,
      O => mac_control_Mmux_n0017_Result_30_77_1
    );
  mac_control_Mmux_n0017_Result_30_77_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_30_77_1_GROM,
      O => mac_control_Mmux_n0017_Result_21_80_1
    );
  mac_control_Mmux_n0017_Result_25_42_1_1688 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cnt(25),
      ADR1 => mac_control_n0084,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_25_42_1_FROM
    );
  mac_control_Mmux_n0017_Result_30_42_1_1689 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0084,
      ADR2 => mac_control_rxcrcerr_cnt(30),
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_25_42_1_GROM
    );
  mac_control_Mmux_n0017_Result_25_42_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_25_42_1_FROM,
      O => mac_control_Mmux_n0017_Result_25_42_1
    );
  mac_control_Mmux_n0017_Result_25_42_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_25_42_1_GROM,
      O => mac_control_Mmux_n0017_Result_30_42_1
    );
  mac_control_Mmux_n0017_Result_28_42_1_1690 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cnt(28),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_n0084,
      O => mac_control_Mmux_n0017_Result_28_42_1_FROM
    );
  mac_control_Mmux_n0017_Result_22_42_1_1691 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cnt(22),
      ADR1 => VCC,
      ADR2 => mac_control_n0084,
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_28_42_1_GROM
    );
  mac_control_Mmux_n0017_Result_28_42_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_28_42_1_FROM,
      O => mac_control_Mmux_n0017_Result_28_42_1
    );
  mac_control_Mmux_n0017_Result_28_42_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_28_42_1_GROM,
      O => mac_control_Mmux_n0017_Result_22_42_1
    );
  tx_output_crc_loigc_Mxor_CO_28_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0104(0),
      ADR1 => tx_output_crc_loigc_n0118(0),
      ADR2 => tx_output_crc_loigc_n0118(1),
      ADR3 => tx_output_crcl(20),
      O => tx_output_crcl_28_FROM
    );
  tx_output_n0034_28_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crc_28_Q,
      O => tx_output_n0034(28)
    );
  tx_output_crcl_28_XUSED : X_BUF
    port map (
      I => tx_output_crcl_28_FROM,
      O => tx_output_crc_28_Q
    );
  mac_control_Mmux_n0017_Result_25_77_1_1692 : X_LUT4
    generic map(
      INIT => X"FF55"
    )
    port map (
      ADR0 => mac_control_dout(24),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_n0060,
      O => mac_control_Mmux_n0017_Result_25_77_1_FROM
    );
  mac_control_Mmux_n0017_Result_22_77_1_1693 : X_LUT4
    generic map(
      INIT => X"F0FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_dout(21),
      O => mac_control_Mmux_n0017_Result_25_77_1_GROM
    );
  mac_control_Mmux_n0017_Result_25_77_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_25_77_1_FROM,
      O => mac_control_Mmux_n0017_Result_25_77_1
    );
  mac_control_Mmux_n0017_Result_25_77_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_25_77_1_GROM,
      O => mac_control_Mmux_n0017_Result_22_77_1
    );
  rx_input_memio_crccomb_Mxor_CO_23_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_datal(7),
      ADR1 => rx_input_memio_crcl(25),
      ADR2 => rx_input_memio_crcl(24),
      ADR3 => rx_input_memio_datal(6),
      O => rx_input_memio_crcl_23_FROM
    );
  rx_input_memio_n0048_23_1 : X_LUT4
    generic map(
      INIT => X"AFFA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1_2,
      ADR3 => rx_input_memio_crccomb_Mxor_CO_23_Xo(0),
      O => rx_input_memio_n0048(23)
    );
  rx_input_memio_crcl_23_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_23_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_23_Xo(0)
    );
  rx_input_memio_crccomb_Mxor_CO_15_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_Mxor_CO_13_Xo(2),
      ADR1 => rx_input_memio_crccomb_n0115(0),
      ADR2 => rx_input_memio_crcl(7),
      ADR3 => rx_input_memio_crccomb_n0118(0),
      O => rx_input_memio_crcl_15_FROM
    );
  rx_input_memio_n0048_15_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_15_Q,
      O => rx_input_memio_n0048(15)
    );
  rx_input_memio_crcl_15_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_15_FROM,
      O => rx_input_memio_crc_15_Q
    );
  mac_control_Mmux_n0017_Result_16_80_1_1694 : X_LUT4
    generic map(
      INIT => X"FF0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_dout(15),
      ADR3 => mac_control_n0060,
      O => mac_control_Mmux_n0017_Result_16_80_1_FROM
    );
  mac_control_Mmux_n0017_Result_24_80_1_1695 : X_LUT4
    generic map(
      INIT => X"F5F5"
    )
    port map (
      ADR0 => mac_control_dout(23),
      ADR1 => VCC,
      ADR2 => mac_control_n0060,
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_16_80_1_GROM
    );
  mac_control_Mmux_n0017_Result_16_80_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_16_80_1_FROM,
      O => mac_control_Mmux_n0017_Result_16_80_1
    );
  mac_control_Mmux_n0017_Result_16_80_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_16_80_1_GROM,
      O => mac_control_Mmux_n0017_Result_24_80_1
    );
  rx_input_memio_addrchk_rxallfl_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_rxallfl_CEMUXNOT
    );
  memcontroller_Q3_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(7),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_7_FFX_RST,
      O => q3(7)
    );
  q3_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_7_FFX_RST
    );
  mac_control_Mmux_n0017_Result_28_77_1_1696 : X_LUT4
    generic map(
      INIT => X"F3F3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_dout(27),
      ADR2 => mac_control_n0060,
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_28_77_1_FROM
    );
  mac_control_Mmux_n0017_Result_17_80_1_1697 : X_LUT4
    generic map(
      INIT => X"CFCF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0060,
      ADR2 => mac_control_dout(16),
      ADR3 => VCC,
      O => mac_control_Mmux_n0017_Result_28_77_1_GROM
    );
  mac_control_Mmux_n0017_Result_28_77_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_28_77_1_FROM,
      O => mac_control_Mmux_n0017_Result_28_77_1
    );
  mac_control_Mmux_n0017_Result_28_77_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_28_77_1_GROM,
      O => mac_control_Mmux_n0017_Result_17_80_1
    );
  mac_control_Mmux_n0017_Result_29_42_1_1698 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0084,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(29),
      O => mac_control_Mmux_n0017_Result_29_42_1_FROM
    );
  mac_control_Mmux_n0017_Result_26_42_1_1699 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0084,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(26),
      O => mac_control_Mmux_n0017_Result_29_42_1_GROM
    );
  mac_control_Mmux_n0017_Result_29_42_1_XUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_29_42_1_FROM,
      O => mac_control_Mmux_n0017_Result_29_42_1
    );
  mac_control_Mmux_n0017_Result_29_42_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_29_42_1_GROM,
      O => mac_control_Mmux_n0017_Result_26_42_1
    );
  mac_control_n001220_SW0_1_1700 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => mac_control_bitcnt_109,
      ADR1 => VCC,
      ADR2 => mac_control_sclkdeltall,
      ADR3 => VCC,
      O => mac_control_n001220_SW0_1_GROM
    );
  mac_control_n001220_SW0_1_YUSED : X_BUF
    port map (
      I => mac_control_n001220_SW0_1_GROM,
      O => mac_control_n001220_SW0_1
    );
  mac_control_Mmux_n0017_Result_29_77_1_1701 : X_LUT4
    generic map(
      INIT => X"F0FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_dout(28),
      O => mac_control_Mmux_n0017_Result_29_77_1_GROM
    );
  mac_control_Mmux_n0017_Result_29_77_1_YUSED : X_BUF
    port map (
      I => mac_control_Mmux_n0017_Result_29_77_1_GROM,
      O => mac_control_Mmux_n0017_Result_29_77_1
    );
  tx_output_crc_loigc_Mxor_CO_29_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0104(0),
      ADR1 => tx_output_crc_loigc_n0124(0),
      ADR2 => tx_output_crc_loigc_n0124(1),
      ADR3 => tx_output_crcl(21),
      O => tx_output_crcl_29_FROM
    );
  tx_output_n0034_29_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16,
      ADR2 => VCC,
      ADR3 => tx_output_crc_29_Q,
      O => tx_output_n0034(29)
    );
  tx_output_crcl_29_XUSED : X_BUF
    port map (
      I => tx_output_crcl_29_FROM,
      O => tx_output_crc_29_Q
    );
  rx_input_memio_crcll_11_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_11_CEMUXNOT
    );
  rx_output_FBBP_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(13),
      CE => rxfbbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_13_FFX_RST,
      O => rxfbbp(13)
    );
  rxfbbp_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_13_FFX_RST
    );
  rx_input_memio_crcll_13_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_13_CEMUXNOT
    );
  rx_input_memio_crcll_21_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_21_CEMUXNOT
    );
  rx_input_memio_crcll_15_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_15_CEMUXNOT
    );
  rx_input_memio_crcll_31_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_31_CEMUXNOT
    );
  rx_input_memio_crcll_23_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_23_CEMUXNOT
    );
  rx_input_memio_crcll_17_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_17_CEMUXNOT
    );
  rx_input_memio_crcll_25_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_25_CEMUXNOT
    );
  rx_input_memio_crcll_27_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_27_CEMUXNOT
    );
  rx_input_memio_crcll_19_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_19_CEMUXNOT
    );
  rx_input_memio_crcll_29_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_crcll_29_CEMUXNOT
    );
  rx_input_memio_crccomb_Mxor_CO_24_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0118(1),
      ADR1 => rx_input_memio_crccomb_n0122(0),
      ADR2 => rx_input_memio_crcl(16),
      ADR3 => rx_input_memio_crccomb_n0124(0),
      O => rx_input_memio_crcl_24_FROM
    );
  rx_input_memio_n0048_24_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_24_Q,
      O => rx_input_memio_n0048(24)
    );
  rx_input_memio_crcl_24_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_24_FROM,
      O => rx_input_memio_crc_24_Q
    );
  rx_input_memio_crccomb_Mxor_CO_16_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0115(0),
      ADR1 => rx_input_memio_crcl(8),
      ADR2 => rx_input_memio_crccomb_n0122(1),
      ADR3 => rx_input_memio_crccomb_n0118(0),
      O => rx_input_memio_crcl_16_FROM
    );
  rx_input_memio_n0048_16_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_16_Q,
      O => rx_input_memio_n0048(16)
    );
  rx_input_memio_crcl_16_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_16_FROM,
      O => rx_input_memio_crc_16_Q
    );
  mac_control_Ker521301 : X_LUT4
    generic map(
      INIT => X"1100"
    )
    port map (
      ADR0 => mac_control_addr(2),
      ADR1 => mac_control_addr(4),
      ADR2 => VCC,
      ADR3 => mac_control_addr(3),
      O => mac_control_N52132_FROM
    );
  mac_control_n00251 : X_LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_N52100,
      ADR3 => mac_control_N52132,
      O => mac_control_N52132_GROM
    );
  mac_control_N52132_XUSED : X_BUF
    port map (
      I => mac_control_N52132_FROM,
      O => mac_control_N52132
    );
  mac_control_N52132_YUSED : X_BUF
    port map (
      I => mac_control_N52132_GROM,
      O => mac_control_n0025
    );
  memcontroller_Q3_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(9),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_9_FFX_RST,
      O => q3(9)
    );
  q3_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_9_FFX_RST
    );
  mac_control_Ker521231 : X_LUT4
    generic map(
      INIT => X"0101"
    )
    port map (
      ADR0 => mac_control_addr(3),
      ADR1 => mac_control_addr(4),
      ADR2 => mac_control_addr(2),
      ADR3 => VCC,
      O => mac_control_N52125_FROM
    );
  mac_control_Ker520791 : X_LUT4
    generic map(
      INIT => X"C300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_addr(1),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_N52125,
      O => mac_control_N52125_GROM
    );
  mac_control_N52125_XUSED : X_BUF
    port map (
      I => mac_control_N52125_FROM,
      O => mac_control_N52125
    );
  mac_control_N52125_YUSED : X_BUF
    port map (
      I => mac_control_N52125_GROM,
      O => mac_control_N52081
    );
  mac_control_Ker521161 : X_LUT4
    generic map(
      INIT => X"0404"
    )
    port map (
      ADR0 => mac_control_addr(3),
      ADR1 => mac_control_addr(4),
      ADR2 => mac_control_addr(2),
      ADR3 => VCC,
      O => mac_control_N52118_FROM
    );
  mac_control_Mmux_n0017_Result_1_31 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_N52132,
      ADR1 => mac_control_phydi(1),
      ADR2 => mac_control_txf_cnt(1),
      ADR3 => mac_control_N52118,
      O => mac_control_N52118_GROM
    );
  mac_control_N52118_XUSED : X_BUF
    port map (
      I => mac_control_N52118_FROM,
      O => mac_control_N52118
    );
  mac_control_N52118_YUSED : X_BUF
    port map (
      I => mac_control_N52118_GROM,
      O => mac_control_CHOICE2239
    );
  mac_control_Ker521411 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_addr(3),
      ADR2 => mac_control_addr(2),
      ADR3 => mac_control_addr(4),
      O => mac_control_N52143_FROM
    );
  mac_control_n00311 : X_LUT4
    generic map(
      INIT => X"A000"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => VCC,
      ADR2 => mac_control_N52100,
      ADR3 => mac_control_N52143,
      O => mac_control_N52143_GROM
    );
  mac_control_N52143_XUSED : X_BUF
    port map (
      I => mac_control_N52143_FROM,
      O => mac_control_N52143
    );
  mac_control_N52143_YUSED : X_BUF
    port map (
      I => mac_control_N52143_GROM,
      O => mac_control_n0031
    );
  mac_control_Ker521091 : X_LUT4
    generic map(
      INIT => X"3000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_addr(3),
      ADR2 => mac_control_addr(4),
      ADR3 => mac_control_addr(2),
      O => mac_control_N52111_FROM
    );
  mac_control_Mmux_n0017_Result_2_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_N52118,
      ADR1 => mac_control_rxf_cnt(2),
      ADR2 => mac_control_rxoferr_cnt(2),
      ADR3 => mac_control_N52111,
      O => mac_control_N52111_GROM
    );
  mac_control_N52111_XUSED : X_BUF
    port map (
      I => mac_control_N52111_FROM,
      O => mac_control_N52111
    );
  mac_control_N52111_YUSED : X_BUF
    port map (
      I => mac_control_N52111_GROM,
      O => mac_control_CHOICE2271
    );
  mac_control_Ker522341 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_addr(1),
      O => mac_control_N52236_FROM
    );
  mac_control_n00281 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_N52100,
      ADR1 => mac_control_addr(2),
      ADR2 => mac_control_N52268,
      ADR3 => mac_control_N52236,
      O => mac_control_N52236_GROM
    );
  mac_control_N52236_XUSED : X_BUF
    port map (
      I => mac_control_N52236_FROM,
      O => mac_control_N52236
    );
  mac_control_N52236_YUSED : X_BUF
    port map (
      I => mac_control_N52236_GROM,
      O => mac_control_n0028
    );
  mac_control_Ker522261 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_addr(1),
      O => mac_control_N52228_FROM
    );
  mac_control_n00261 : X_LUT4
    generic map(
      INIT => X"0080"
    )
    port map (
      ADR0 => mac_control_N52228,
      ADR1 => mac_control_N52100,
      ADR2 => mac_control_N52268,
      ADR3 => mac_control_addr(2),
      O => mac_control_N52228_GROM
    );
  mac_control_N52228_XUSED : X_BUF
    port map (
      I => mac_control_N52228_FROM,
      O => mac_control_N52228
    );
  mac_control_N52228_YUSED : X_BUF
    port map (
      I => mac_control_N52228_GROM,
      O => mac_control_n0026
    );
  mac_control_Ker522181 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_addr(0),
      ADR2 => VCC,
      ADR3 => mac_control_addr(1),
      O => mac_control_N52220_FROM
    );
  mac_control_n00781 : X_LUT4
    generic map(
      INIT => X"0400"
    )
    port map (
      ADR0 => mac_control_addr(3),
      ADR1 => mac_control_addr(4),
      ADR2 => mac_control_addr(2),
      ADR3 => mac_control_N52220,
      O => mac_control_N52220_GROM
    );
  mac_control_N52220_XUSED : X_BUF
    port map (
      I => mac_control_N52220_FROM,
      O => mac_control_N52220
    );
  mac_control_N52220_YUSED : X_BUF
    port map (
      I => mac_control_N52220_GROM,
      O => mac_control_n0078
    );
  mac_control_Ker522421 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_addr(1),
      ADR3 => mac_control_addr(0),
      O => mac_control_N52244_FROM
    );
  mac_control_n00271 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => mac_control_addr(2),
      ADR1 => mac_control_N52100,
      ADR2 => mac_control_N52268,
      ADR3 => mac_control_N52244,
      O => mac_control_N52244_GROM
    );
  mac_control_N52244_XUSED : X_BUF
    port map (
      I => mac_control_N52244_FROM,
      O => mac_control_N52244
    );
  mac_control_N52244_YUSED : X_BUF
    port map (
      I => mac_control_N52244_GROM,
      O => mac_control_n0027
    );
  mac_control_Ker522491 : X_LUT4
    generic map(
      INIT => X"0005"
    )
    port map (
      ADR0 => mac_control_bitcnt_108,
      ADR1 => VCC,
      ADR2 => mac_control_bitcnt_107,
      ADR3 => mac_control_bitcnt_109,
      O => mac_control_N52251_FROM
    );
  mac_control_n00111 : X_LUT4
    generic map(
      INIT => X"0020"
    )
    port map (
      ADR0 => mac_control_sclkdelta,
      ADR1 => RESET_IBUF,
      ADR2 => clkslen,
      ADR3 => mac_control_N52251,
      O => mac_control_N52251_GROM
    );
  mac_control_N52251_XUSED : X_BUF
    port map (
      I => mac_control_N52251_FROM,
      O => mac_control_N52251
    );
  mac_control_N52251_YUSED : X_BUF
    port map (
      I => mac_control_N52251_GROM,
      O => mac_control_n0011
    );
  mac_control_Ker520981 : X_LUT4
    generic map(
      INIT => X"0080"
    )
    port map (
      ADR0 => mac_control_newcmd,
      ADR1 => mac_control_addr(7),
      ADR2 => clkslen,
      ADR3 => RESET_IBUF,
      O => mac_control_N52100_GROM
    );
  mac_control_N52100_YUSED : X_BUF
    port map (
      I => mac_control_N52100_GROM,
      O => mac_control_N52100
    );
  mac_control_Ker522661 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_addr(4),
      ADR2 => VCC,
      ADR3 => mac_control_addr(3),
      O => mac_control_N52268_FROM
    );
  mac_control_n00291 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_N52220,
      ADR1 => mac_control_N52100,
      ADR2 => mac_control_addr(2),
      ADR3 => mac_control_N52268,
      O => mac_control_N52268_GROM
    );
  mac_control_N52268_XUSED : X_BUF
    port map (
      I => mac_control_N52268_FROM,
      O => mac_control_N52268
    );
  mac_control_N52268_YUSED : X_BUF
    port map (
      I => mac_control_N52268_GROM,
      O => mac_control_n0029
    );
  rx_output_FBBP_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(15),
      CE => rxfbbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_15_FFX_RST,
      O => rxfbbp(15)
    );
  rxfbbp_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_15_FFX_RST
    );
  mac_control_Ker521961 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => clkslen,
      O => mac_control_N52198_GROM
    );
  mac_control_N52198_YUSED : X_BUF
    port map (
      I => mac_control_N52198_GROM,
      O => mac_control_N52198
    );
  rx_input_memio_cs_FFd3_In_1_1702 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_fifofulll,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_endbyte(2),
      O => rx_input_memio_cs_FFd3_FROM
    );
  rx_input_memio_cs_FFd3_In_1703 : X_LUT4
    generic map(
      INIT => X"F070"
    )
    port map (
      ADR0 => rx_input_memio_crcequal,
      ADR1 => rx_input_memio_destok,
      ADR2 => rx_input_memio_cs_FFd5,
      ADR3 => rx_input_memio_cs_FFd3_In_1,
      O => rx_input_memio_cs_FFd3_In
    );
  rx_input_memio_cs_FFd3_XUSED : X_BUF
    port map (
      I => rx_input_memio_cs_FFd3_FROM,
      O => rx_input_memio_cs_FFd3_In_1
    );
  mac_control_PHY_status_MII_Interface_sout330 : X_LUT4
    generic map(
      INIT => X"88C8"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_CHOICE2562,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR2 => mac_control_PHY_status_MII_Interface_CHOICE2555,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(2),
      O => mac_control_PHY_status_MII_Interface_CHOICE2564_FROM
    );
  mac_control_PHY_status_MII_Interface_sout498 : X_LUT4
    generic map(
      INIT => X"FFFD"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_sout498_2,
      ADR1 => mac_control_PHY_status_MII_Interface_CHOICE2526,
      ADR2 => mac_control_PHY_status_MII_Interface_CHOICE2593,
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE2564,
      O => mac_control_PHY_status_MII_Interface_CHOICE2564_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE2564_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2564_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2564
    );
  mac_control_PHY_status_MII_Interface_CHOICE2564_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2564_GROM,
      O => mac_control_PHY_status_MII_Interface_sout
    );
  mac_control_PHY_status_MII_Interface_sout361 : X_LUT4
    generic map(
      INIT => X"0CAA"
    )
    port map (
      ADR0 => mac_control_PHY_status_miiaddr(3),
      ADR1 => mac_control_PHY_status_din(5),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(4),
      O => mac_control_PHY_status_MII_Interface_CHOICE2574_FROM
    );
  mac_control_PHY_status_MII_Interface_sout365 : X_LUT4
    generic map(
      INIT => X"FFB0"
    )
    port map (
      ADR0 => mac_control_PHY_status_din(1),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE2574,
      O => mac_control_PHY_status_MII_Interface_CHOICE2574_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE2574_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2574_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2574
    );
  mac_control_PHY_status_MII_Interface_CHOICE2574_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2574_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2575
    );
  rx_input_memio_cs_FFd4_In_2_1704 : X_LUT4
    generic map(
      INIT => X"DDFF"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd5,
      ADR1 => rx_input_memio_endbyte(2),
      ADR2 => VCC,
      ADR3 => rx_input_memio_crcequal,
      O => rx_input_memio_cs_FFd4_FROM
    );
  rx_input_memio_cs_FFd4_In_1705 : X_LUT4
    generic map(
      INIT => X"0022"
    )
    port map (
      ADR0 => rx_input_memio_destok,
      ADR1 => rx_input_memio_fifofulll,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd4_In_2,
      O => rx_input_memio_cs_FFd4_In
    );
  rx_input_memio_cs_FFd4_XUSED : X_BUF
    port map (
      I => rx_input_memio_cs_FFd4_FROM,
      O => rx_input_memio_cs_FFd4_In_2
    );
  mac_control_PHY_status_MII_Interface_sout442 : X_LUT4
    generic map(
      INIT => X"5444"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR1 => mac_control_PHY_status_MII_Interface_CHOICE2588,
      ADR2 => mac_control_PHY_status_MII_Interface_CHOICE2575,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(3),
      O => mac_control_PHY_status_MII_Interface_CHOICE2591_FROM
    );
  mac_control_PHY_status_MII_Interface_sout472 : X_LUT4
    generic map(
      INIT => X"CF0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(1),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(5),
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE2591,
      O => mac_control_PHY_status_MII_Interface_CHOICE2591_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE2591_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2591_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2591
    );
  mac_control_PHY_status_MII_Interface_CHOICE2591_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE2591_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2593
    );
  tx_output_bpl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bpl_1_CEMUXNOT
    );
  tx_output_bpl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bpl_3_CEMUXNOT
    );
  tx_output_bpl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bpl_5_CEMUXNOT
    );
  tx_output_bpl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bpl_7_CEMUXNOT
    );
  tx_output_bpl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_bpl_9_CEMUXNOT
    );
  tx_output_addrinc_SW0 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd12,
      ADR3 => tx_output_cs_FFd16,
      O => tx_output_N69282_FROM
    );
  tx_output_addrinc_1706 : X_LUT4
    generic map(
      INIT => X"FEEE"
    )
    port map (
      ADR0 => tx_output_N69282,
      ADR1 => tx_output_cs_FFd7,
      ADR2 => tx_output_n0035,
      ADR3 => tx_output_cs_FFd8,
      O => tx_output_N69282_GROM
    );
  tx_output_N69282_XUSED : X_BUF
    port map (
      I => tx_output_N69282_FROM,
      O => tx_output_N69282
    );
  tx_output_N69282_YUSED : X_BUF
    port map (
      I => tx_output_N69282_GROM,
      O => tx_output_addrinc
    );
  tx_output_bpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(11),
      CE => tx_output_bpl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_11_FFX_RST,
      O => tx_output_bpl(11)
    );
  tx_output_bpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_11_FFX_RST
    );
  tx_output_bpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(13),
      CE => tx_output_bpl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_13_FFX_RST,
      O => tx_output_bpl(13)
    );
  tx_output_bpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_13_FFX_RST
    );
  mac_control_PHY_status_addrl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_addrl_3_FFY_RST
    );
  mac_control_PHY_status_addrl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(2),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_addrl_3_FFY_RST,
      O => mac_control_PHY_status_addrl(2)
    );
  mac_control_PHY_status_addrl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_addrl_4_FFY_RST
    );
  mac_control_PHY_status_addrl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(4),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_addrl_4_FFY_RST,
      O => mac_control_PHY_status_addrl(4)
    );
  tx_input_Ker3448094 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => tx_input_CNT(1),
      ADR1 => tx_input_CNT(0),
      ADR2 => tx_input_CNT(2),
      ADR3 => tx_input_CNT(3),
      O => tx_input_CHOICE1722_FROM
    );
  tx_input_Ker3448012 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_input_CNT(2),
      ADR1 => tx_input_CNT(0),
      ADR2 => tx_input_CNT(3),
      ADR3 => tx_input_CNT(1),
      O => tx_input_CHOICE1722_GROM
    );
  tx_input_CHOICE1722_XUSED : X_BUF
    port map (
      I => tx_input_CHOICE1722_FROM,
      O => tx_input_CHOICE1722
    );
  tx_input_CHOICE1722_YUSED : X_BUF
    port map (
      I => tx_input_CHOICE1722_GROM,
      O => tx_input_CHOICE1695
    );
  tx_input_Ker3448025 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_input_CNT(5),
      ADR1 => tx_input_CNT(6),
      ADR2 => tx_input_CNT(7),
      ADR3 => tx_input_CNT(4),
      O => tx_input_CHOICE1702_GROM
    );
  tx_input_CHOICE1702_YUSED : X_BUF
    port map (
      I => tx_input_CHOICE1702_GROM,
      O => tx_input_CHOICE1702
    );
  tx_output_cs_Out12_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd12,
      ADR1 => tx_output_cs_FFd16,
      ADR2 => tx_output_cs_FFd10,
      ADR3 => tx_output_cs_FFd11,
      O => tx_output_outsell_1_FROM
    );
  tx_output_cs_Out12 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd13,
      ADR1 => tx_output_cs_FFd15,
      ADR2 => tx_output_cs_FFd14,
      ADR3 => tx_output_N70823,
      O => tx_output_outsel_1_Q
    );
  tx_output_outsell_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => tx_output_outsell_1_CEMUXNOT
    );
  tx_output_outsell_1_XUSED : X_BUF
    port map (
      I => tx_output_outsell_1_FROM,
      O => tx_output_N70823
    );
  rx_input_memio_crccomb_Mxor_CO_17_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0104(0),
      ADR1 => rx_input_memio_crcl(9),
      ADR2 => rx_input_memio_crccomb_n0122(0),
      ADR3 => rx_input_memio_crccomb_n0118(0),
      O => rx_input_memio_crcl_17_FROM
    );
  rx_input_memio_n0048_17_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_17_Q,
      O => rx_input_memio_n0048(17)
    );
  rx_input_memio_crcl_17_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_17_FROM,
      O => rx_input_memio_crc_17_Q
    );
  mac_control_PHY_status_n0019_SW0_2_1707 : X_LUT4
    generic map(
      INIT => X"FFCF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_cs_FFd3,
      ADR2 => mac_control_PHY_status_done,
      ADR3 => RESET_IBUF,
      O => mac_control_PHY_status_n0019_SW0_2_FROM
    );
  mac_control_PHY_status_n0019_1708 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_PHY_status_n0019_2,
      ADR1 => mac_control_PHY_status_cs_FFd6,
      ADR2 => mac_control_PHY_status_cs_FFd5,
      ADR3 => mac_control_PHY_status_n0019_SW0_2,
      O => mac_control_PHY_status_n0019_SW0_2_GROM
    );
  mac_control_PHY_status_n0019_SW0_2_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_n0019_SW0_2_FROM,
      O => mac_control_PHY_status_n0019_SW0_2
    );
  mac_control_PHY_status_n0019_SW0_2_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_n0019_SW0_2_GROM,
      O => mac_control_PHY_status_n0019
    );
  tx_input_Ker3448099 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => tx_input_CNT(4),
      ADR1 => tx_input_CNT(5),
      ADR2 => tx_input_CNT(7),
      ADR3 => tx_input_CNT(6),
      O => tx_input_CHOICE1725_FROM
    );
  tx_input_Ker34480137_2_1709 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => tx_input_CHOICE1732,
      ADR1 => tx_input_CHOICE1722,
      ADR2 => tx_input_CHOICE1729,
      ADR3 => tx_input_CHOICE1725,
      O => tx_input_CHOICE1725_GROM
    );
  tx_input_CHOICE1725_XUSED : X_BUF
    port map (
      I => tx_input_CHOICE1725_FROM,
      O => tx_input_CHOICE1725
    );
  tx_input_CHOICE1725_YUSED : X_BUF
    port map (
      I => tx_input_CHOICE1725_GROM,
      O => tx_input_Ker34480137_2
    );
  tx_output_bpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(15),
      CE => tx_output_bpl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_15_FFX_RST,
      O => tx_output_bpl(15)
    );
  tx_output_bpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_15_FFX_RST
    );
  memcontroller_oel_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_oel_CEMUXNOT
    );
  memcontroller_oel_BYMUX : X_INV
    port map (
      I => memcontroller_oe,
      O => memcontroller_oel_BYMUXNOT
    );
  slowclock_clkcnt_Madd_n0000_Mxor_Result_1_Result1 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => slowclock_clkcnt(0),
      ADR1 => VCC,
      ADR2 => slowclock_clkcnt(1),
      ADR3 => VCC,
      O => slowclock_clkcnt_n0000(1)
    );
  slowclock_clkcnt_0_BXMUX : X_INV
    port map (
      I => slowclock_clkcnt(0),
      O => slowclock_clkcnt_0_BXMUXNOT
    );
  slowclock_RXOFERRSR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_rxoferrl,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxoferrsr_FFY_RST,
      O => rxoferrsr
    );
  rxoferrsr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxoferrsr_FFY_RST
    );
  mac_control_PHY_status_cs_Out51 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_cs_FFd6,
      ADR2 => mac_control_PHY_status_cs_FFd8,
      ADR3 => mac_control_PHY_status_cs_FFd3,
      O => mac_control_PHY_status_MII_Interface_cs_FFd6_FROM
    );
  mac_control_PHY_status_MII_Interface_cs_FFd6_In1 : X_LUT4
    generic map(
      INIT => X"F0FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd6,
      ADR2 => mac_control_PHY_status_done,
      ADR3 => mac_control_PHY_status_start,
      O => mac_control_PHY_status_MII_Interface_cs_FFd6_In
    );
  mac_control_PHY_status_MII_Interface_cs_FFd6_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd6_FROM,
      O => mac_control_PHY_status_start
    );
  rx_input_memio_crccomb_Mxor_CO_18_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(30),
      ADR1 => rx_input_memio_crcl(26),
      ADR2 => rx_input_memio_datal(5),
      ADR3 => rx_input_memio_datal(1),
      O => rx_input_memio_crcl_18_FROM
    );
  rx_input_memio_n0048_18_1 : X_LUT4
    generic map(
      INIT => X"BBEE"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1_2,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crccomb_Mxor_CO_18_Xo(0),
      O => rx_input_memio_n0048(18)
    );
  rx_input_memio_crcl_18_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_18_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_18_Xo(0)
    );
  rx_input_memio_crccomb_Mxor_CO_26_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(18),
      ADR1 => rx_input_memio_crccomb_n0104(0),
      ADR2 => rx_input_memio_crccomb_n0124(1),
      ADR3 => rx_input_memio_crccomb_Mxor_CO_26_Xo(1),
      O => rx_input_memio_crcl_26_FROM
    );
  rx_input_memio_n0048_26_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_26_Q,
      O => rx_input_memio_n0048(26)
    );
  rx_input_memio_crcl_26_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_26_FROM,
      O => rx_input_memio_crc_26_Q
    );
  memcontroller_n01161 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => memcontroller_clknum(0),
      O => memcontroller_clknum_0_GROM
    );
  memcontroller_clknum_0_BXMUX : X_INV
    port map (
      I => memcontroller_clknum(0),
      O => memcontroller_clknum_0_BXMUXNOT
    );
  memcontroller_clknum_0_YUSED : X_BUF
    port map (
      I => memcontroller_clknum_0_GROM,
      O => memcontroller_n0116
    );
  slowclock_txfifowerrl_1710 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_txfifowerrl_GROM,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => txfifowerr,
      SRST => slowclock_txfifowerrl_LOGIC_ZERO,
      O => slowclock_txfifowerrl
    );
  slowclock_rxfifowerrl_LOGIC_ZERO_1711 : X_ZERO
    port map (
      O => slowclock_rxfifowerrl_LOGIC_ZERO
    );
  slowclock_rxfifowerrl_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => slowclock_rxfifowerrl_GROM
    );
  txfbbp_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => txfbbp_1_CEMUXNOT
    );
  txfbbp_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => txfbbp_3_CEMUXNOT
    );
  txfbbp_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => txfbbp_5_CEMUXNOT
    );
  txfbbp_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => txfbbp_7_CEMUXNOT
    );
  txfbbp_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => txfbbp_9_CEMUXNOT
    );
  tx_output_outsell_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd9,
      CE => tx_output_outsell_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outsell_2_FFX_RST,
      O => tx_output_outsell(2)
    );
  tx_output_outsell_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outsell_2_FFX_RST
    );
  rx_input_fifo_control_d0_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_3_FFY_RST
    );
  rx_input_fifo_control_d0_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(2),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_3_FFY_RST,
      O => rx_input_fifo_control_d0(2)
    );
  rx_input_fifo_control_d0_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_5_FFY_RST
    );
  rx_input_fifo_control_d0_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(4),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_5_FFY_RST,
      O => rx_input_fifo_control_d0(4)
    );
  rx_input_fifo_control_d1_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_1_FFY_RST
    );
  rx_input_fifo_control_d1_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(0),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_1_FFY_RST,
      O => rx_input_fifo_control_d1(0)
    );
  rx_input_fifo_control_d1_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_3_FFY_RST
    );
  rx_input_fifo_control_d1_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(2),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_3_FFY_RST,
      O => rx_input_fifo_control_d1(2)
    );
  rx_input_fifo_control_d0_9_LOGIC_ZERO_1712 : X_ZERO
    port map (
      O => rx_input_fifo_control_d0_9_LOGIC_ZERO
    );
  rx_input_fifo_control_dinl_9_rt_1713 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_control_dinl(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_control_dinl_9_rt
    );
  rx_input_fifo_control_d1_9_LOGIC_ZERO_1714 : X_ZERO
    port map (
      O => rx_input_fifo_control_d1_9_LOGIC_ZERO
    );
  rx_input_fifo_control_d0_9_rt_1715 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_control_d0(9),
      O => rx_input_fifo_control_d0_9_rt
    );
  rx_input_fifo_control_d2_9_LOGIC_ZERO_1716 : X_ZERO
    port map (
      O => rx_input_fifo_control_d2_9_LOGIC_ZERO
    );
  rx_input_fifo_control_d1_9_rt_1717 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_control_d1(9),
      O => rx_input_fifo_control_d1_9_rt
    );
  rx_input_memio_endbyte_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_endbyte_1_FFX_RST,
      O => rx_input_memio_endbyte(1)
    );
  rx_input_memio_endbyte_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_endbyte_1_FFX_RST
    );
  rx_input_fifo_control_d3_9_LOGIC_ZERO_1718 : X_ZERO
    port map (
      O => rx_input_fifo_control_d3_9_LOGIC_ZERO
    );
  rx_input_fifo_control_d2_9_rt_1719 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_control_d2(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_control_d2_9_rt
    );
  rx_input_memio_crccomb_Mxor_CO_27_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0124(0),
      ADR1 => rx_input_memio_crcl(19),
      ADR2 => rx_input_memio_crccomb_n0118(0),
      ADR3 => rx_input_memio_crccomb_Mxor_CO_9_Xo(0),
      O => rx_input_memio_crcl_27_FROM
    );
  rx_input_memio_n0048_27_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_27_Q,
      O => rx_input_memio_n0048(27)
    );
  rx_input_memio_crcl_27_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_27_FROM,
      O => rx_input_memio_crc_27_Q
    );
  mac_control_PHY_status_miirw1 : X_LUT4
    generic map(
      INIT => X"0008"
    )
    port map (
      ADR0 => mac_control_PHY_status_rwl,
      ADR1 => mac_control_PHY_status_N41765,
      ADR2 => mac_control_PHY_status_cs_FFd6,
      ADR3 => mac_control_PHY_status_cs_FFd5,
      O => mac_control_PHY_status_miirw_FROM
    );
  mac_control_PHY_status_MII_Interface_sout273_SW2 : X_LUT4
    generic map(
      INIT => X"3120"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR2 => mac_control_PHY_status_din(12),
      ADR3 => mac_control_PHY_status_miirw,
      O => mac_control_PHY_status_miirw_GROM
    );
  mac_control_PHY_status_miirw_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miirw_FROM,
      O => mac_control_PHY_status_miirw
    );
  mac_control_PHY_status_miirw_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miirw_GROM,
      O => mac_control_PHY_status_MII_Interface_N82069
    );
  rx_input_fifo_control_cell_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_cell_CEMUXNOT
    );
  rx_input_memio_crccomb_Mxor_CO_28_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(20),
      ADR1 => rx_input_memio_crccomb_n0104(0),
      ADR2 => rx_input_memio_crccomb_n0118(1),
      ADR3 => rx_input_memio_crccomb_n0118(0),
      O => rx_input_memio_crcl_28_FROM
    );
  rx_input_memio_n0048_28_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_28_Q,
      O => rx_input_memio_n0048(28)
    );
  rx_input_memio_crcl_28_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_28_FROM,
      O => rx_input_memio_crc_28_Q
    );
  mac_control_PHY_status_Ker417711 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_cs_FFd5,
      ADR2 => mac_control_PHY_status_cs_FFd6,
      ADR3 => VCC,
      O => mac_control_PHY_status_N41773_FROM
    );
  mac_control_PHY_status_n00201 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => mac_control_PHY_status_done,
      ADR1 => RESET_IBUF,
      ADR2 => clkslen,
      ADR3 => mac_control_PHY_status_N41773,
      O => mac_control_PHY_status_N41773_GROM
    );
  mac_control_PHY_status_N41773_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_N41773_FROM,
      O => mac_control_PHY_status_N41773
    );
  mac_control_PHY_status_N41773_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_N41773_GROM,
      O => mac_control_PHY_status_n0020
    );
  mac_control_PHY_status_Ker417631 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd3,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_cs_FFd2,
      ADR3 => mac_control_PHY_status_cs_FFd4,
      O => mac_control_PHY_status_N41765_FROM
    );
  mac_control_PHY_status_n00211 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => mac_control_PHY_status_done,
      ADR1 => RESET_IBUF,
      ADR2 => clkslen,
      ADR3 => mac_control_PHY_status_N41765,
      O => mac_control_PHY_status_N41765_GROM
    );
  mac_control_PHY_status_N41765_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_N41765_FROM,
      O => mac_control_PHY_status_N41765
    );
  mac_control_PHY_status_N41765_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_N41765_GROM,
      O => mac_control_PHY_status_n0021
    );
  rx_input_memio_crccomb_Mxor_CO_14_Xo_3_1_SW0 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(30),
      ADR1 => rx_input_memio_crccomb_Mxor_CO_13_Xo(2),
      ADR2 => rx_input_memio_crcl(6),
      ADR3 => rx_input_memio_datal(1),
      O => rx_input_memio_crcl_14_FROM
    );
  rx_input_memio_n0048_14_1 : X_LUT4
    generic map(
      INIT => X"F3FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crccomb_Mxor_CO_14_Xo_3_1_2,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crccomb_N82101,
      O => rx_input_memio_n0048(14)
    );
  rx_input_memio_crcl_14_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_14_FROM,
      O => rx_input_memio_crccomb_N82101
    );
  mac_control_PHY_status_miiaddr_3_1 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_PHY_status_N41765,
      ADR1 => mac_control_PHY_status_addrl(3),
      ADR2 => mac_control_PHY_status_cs_FFd6,
      ADR3 => mac_control_PHY_status_cs_FFd5,
      O => mac_control_PHY_status_miiaddr_3_FROM
    );
  mac_control_PHY_status_miiaddr_0_1 : X_LUT4
    generic map(
      INIT => X"FFEF"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd5,
      ADR1 => mac_control_PHY_status_addrl(0),
      ADR2 => mac_control_PHY_status_N41765,
      ADR3 => mac_control_PHY_status_cs_FFd6,
      O => mac_control_PHY_status_miiaddr_3_GROM
    );
  mac_control_PHY_status_miiaddr_3_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_3_FROM,
      O => mac_control_PHY_status_miiaddr(3)
    );
  mac_control_PHY_status_miiaddr_3_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_3_GROM,
      O => mac_control_PHY_status_miiaddr(0)
    );
  mac_control_PHY_status_miiaddr_1_1 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_PHY_status_addrl(1),
      ADR1 => mac_control_PHY_status_N41765,
      ADR2 => mac_control_PHY_status_cs_FFd6,
      ADR3 => mac_control_PHY_status_cs_FFd5,
      O => mac_control_PHY_status_miiaddr_1_GROM
    );
  mac_control_PHY_status_miiaddr_1_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_1_GROM,
      O => mac_control_PHY_status_miiaddr(1)
    );
  mac_control_PHY_status_miiaddr_2_1 : X_LUT4
    generic map(
      INIT => X"FEEE"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd5,
      ADR1 => mac_control_PHY_status_cs_FFd6,
      ADR2 => mac_control_PHY_status_N41765,
      ADR3 => mac_control_PHY_status_addrl(2),
      O => mac_control_PHY_status_miiaddr_2_FROM
    );
  mac_control_PHY_status_MII_Interface_sout178 : X_LUT4
    generic map(
      INIT => X"8A80"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_din(4),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR3 => mac_control_PHY_status_miiaddr(2),
      O => mac_control_PHY_status_miiaddr_2_GROM
    );
  mac_control_PHY_status_miiaddr_2_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_2_FROM,
      O => mac_control_PHY_status_miiaddr(2)
    );
  mac_control_PHY_status_miiaddr_2_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_2_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2532
    );
  mac_control_PHY_status_miiaddr_4_1 : X_LUT4
    generic map(
      INIT => X"1011"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd6,
      ADR1 => mac_control_PHY_status_cs_FFd5,
      ADR2 => mac_control_PHY_status_addrl(4),
      ADR3 => mac_control_PHY_status_N41765,
      O => mac_control_PHY_status_miiaddr_4_FROM
    );
  mac_control_PHY_status_MII_Interface_sout222 : X_LUT4
    generic map(
      INIT => X"D580"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR1 => mac_control_PHY_status_din(6),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR3 => mac_control_PHY_status_miiaddr(4),
      O => mac_control_PHY_status_miiaddr_4_GROM
    );
  mac_control_PHY_status_miiaddr_4_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_4_FROM,
      O => mac_control_PHY_status_miiaddr(4)
    );
  mac_control_PHY_status_miiaddr_4_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_4_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE2546
    );
  tx_fifocheck_n000212 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(1),
      ADR1 => tx_fifocheck_diff(3),
      ADR2 => tx_fifocheck_diff(2),
      ADR3 => tx_fifocheck_diff(0),
      O => tx_fifocheck_CHOICE1742_GROM
    );
  tx_fifocheck_CHOICE1742_YUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1742_GROM,
      O => tx_fifocheck_CHOICE1742
    );
  rx_input_memio_crccomb_Mxor_CO_29_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0104(0),
      ADR1 => rx_input_memio_crcl(21),
      ADR2 => rx_input_memio_crccomb_n0124(0),
      ADR3 => rx_input_memio_crccomb_n0124(1),
      O => rx_input_memio_crcl_29_FROM
    );
  rx_input_memio_n0048_29_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_29_Q,
      O => rx_input_memio_n0048(29)
    );
  rx_input_memio_crcl_29_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_29_FROM,
      O => rx_input_memio_crc_29_Q
    );
  tx_fifocheck_n000225 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(6),
      ADR1 => tx_fifocheck_diff(7),
      ADR2 => tx_fifocheck_diff(5),
      ADR3 => tx_fifocheck_diff(4),
      O => tx_fifocheck_CHOICE1749_GROM
    );
  tx_fifocheck_CHOICE1749_YUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1749_GROM,
      O => tx_fifocheck_CHOICE1749
    );
  tx_fifocheck_n000262 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(12),
      ADR1 => tx_fifocheck_diff(13),
      ADR2 => tx_fifocheck_diff(14),
      ADR3 => tx_fifocheck_diff(15),
      O => tx_fifocheck_CHOICE1764_GROM
    );
  tx_fifocheck_CHOICE1764_YUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1764_GROM,
      O => tx_fifocheck_CHOICE1764
    );
  tx_fifocheck_n000263 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_fifocheck_CHOICE1757,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_CHOICE1764,
      O => tx_fifocheck_CHOICE1765_FROM
    );
  tx_fifocheck_n000292 : X_LUT4
    generic map(
      INIT => X"ECCC"
    )
    port map (
      ADR0 => tx_fifocheck_CHOICE1749,
      ADR1 => tx_fifocheck_n0003,
      ADR2 => tx_fifocheck_CHOICE1742,
      ADR3 => tx_fifocheck_CHOICE1765,
      O => tx_fifocheck_CHOICE1765_GROM
    );
  tx_fifocheck_CHOICE1765_XUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1765_FROM,
      O => tx_fifocheck_CHOICE1765
    );
  tx_fifocheck_CHOICE1765_YUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1765_GROM,
      O => tx_fifocheck_N73964
    );
  tx_fifocheck_n000249 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(11),
      ADR1 => tx_fifocheck_diff(8),
      ADR2 => tx_fifocheck_diff(10),
      ADR3 => tx_fifocheck_diff(9),
      O => tx_fifocheck_CHOICE1757_GROM
    );
  tx_fifocheck_CHOICE1757_YUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1757_GROM,
      O => tx_fifocheck_CHOICE1757
    );
  rx_input_fifo_control_celll_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_celll_CEMUXNOT
    );
  mac_control_addr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(0),
      CE => mac_control_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_addr_1_FFX_RST,
      O => mac_control_addr(1)
    );
  mac_control_addr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_1_FFX_RST
    );
  rx_input_memio_addrchk_validmcast_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_validmcast_CEMUXNOT
    );
  rx_input_memio_cs_Out910 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd6,
      ADR1 => rx_input_memio_cs_FFd8,
      ADR2 => rx_input_memio_cs_FFd13,
      ADR3 => rx_input_memio_cs_FFd7,
      O => rx_input_memio_CHOICE1570_GROM
    );
  rx_input_memio_CHOICE1570_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1570_GROM,
      O => rx_input_memio_CHOICE1570
    );
  mac_control_addr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(2),
      CE => mac_control_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_addr_3_FFX_RST,
      O => mac_control_addr(3)
    );
  mac_control_addr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_3_FFX_RST
    );
  rx_input_memio_cs_Out8_2_1720 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd10,
      ADR2 => rx_input_memio_cs_FFd15,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_fifo_rd_en_FROM
    );
  rx_input_memio_cs_Out8 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd14,
      ADR2 => rx_input_memio_cs_FFd12,
      ADR3 => rx_input_memio_cs_Out8_2,
      O => rx_input_fifo_rd_en_GROM
    );
  rx_input_fifo_rd_en_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_rd_en_CEMUXNOT
    );
  rx_input_fifo_rd_en_XUSED : X_BUF
    port map (
      I => rx_input_fifo_rd_en_FROM,
      O => rx_input_memio_cs_Out8_2
    );
  rx_input_fifo_rd_en_YUSED : X_BUF
    port map (
      I => rx_input_fifo_rd_en_GROM,
      O => rx_input_ce
    );
  rxfifofull_LOGIC_ONE_1721 : X_ONE
    port map (
      O => rxfifofull_LOGIC_ONE
    );
  rx_input_memio_addrchk_rxbcastl_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_rxbcastl_CEMUXNOT
    );
  mac_control_addr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(4),
      CE => mac_control_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_addr_5_FFX_RST,
      O => mac_control_addr(5)
    );
  mac_control_addr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_5_FFX_RST
    );
  rx_output_n0046_10_SW0 : X_LUT4
    generic map(
      INIT => X"11DD"
    )
    port map (
      ADR0 => rx_output_len(10),
      ADR1 => rx_output_len(1),
      ADR2 => VCC,
      ADR3 => rx_output_n0070(10),
      O => rx_output_lenr_10_FROM
    );
  rx_output_n0046_10_Q : X_LUT4
    generic map(
      INIT => X"A0F5"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => VCC,
      ADR2 => rx_output_n0060(10),
      ADR3 => rx_output_N70216,
      O => rx_output_n0046(10)
    );
  rx_output_lenr_10_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_10_CEMUXNOT
    );
  rx_output_lenr_10_XUSED : X_BUF
    port map (
      I => rx_output_lenr_10_FROM,
      O => rx_output_N70216
    );
  rx_output_n0046_11_SW0 : X_LUT4
    generic map(
      INIT => X"5533"
    )
    port map (
      ADR0 => rx_output_n0070(11),
      ADR1 => rx_output_len(11),
      ADR2 => VCC,
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_11_FROM
    );
  rx_output_n0046_11_Q : X_LUT4
    generic map(
      INIT => X"88BB"
    )
    port map (
      ADR0 => rx_output_n0060(11),
      ADR1 => rx_output_len(0),
      ADR2 => VCC,
      ADR3 => rx_output_N70268,
      O => rx_output_n0046(11)
    );
  rx_output_lenr_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_11_CEMUXNOT
    );
  rx_output_lenr_11_XUSED : X_BUF
    port map (
      I => rx_output_lenr_11_FROM,
      O => rx_output_N70268
    );
  rx_output_n0046_12_SW0 : X_LUT4
    generic map(
      INIT => X"05F5"
    )
    port map (
      ADR0 => rx_output_len(12),
      ADR1 => VCC,
      ADR2 => rx_output_len(1),
      ADR3 => rx_output_n0070(12),
      O => rx_output_lenr_12_FROM
    );
  rx_output_n0046_12_Q : X_LUT4
    generic map(
      INIT => X"A0F5"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => VCC,
      ADR2 => rx_output_n0060(12),
      ADR3 => rx_output_N70320,
      O => rx_output_n0046(12)
    );
  rx_output_lenr_12_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_12_CEMUXNOT
    );
  rx_output_lenr_12_XUSED : X_BUF
    port map (
      I => rx_output_lenr_12_FROM,
      O => rx_output_N70320
    );
  rx_output_n0046_13_SW0 : X_LUT4
    generic map(
      INIT => X"5533"
    )
    port map (
      ADR0 => rx_output_n0070(13),
      ADR1 => rx_output_len(13),
      ADR2 => VCC,
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_13_FROM
    );
  rx_output_n0046_13_Q : X_LUT4
    generic map(
      INIT => X"88DD"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => rx_output_n0060(13),
      ADR2 => VCC,
      ADR3 => rx_output_N69748,
      O => rx_output_n0046(13)
    );
  rx_output_lenr_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_13_CEMUXNOT
    );
  rx_output_lenr_13_XUSED : X_BUF
    port map (
      I => rx_output_lenr_13_FROM,
      O => rx_output_N69748
    );
  mac_control_n0033102 : X_LUT4
    generic map(
      INIT => X"0F0D"
    )
    port map (
      ADR0 => mac_control_N81729,
      ADR1 => mac_control_CHOICE2963,
      ADR2 => mac_control_phyrstcnt_141,
      ADR3 => mac_control_CHOICE2960,
      O => mac_control_CHOICE2986_FROM
    );
  mac_control_n0033124 : X_LUT4
    generic map(
      INIT => X"3020"
    )
    port map (
      ADR0 => mac_control_N52153,
      ADR1 => RESET_IBUF,
      ADR2 => clkslen,
      ADR3 => mac_control_CHOICE2986,
      O => mac_control_CHOICE2986_GROM
    );
  mac_control_CHOICE2986_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2986_FROM,
      O => mac_control_CHOICE2986
    );
  mac_control_CHOICE2986_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2986_GROM,
      O => mac_control_N80441
    );
  rx_output_n0046_14_SW0 : X_LUT4
    generic map(
      INIT => X"0F55"
    )
    port map (
      ADR0 => rx_output_len(14),
      ADR1 => VCC,
      ADR2 => rx_output_n0070(14),
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_14_FROM
    );
  rx_output_n0046_14_Q : X_LUT4
    generic map(
      INIT => X"A0F5"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => VCC,
      ADR2 => rx_output_n0060(14),
      ADR3 => rx_output_N70372,
      O => rx_output_n0046(14)
    );
  rx_output_lenr_14_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_14_CEMUXNOT
    );
  rx_output_lenr_14_XUSED : X_BUF
    port map (
      I => rx_output_lenr_14_FROM,
      O => rx_output_N70372
    );
  rx_output_n0046_15_SW0 : X_LUT4
    generic map(
      INIT => X"05F5"
    )
    port map (
      ADR0 => rx_output_len(15),
      ADR1 => VCC,
      ADR2 => rx_output_len(1),
      ADR3 => rx_output_n0070(15),
      O => rx_output_lenr_15_FROM
    );
  rx_output_n0046_15_Q : X_LUT4
    generic map(
      INIT => X"88DD"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => rx_output_n0060(15),
      ADR2 => VCC,
      ADR3 => rx_output_N69696,
      O => rx_output_n0046(15)
    );
  rx_output_lenr_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_15_CEMUXNOT
    );
  rx_output_lenr_15_XUSED : X_BUF
    port map (
      I => rx_output_lenr_15_FROM,
      O => rx_output_N69696
    );
  tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_SW0 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(6),
      ADR1 => tx_output_crc_loigc_n0104(0),
      ADR2 => tx_output_data(3),
      ADR3 => tx_output_crc_loigc_Mxor_CO_13_Xo(2),
      O => tx_output_crcl_14_FROM
    );
  tx_output_n0034_14_1 : X_LUT4
    generic map(
      INIT => X"BBEE"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_2,
      ADR2 => VCC,
      ADR3 => tx_output_crc_loigc_N81880,
      O => tx_output_n0034(14)
    );
  tx_output_crcl_14_XUSED : X_BUF
    port map (
      I => tx_output_crcl_14_FROM,
      O => tx_output_crc_loigc_N81880
    );
  mac_control_addr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(6),
      CE => mac_control_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_addr_7_FFX_RST,
      O => mac_control_addr(7)
    );
  mac_control_addr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_7_FFX_RST
    );
  rx_input_memio_addrchk_rxmcastl_CEMUX : X_INV
    port map (
      I => rx_input_RESET_1,
      O => rx_input_memio_addrchk_rxmcastl_CEMUXNOT
    );
  rx_input_fifo_control_dinl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_dinl_1_CEMUXNOT
    );
  rx_input_fifo_control_dinl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_dinl_3_CEMUXNOT
    );
  rx_input_fifo_control_dinl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_dinl_5_CEMUXNOT
    );
  rx_input_fifo_control_dinl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_dinl_7_CEMUXNOT
    );
  tx_input_cs_FFd10_1722 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd10_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd10_FFY_RST,
      O => tx_input_cs_FFd10
    );
  tx_input_cs_FFd10_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd10_FFY_RST
    );
  mac_control_din_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_11_FFX_RST,
      O => mac_control_din(11)
    );
  mac_control_din_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_11_FFX_RST
    );
  mac_control_din_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_13_FFY_RST,
      O => mac_control_din(12)
    );
  mac_control_din_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_13_FFY_RST
    );
  mac_control_din_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_13_FFX_RST,
      O => mac_control_din(13)
    );
  mac_control_din_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_13_FFX_RST
    );
  mac_control_din_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(19),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_21_FFY_RST,
      O => mac_control_din(20)
    );
  mac_control_din_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_21_FFY_RST
    );
  mac_control_din_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(20),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_21_FFX_RST,
      O => mac_control_din(21)
    );
  mac_control_din_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_21_FFX_RST
    );
  mac_control_din_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_15_FFX_RST,
      O => mac_control_din(15)
    );
  mac_control_din_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_15_FFX_RST
    );
  mac_control_din_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(21),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_23_FFY_RST,
      O => mac_control_din(22)
    );
  mac_control_din_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_23_FFY_RST
    );
  mac_control_din_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(22),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_23_FFX_RST,
      O => mac_control_din(23)
    );
  mac_control_din_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_23_FFX_RST
    );
  mac_control_din_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(30),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_31_FFX_RST,
      O => mac_control_din(31)
    );
  mac_control_din_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_31_FFX_RST
    );
  mac_control_din_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(23),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_25_FFY_RST,
      O => mac_control_din(24)
    );
  mac_control_din_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_25_FFY_RST
    );
  mac_control_din_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(16),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_17_FFX_RST,
      O => mac_control_din(17)
    );
  mac_control_din_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_17_FFX_RST
    );
  rx_output_FBBP_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(7),
      CE => rxfbbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_7_FFX_RST,
      O => rxfbbp(7)
    );
  rxfbbp_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_7_FFX_RST
    );
  rx_output_FBBP_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(9),
      CE => rxfbbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_9_FFX_RST,
      O => rxfbbp(9)
    );
  rxfbbp_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_9_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(0),
      CE => rx_input_memio_addrchk_macaddrl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_1_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(0)
    );
  rx_input_memio_addrchk_macaddrl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_1_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(1),
      CE => rx_input_memio_addrchk_macaddrl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_1_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(1)
    );
  rx_input_memio_addrchk_macaddrl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_1_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(3),
      CE => rx_input_memio_addrchk_macaddrl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_3_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(3)
    );
  rx_input_memio_addrchk_macaddrl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_3_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(5),
      CE => rx_input_memio_addrchk_macaddrl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_5_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(5)
    );
  rx_input_memio_addrchk_macaddrl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_5_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(7),
      CE => rx_input_memio_addrchk_macaddrl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_7_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(7)
    );
  rx_input_memio_addrchk_macaddrl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_7_FFX_RST
    );
  rx_input_memio_crcl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(4),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_4_FFY_RST,
      O => rx_input_memio_crcl(4)
    );
  rx_input_memio_crcl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_4_FFY_RST
    );
  tx_output_ncrcbytel_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(4),
      CE => tx_output_ncrcbytel_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_4_FFY_RST,
      O => tx_output_ncrcbytel(4)
    );
  tx_output_ncrcbytel_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_4_FFY_RST
    );
  tx_output_crcl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(25),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_25_FFY_RST,
      O => tx_output_crcl(25)
    );
  tx_output_crcl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_25_FFY_RST
    );
  tx_output_ncrcbytel_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(5),
      CE => tx_output_ncrcbytel_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_5_FFY_RST,
      O => tx_output_ncrcbytel(5)
    );
  tx_output_ncrcbytel_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_5_FFY_RST
    );
  tx_output_ncrcbytel_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(6),
      CE => tx_output_ncrcbytel_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_6_FFY_RST,
      O => tx_output_ncrcbytel(6)
    );
  tx_output_ncrcbytel_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_6_FFY_RST
    );
  rx_input_memio_addrchk_validbcast_1723 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_n0051,
      CE => rx_input_memio_addrchk_validbcast_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_validbcast_FFY_RST,
      O => rx_input_memio_addrchk_validbcast
    );
  rx_input_memio_addrchk_validbcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_validbcast_FFY_RST
    );
  tx_output_ncrcbytel_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(7),
      CE => tx_output_ncrcbytel_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_7_FFY_RST,
      O => tx_output_ncrcbytel(7)
    );
  tx_output_ncrcbytel_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_7_FFY_RST
    );
  rx_output_cs_FFd12_1724 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd13,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd12_FFX_RST,
      O => rx_output_cs_FFd12
    );
  rx_output_cs_FFd12_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd12_FFX_RST
    );
  rx_output_cs_FFd14_1725 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd15,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd14_FFX_RST,
      O => rx_output_cs_FFd14
    );
  rx_output_cs_FFd14_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd14_FFX_RST
    );
  rx_output_ceinl_1726 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cein,
      CE => rx_output_ceinl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_ceinl_FFX_RST,
      O => rx_output_ceinl
    );
  rx_output_ceinl_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_ceinl_FFX_RST
    );
  rx_output_cs_FFd16_1727 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd17,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd16_FFX_RST,
      O => rx_output_cs_FFd16
    );
  rx_output_cs_FFd16_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd16_FFX_RST
    );
  mac_control_rxf_cross_1728 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfsr,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_rxf_cross_FFY_RST,
      O => mac_control_rxf_cross
    );
  mac_control_rxf_cross_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cross_FFY_RST
    );
  tx_input_cs_FFd6_1729 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd6_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd6_FFX_RST,
      O => tx_input_cs_FFd6
    );
  tx_input_cs_FFd6_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd6_FFX_RST
    );
  rx_input_memio_addrchk_bcast_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(2),
      CE => rx_input_memio_addrchk_bcast_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_2_FFY_RST,
      O => rx_input_memio_addrchk_bcast(2)
    );
  rx_input_memio_addrchk_bcast_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_2_FFY_RST
    );
  rx_input_memio_addrchk_bcast_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(4),
      CE => rx_input_memio_addrchk_bcast_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_4_FFY_RST,
      O => rx_input_memio_addrchk_bcast(4)
    );
  rx_input_memio_addrchk_bcast_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_4_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(0),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_0_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(0)
    );
  mac_control_PHY_status_MII_Interface_statecnt_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_0_FFX_RST
    );
  rx_input_memio_addrchk_bcast_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(1),
      CE => rx_input_memio_addrchk_bcast_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_1_FFY_RST,
      O => rx_input_memio_addrchk_bcast(1)
    );
  rx_input_memio_addrchk_bcast_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_1_FFY_RST
    );
  rx_output_ldouten2_1730 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_denll,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_output_invalid,
      O => rx_output_ldouten2
    );
  tx_output_cs_FFd11_1731 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd12,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd12_FFY_RST,
      O => tx_output_cs_FFd11
    );
  tx_output_cs_FFd12_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd12_FFY_RST
    );
  tx_output_cs_FFd16_1732 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd16_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd15_FFY_RST,
      O => tx_output_cs_FFd16
    );
  tx_output_cs_FFd15_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd15_FFY_RST
    );
  tx_output_cs_FFd12_1733 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd13,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd12_FFX_RST,
      O => tx_output_cs_FFd12
    );
  tx_output_cs_FFd12_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd12_FFX_RST
    );
  tx_output_cs_FFd13_1734 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd14,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd14_FFY_RST,
      O => tx_output_cs_FFd13
    );
  tx_output_cs_FFd14_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd14_FFY_RST
    );
  tx_output_cs_FFd14_1735 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd15,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd14_FFX_RST,
      O => tx_output_cs_FFd14
    );
  tx_output_cs_FFd14_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd14_FFX_RST
    );
  mac_control_din_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(25),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_27_FFY_RST,
      O => mac_control_din(26)
    );
  mac_control_din_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_27_FFY_RST
    );
  mac_control_din_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(24),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_25_FFX_RST,
      O => mac_control_din(25)
    );
  mac_control_din_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_25_FFX_RST
    );
  mac_control_din_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(18),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_19_FFX_RST,
      O => mac_control_din(19)
    );
  mac_control_din_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_19_FFX_RST
    );
  mac_control_din_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(26),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_27_FFX_RST,
      O => mac_control_din(27)
    );
  mac_control_din_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_27_FFX_RST
    );
  mac_control_din_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(28),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_29_FFX_RST,
      O => mac_control_din(29)
    );
  mac_control_din_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_29_FFX_RST
    );
  rx_input_memio_cs_FFd15_1736 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd15_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd15_FFY_RST,
      O => rx_input_memio_cs_FFd15
    );
  rx_input_memio_cs_FFd15_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd15_FFY_RST
    );
  tx_output_crcl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(3),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_3_FFY_RST,
      O => tx_output_crcl(3)
    );
  tx_output_crcl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_3_FFY_RST
    );
  mac_control_PHY_status_din_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(1),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_1_FFX_RST,
      O => mac_control_PHY_status_din(1)
    );
  mac_control_PHY_status_din_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_1_FFX_RST
    );
  mac_control_PHY_status_din_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(0),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_1_FFY_RST,
      O => mac_control_PHY_status_din(0)
    );
  mac_control_PHY_status_din_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_1_FFY_RST
    );
  mac_control_PHY_status_din_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(3),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_3_FFX_RST,
      O => mac_control_PHY_status_din(3)
    );
  mac_control_PHY_status_din_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_3_FFX_RST
    );
  mac_control_PHY_status_din_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(5),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_5_FFX_RST,
      O => mac_control_PHY_status_din(5)
    );
  mac_control_PHY_status_din_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_5_FFX_RST
    );
  mac_control_PHY_status_din_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(7),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_7_FFX_RST,
      O => mac_control_PHY_status_din(7)
    );
  mac_control_PHY_status_din_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_7_FFX_RST
    );
  mac_control_PHY_status_din_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(9),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_9_FFX_RST,
      O => mac_control_PHY_status_din(9)
    );
  mac_control_PHY_status_din_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_9_FFX_RST
    );
  rx_output_fifo_nearfull_1737 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_wrcount(1),
      CE => rx_output_fifo_nearfull_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_nearfull_FFY_RST,
      O => rx_output_fifo_nearfull
    );
  rx_output_fifo_nearfull_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifo_nearfull_FFY_RST
    );
  tx_input_MA_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_16,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_1_FFY_RST,
      O => addr4ext(0)
    );
  addr4ext_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_1_FFY_RST
    );
  tx_input_MA_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_17,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_1_FFX_RST,
      O => addr4ext(1)
    );
  addr4ext_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_1_FFX_RST
    );
  tx_input_MA_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_19,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_3_FFX_RST,
      O => addr4ext(3)
    );
  addr4ext_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_3_FFX_RST
    );
  tx_input_MA_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_21,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_5_FFX_RST,
      O => addr4ext(5)
    );
  addr4ext_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_5_FFX_RST
    );
  tx_input_MA_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_23,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_7_FFX_RST,
      O => addr4ext(7)
    );
  addr4ext_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_7_FFX_RST
    );
  tx_input_MD_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(0),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_1_FFY_RST,
      O => d4(0)
    );
  d4_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_1_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(2),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_4_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(3)
    );
  mac_control_PHY_status_MII_Interface_dreg_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_4_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(0),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_2_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(1)
    );
  mac_control_PHY_status_MII_Interface_dreg_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_2_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(1),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_2_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(2)
    );
  mac_control_PHY_status_MII_Interface_dreg_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_2_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(3),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_4_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(4)
    );
  mac_control_PHY_status_MII_Interface_dreg_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_4_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(4),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_6_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(5)
    );
  mac_control_PHY_status_MII_Interface_dreg_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_6_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(5),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_6_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(6)
    );
  mac_control_PHY_status_MII_Interface_dreg_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_6_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(6),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_8_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(7)
    );
  mac_control_PHY_status_MII_Interface_dreg_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_8_FFY_RST
    );
  rx_input_memio_bpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(15),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_15_FFX_RST,
      O => rx_input_memio_bpl(15)
    );
  rx_input_memio_bpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_15_FFX_RST
    );
  rx_input_memio_RXF : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd1,
      CE => rxf_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxf_FFY_RST,
      O => rxf
    );
  rxf_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxf_FFY_RST
    );
  mac_control_phyaddr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_1_FFY_RST,
      O => mac_control_phyaddr(0)
    );
  mac_control_phyaddr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_1_FFY_RST
    );
  mac_control_phyaddr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_1_FFX_RST,
      O => mac_control_phyaddr(1)
    );
  mac_control_phyaddr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_1_FFX_RST
    );
  mac_control_phyaddr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_3_FFX_RST,
      O => mac_control_phyaddr(3)
    );
  mac_control_phyaddr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_3_FFX_RST
    );
  mac_control_phyaddr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_5_FFX_RST,
      O => mac_control_phyaddr(5)
    );
  mac_control_phyaddr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_5_FFX_RST
    );
  mac_control_phyaddr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_7_FFX_RST,
      O => mac_control_phyaddr(7)
    );
  mac_control_phyaddr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_7_FFX_RST
    );
  rx_input_memio_BPOUT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_3_66,
      CE => rxbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_3_FFX_RST,
      O => rxbp(3)
    );
  rxbp_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_3_FFX_RST
    );
  rx_input_memio_BPOUT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_5_64,
      CE => rxbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_5_FFX_RST,
      O => rxbp(5)
    );
  rxbp_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_5_FFX_RST
    );
  rx_input_memio_BPOUT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_7_62,
      CE => rxbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_7_FFX_RST,
      O => rxbp(7)
    );
  rxbp_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_7_FFX_RST
    );
  rx_input_memio_BPOUT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_9_60,
      CE => rxbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_9_FFX_RST,
      O => rxbp(9)
    );
  rxbp_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_9_FFX_RST
    );
  rx_output_FBBP_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(1),
      CE => rxfbbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_1_FFX_RST,
      O => rxfbbp(1)
    );
  rxfbbp_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_1_FFX_RST
    );
  rx_output_FBBP_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(3),
      CE => rxfbbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_3_FFX_RST,
      O => rxfbbp(3)
    );
  rxfbbp_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_3_FFX_RST
    );
  rx_output_FBBP_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(6),
      CE => rxfbbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_7_FFY_RST,
      O => rxfbbp(6)
    );
  rxfbbp_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_7_FFY_RST
    );
  rx_output_FBBP_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(5),
      CE => rxfbbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_5_FFX_RST,
      O => rxfbbp(5)
    );
  rxfbbp_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_5_FFX_RST
    );
  rx_input_memio_cs_FFd7_1738 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd13,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd8_FFY_RST,
      O => rx_input_memio_cs_FFd7
    );
  rx_input_memio_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd8_FFY_RST
    );
  rx_input_memio_cs_FFd8_1739 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd8_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd8_FFX_RST,
      O => rx_input_memio_cs_FFd8
    );
  rx_input_memio_cs_FFd8_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd8_FFX_RST
    );
  rx_input_memio_crcl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(5),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_5_FFX_RST,
      O => rx_input_memio_crcl(5)
    );
  rx_input_memio_crcl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_5_FFX_RST
    );
  tx_input_dh_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(1),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_1_FFX_RST,
      O => tx_input_dh(1)
    );
  tx_input_dh_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_1_FFX_RST
    );
  tx_input_dh_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(3),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_3_FFX_RST,
      O => tx_input_dh(3)
    );
  tx_input_dh_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_3_FFX_RST
    );
  tx_input_dh_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(5),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_5_FFX_RST,
      O => tx_input_dh(5)
    );
  tx_input_dh_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_5_FFX_RST
    );
  tx_input_dh_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(6),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_7_FFY_RST,
      O => tx_input_dh(6)
    );
  tx_input_dh_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_7_FFY_RST
    );
  tx_input_dh_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(7),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_7_FFX_RST,
      O => tx_input_dh(7)
    );
  tx_input_dh_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_7_FFX_RST
    );
  tx_input_dh_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(9),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_9_FFX_RST,
      O => tx_input_dh(9)
    );
  tx_input_dh_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_9_FFX_RST
    );
  tx_input_dl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(1),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_1_FFX_RST,
      O => tx_input_dl(1)
    );
  tx_input_dl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_1_FFX_RST
    );
  tx_input_bp_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_16,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_1_FFY_RST,
      O => txbp(0)
    );
  txbp_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_1_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(0),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_1_FFY_RST,
      O => mac_control_PHY_status_dout(0)
    );
  mac_control_PHY_status_dout_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_1_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(1),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_1_FFX_RST,
      O => mac_control_PHY_status_dout(1)
    );
  mac_control_PHY_status_dout_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_1_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(3),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_3_FFX_RST,
      O => mac_control_PHY_status_dout(3)
    );
  mac_control_PHY_status_dout_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_3_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(5),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_5_FFX_RST,
      O => mac_control_PHY_status_dout(5)
    );
  mac_control_PHY_status_dout_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_5_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(7),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_7_FFX_RST,
      O => mac_control_PHY_status_dout(7)
    );
  mac_control_PHY_status_dout_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_7_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(9),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_9_FFX_RST,
      O => mac_control_PHY_status_dout(9)
    );
  mac_control_PHY_status_dout_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_9_FFX_RST
    );
  rx_input_memio_bpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(10),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_11_FFY_RST,
      O => rx_input_memio_bpl(10)
    );
  rx_input_memio_bpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_11_FFY_RST
    );
  rx_input_memio_bpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(11),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_11_FFX_RST,
      O => rx_input_memio_bpl(11)
    );
  rx_input_memio_bpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_11_FFX_RST
    );
  rx_input_memio_bpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(14),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_15_FFY_RST,
      O => rx_input_memio_bpl(14)
    );
  rx_input_memio_bpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_15_FFY_RST
    );
  rx_input_memio_bpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(13),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_13_FFX_RST,
      O => rx_input_memio_bpl(13)
    );
  rx_input_memio_bpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_13_FFX_RST
    );
  tx_input_bp_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_17,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_1_FFX_RST,
      O => txbp(1)
    );
  txbp_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_1_FFX_RST
    );
  tx_input_dl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(3),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_3_FFX_RST,
      O => tx_input_dl(3)
    );
  tx_input_dl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_3_FFX_RST
    );
  tx_input_bp_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_18,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_3_FFY_RST,
      O => txbp(2)
    );
  txbp_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_3_FFY_RST
    );
  tx_input_bp_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_19,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_3_FFX_RST,
      O => txbp(3)
    );
  txbp_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_3_FFX_RST
    );
  tx_input_dl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(5),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_5_FFX_RST,
      O => tx_input_dl(5)
    );
  tx_input_dl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_5_FFX_RST
    );
  tx_input_bp_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_20,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_5_FFY_RST,
      O => txbp(4)
    );
  txbp_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_5_FFY_RST
    );
  tx_input_bp_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_21,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_5_FFX_RST,
      O => txbp(5)
    );
  txbp_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_5_FFX_RST
    );
  tx_input_dl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(7),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_7_FFX_RST,
      O => tx_input_dl(7)
    );
  tx_input_dl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_7_FFX_RST
    );
  tx_input_bp_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_22,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_7_FFY_RST,
      O => txbp(6)
    );
  txbp_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_7_FFY_RST
    );
  tx_input_bp_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_23,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_7_FFX_RST,
      O => txbp(7)
    );
  txbp_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_7_FFX_RST
    );
  tx_input_dl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(9),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_9_FFX_RST,
      O => tx_input_dl(9)
    );
  tx_input_dl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_9_FFX_RST
    );
  tx_input_bp_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_24,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_9_FFY_RST,
      O => txbp(8)
    );
  txbp_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_9_FFY_RST
    );
  rx_input_memio_dout_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_5_FFX_RST,
      O => rx_input_memio_dout(5)
    );
  rx_input_memio_dout_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_5_FFX_RST
    );
  tx_output_FBBP_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(15),
      CE => txfbbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_15_FFX_RST,
      O => txfbbp(15)
    );
  txfbbp_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_15_FFX_RST
    );
  rx_input_memio_dout_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_7_FFX_RST,
      O => rx_input_memio_dout(7)
    );
  rx_input_memio_dout_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_7_FFX_RST
    );
  rx_input_memio_dout_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_9_FFX_RST,
      O => rx_input_memio_dout(9)
    );
  rx_input_memio_dout_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_9_FFX_RST
    );
  rx_input_fifo_control_DATA_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(0),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_0_FFY_RST,
      O => rx_input_data(0)
    );
  rx_input_data_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_0_FFY_RST
    );
  rx_output_cs_FFd9_1740 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd9_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd9_FFY_RST,
      O => rx_output_cs_FFd9
    );
  rx_output_cs_FFd9_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd9_FFY_RST
    );
  tx_output_crcl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(5),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_5_FFX_RST,
      O => tx_output_crcl(5)
    );
  tx_output_crcl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_5_FFX_RST
    );
  tx_output_crcl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(4),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_4_FFY_RST,
      O => tx_output_crcl(4)
    );
  tx_output_crcl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_4_FFY_RST
    );
  tx_output_outsell_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => tx_output_outsel_0_Q,
      CE => tx_output_outsell_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => tx_output_outsell_0_FFY_SET,
      RST => GND,
      O => tx_output_outsell(0)
    );
  tx_output_outsell_0_FFY_SETOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outsell_0_FFY_SET
    );
  mac_control_PHY_status_rwl_1741 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(5),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_rwl_FFY_RST,
      O => mac_control_PHY_status_rwl
    );
  mac_control_PHY_status_rwl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_rwl_FFY_RST
    );
  rx_input_GMII_rx_of_1742 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_rx_nearf,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_GMII_rx_of_FFY_RST,
      O => rx_input_GMII_rx_of
    );
  rx_input_GMII_rx_of_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_GMII_rx_of_FFY_RST
    );
  mac_control_phyaddr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_9_FFX_RST,
      O => mac_control_phyaddr(9)
    );
  mac_control_phyaddr_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_9_FFX_RST
    );
  rx_input_memio_crcrst_1743 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd16,
      CE => rx_input_memio_crcrst_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcrst_FFY_RST,
      O => rx_input_memio_crcrst
    );
  rx_input_memio_crcrst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcrst_FFY_RST
    );
  mac_control_sclkll_1744 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_sclkl,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_sclkll_FFY_RST,
      O => mac_control_sclkll
    );
  mac_control_sclkll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_sclkll_FFY_RST
    );
  rx_input_memio_dout_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_1_FFX_RST,
      O => rx_input_memio_dout(1)
    );
  rx_input_memio_dout_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_1_FFX_RST
    );
  tx_output_FBBP_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(11),
      CE => txfbbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_11_FFX_RST,
      O => txfbbp(11)
    );
  txfbbp_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_11_FFX_RST
    );
  rx_input_memio_dout_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_3_FFX_RST,
      O => rx_input_memio_dout(3)
    );
  rx_input_memio_dout_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_3_FFX_RST
    );
  rx_input_memio_dout_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_5_FFY_RST,
      O => rx_input_memio_dout(4)
    );
  rx_input_memio_dout_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_5_FFY_RST
    );
  tx_output_FBBP_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(13),
      CE => txfbbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_13_FFX_RST,
      O => txfbbp(13)
    );
  txfbbp_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_13_FFX_RST
    );
  rx_input_fifo_control_DATA_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(1),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_1_FFY_RST,
      O => rx_input_data(1)
    );
  rx_input_data_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_1_FFY_RST
    );
  rx_input_fifo_control_DATA_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(2),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_2_FFY_RST,
      O => rx_input_data(2)
    );
  rx_input_data_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_2_FFY_RST
    );
  rx_input_fifo_control_DATA_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(3),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_3_FFY_RST,
      O => rx_input_data(3)
    );
  rx_input_data_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_3_FFY_RST
    );
  rx_input_fifo_control_DATA_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(4),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_4_FFY_RST,
      O => rx_input_data(4)
    );
  rx_input_data_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_4_FFY_RST
    );
  rx_input_fifo_control_DATA_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(5),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_5_FFY_RST,
      O => rx_input_data(5)
    );
  rx_input_data_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_5_FFY_RST
    );
  rx_input_fifo_control_DATA_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(6),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_6_FFY_RST,
      O => rx_input_data(6)
    );
  rx_input_data_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_6_FFY_RST
    );
  rx_input_fifo_control_DATA_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(7),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_7_FFY_RST,
      O => rx_input_data(7)
    );
  rx_input_data_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_7_FFY_RST
    );
  rx_input_fifo_control_ENDF : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(8),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_endf_FFY_RST,
      O => rx_input_endf
    );
  rx_input_endf_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_endf_FFY_RST
    );
  rx_input_fifo_control_INVALID : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(9),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_invalid_FFY_RST,
      O => rx_input_invalid
    );
  rx_input_invalid_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_invalid_FFY_RST
    );
  tx_input_fifofulll_1745 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfifofull,
      CE => tx_input_fifofulll_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_fifofulll_FFY_RST,
      O => tx_input_fifofulll
    );
  tx_input_fifofulll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_fifofulll_FFY_RST
    );
  rx_input_memio_crcequal_1746 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_N80267,
      CE => rx_input_memio_crcequal_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcequal_FFY_RST,
      O => rx_input_memio_crcequal
    );
  rx_input_memio_crcequal_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcequal_FFY_RST
    );
  mac_control_dout_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N77583,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_10_FFY_RST,
      O => mac_control_dout(10)
    );
  mac_control_dout_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_10_FFY_RST
    );
  mac_control_PHY_status_phyaddrws_1747 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_phyaddrws_BYMUXNOT,
      CE => mac_control_PHY_status_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_phyaddrws_FFY_RST,
      O => mac_control_PHY_status_phyaddrws
    );
  mac_control_PHY_status_phyaddrws_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_phyaddrws_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(9),
      CE => rx_input_memio_addrchk_macaddrl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_9_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(9)
    );
  rx_input_memio_addrchk_macaddrl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_9_FFX_RST
    );
  rx_output_lenr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(2),
      CE => rx_output_lenr_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_2_FFY_RST,
      O => rx_output_lenr(2)
    );
  rx_output_lenr_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_2_FFY_RST
    );
  rx_input_memio_crcl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(25),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_25_FFY_RST,
      O => rx_input_memio_crcl(25)
    );
  rx_input_memio_crcl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_25_FFY_RST
    );
  mac_control_txf_cross_1748 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfsr,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_txf_cross_FFY_RST,
      O => mac_control_txf_cross
    );
  mac_control_txf_cross_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cross_FFY_RST
    );
  rx_output_lenr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(3),
      CE => rx_output_lenr_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_3_FFY_RST,
      O => rx_output_lenr(3)
    );
  rx_output_lenr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_3_FFY_RST
    );
  rx_output_fifo_BU378 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1553,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1585_FFX_RST,
      O => rx_output_fifo_N1585
    );
  rx_output_fifo_N1585_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1585_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(7),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_23_FFX_RST,
      O => mac_control_phystat(23)
    );
  mac_control_phystat_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_23_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(15),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_31_FFX_RST,
      O => mac_control_phystat(31)
    );
  mac_control_phystat_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_31_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(14),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_15_FFY_RST,
      O => mac_control_phystat(14)
    );
  mac_control_phystat_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_15_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(15),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_15_FFX_RST,
      O => mac_control_phystat(15)
    );
  mac_control_phystat_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_15_FFX_RST
    );
  rx_output_fifo_BU346 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1563,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1571_FFX_RST,
      O => rx_output_fifo_N1571
    );
  rx_output_fifo_N1571_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1571_FFX_RST
    );
  memcontroller_Q2_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(29),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_29_FFX_RST,
      O => q2(29)
    );
  q2_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_29_FFX_RST
    );
  memcontroller_Q3_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(21),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_21_FFX_RST,
      O => q3(21)
    );
  q3_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_21_FFX_RST
    );
  memcontroller_Q3_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(13),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_13_FFX_RST,
      O => q3(13)
    );
  q3_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_13_FFX_RST
    );
  rx_output_fifo_BU470 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1578,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1586_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1586
    );
  rx_output_fifo_N1586_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1586_FFX_SET
    );
  tx_input_MA_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_25,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_9_FFX_RST,
      O => addr4ext(9)
    );
  addr4ext_9_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_9_FFX_RST
    );
  tx_input_MD_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(1),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_1_FFX_RST,
      O => d4(1)
    );
  d4_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_1_FFX_RST
    );
  tx_input_MD_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(3),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_3_FFX_RST,
      O => d4(3)
    );
  d4_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_3_FFX_RST
    );
  tx_input_MD_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(5),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_5_FFX_RST,
      O => d4(5)
    );
  d4_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_5_FFX_RST
    );
  tx_input_MD_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(7),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_7_FFX_RST,
      O => d4(7)
    );
  d4_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_7_FFX_RST
    );
  tx_input_MD_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(9),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_9_FFX_RST,
      O => d4(9)
    );
  d4_9_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_9_FFX_RST
    );
  tx_fifocheck_fbbpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_11_FFX_RST,
      O => tx_fifocheck_fbbpl(11)
    );
  tx_fifocheck_fbbpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_11_FFX_RST
    );
  tx_fifocheck_fbbpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_13_FFX_RST,
      O => tx_fifocheck_fbbpl(13)
    );
  tx_fifocheck_fbbpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_13_FFX_RST
    );
  tx_fifocheck_fbbpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_15_FFX_RST,
      O => tx_fifocheck_fbbpl(15)
    );
  tx_fifocheck_fbbpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_15_FFX_RST
    );
  rx_output_fifo_BU368 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N5,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1605_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1605
    );
  rx_output_fifo_N1605_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1605_FFX_SET
    );
  rx_output_fifo_BU360 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N9,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1609_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1609
    );
  rx_output_fifo_N1609_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1609_FFX_SET
    );
  mac_control_PHY_status_PHYSTAT_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(5),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_21_FFX_RST,
      O => mac_control_phystat(21)
    );
  mac_control_phystat_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_21_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(13),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_13_FFX_RST,
      O => mac_control_phystat(13)
    );
  mac_control_phystat_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_13_FFX_RST
    );
  memcontroller_Q2_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(27),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_27_FFX_RST,
      O => q2(27)
    );
  q2_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_27_FFX_RST
    );
  memcontroller_Q2_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(19),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_19_FFX_RST,
      O => q2(19)
    );
  q2_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_19_FFX_RST
    );
  memcontroller_Q3_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(11),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_11_FFX_RST,
      O => q3(11)
    );
  q3_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_11_FFX_RST
    );
  rx_input_memio_addrchk_cs_FFd2_1749 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd2_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd2_FFX_RST,
      O => rx_input_memio_addrchk_cs_FFd2
    );
  rx_input_memio_addrchk_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd2_FFX_RST
    );
  tx_output_crcl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(6),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_6_FFY_RST,
      O => tx_output_crcl(6)
    );
  tx_output_crcl_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_6_FFY_RST
    );
  rx_input_memio_addrchk_cs_FFd6_1750 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd6_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd6_FFY_RST,
      O => rx_input_memio_addrchk_cs_FFd6
    );
  rx_input_memio_addrchk_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd6_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd2_1751 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd2_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_cs_FFd2_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_cs_FFd2
    );
  mac_control_PHY_status_MII_Interface_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_MII_Interface_cs_FFd2_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(1),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_1_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(1)
    );
  mac_control_PHY_status_MII_Interface_statecnt_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_1_FFY_RST
    );
  mac_control_MACADDR_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(0),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_1_FFY_RST,
      O => macaddr(0)
    );
  macaddr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_1_FFY_RST
    );
  mac_control_MACADDR_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(1),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_1_FFX_RST,
      O => macaddr(1)
    );
  macaddr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_1_FFX_RST
    );
  mac_control_MACADDR_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(3),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_3_FFX_RST,
      O => macaddr(3)
    );
  macaddr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_3_FFX_RST
    );
  mac_control_MACADDR_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(5),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_5_FFX_RST,
      O => macaddr(5)
    );
  macaddr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_5_FFX_RST
    );
  mac_control_MACADDR_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(7),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_7_FFX_RST,
      O => macaddr(7)
    );
  macaddr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_7_FFX_RST
    );
  mac_control_MACADDR_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(9),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_9_FFX_RST,
      O => macaddr(9)
    );
  macaddr_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_9_FFX_RST
    );
  tx_output_crcl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(7),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_7_FFY_RST,
      O => tx_output_crcl(7)
    );
  tx_output_crcl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_7_FFY_RST
    );
  rx_output_mdl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(25),
      CE => rx_output_mdl_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_25_FFX_RST,
      O => rx_output_mdl(25)
    );
  rx_output_mdl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_25_FFX_RST
    );
  rx_output_mdl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(17),
      CE => rx_output_mdl_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_17_FFX_RST,
      O => rx_output_mdl(17)
    );
  rx_output_mdl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_17_FFX_RST
    );
  rx_output_mdl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(26),
      CE => rx_output_mdl_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_27_FFY_RST,
      O => rx_output_mdl(26)
    );
  rx_output_mdl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_27_FFY_RST
    );
  rx_output_mdl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(27),
      CE => rx_output_mdl_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_27_FFX_RST,
      O => rx_output_mdl(27)
    );
  rx_output_mdl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_27_FFX_RST
    );
  rx_output_mdl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(19),
      CE => rx_output_mdl_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_19_FFX_RST,
      O => rx_output_mdl(19)
    );
  rx_output_mdl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_19_FFX_RST
    );
  rx_output_mdl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(29),
      CE => rx_output_mdl_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_29_FFX_RST,
      O => rx_output_mdl(29)
    );
  rx_output_mdl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_29_FFX_RST
    );
  tx_output_cs_FFd1_1752 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd2,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd2_FFY_RST,
      O => tx_output_cs_FFd1
    );
  tx_output_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd2_FFY_RST
    );
  tx_output_cs_FFd4_1753 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd3_FFY_RST,
      O => tx_output_cs_FFd4
    );
  tx_output_cs_FFd3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd3_FFY_RST
    );
  memcontroller_dnl1_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(5),
      CE => memcontroller_dnl1_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_5_FFX_RST,
      O => memcontroller_dnl1(5)
    );
  memcontroller_dnl1_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_5_FFX_RST
    );
  memcontroller_dnl1_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(13),
      CE => memcontroller_dnl1_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_13_FFX_RST,
      O => memcontroller_dnl1(13)
    );
  memcontroller_dnl1_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_13_FFX_RST
    );
  memcontroller_dnl1_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(14),
      CE => memcontroller_dnl1_14_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_14_FFX_RST,
      O => memcontroller_dnl1(14)
    );
  memcontroller_dnl1_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_14_FFX_RST
    );
  memcontroller_dnl1_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(6),
      CE => memcontroller_dnl1_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_6_FFX_RST,
      O => memcontroller_dnl1(6)
    );
  memcontroller_dnl1_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_6_FFX_RST
    );
  memcontroller_dnl1_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(7),
      CE => memcontroller_dnl1_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_7_FFX_RST,
      O => memcontroller_dnl1(7)
    );
  memcontroller_dnl1_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_7_FFX_RST
    );
  memcontroller_dnout_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_5_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_5_OFF_RST,
      O => memcontroller_dnout(5)
    );
  MD_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_5_OFF_RST
    );
  memcontroller_ts_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_5_TFF_RST,
      O => memcontroller_ts(5)
    );
  MD_5_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_5_TFF_RST
    );
  memcontroller_dnout_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_6_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_6_OFF_RST,
      O => memcontroller_dnout(6)
    );
  MD_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_6_OFF_RST
    );
  memcontroller_ts_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_6_TFF_RST,
      O => memcontroller_ts(6)
    );
  MD_6_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_6_TFF_RST
    );
  memcontroller_qn_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_7_IFF_RST,
      O => memcontroller_qn(7)
    );
  MD_7_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_7_IFF_RST
    );
  memcontroller_dnout_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_7_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_7_OFF_RST,
      O => memcontroller_dnout(7)
    );
  MD_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_7_OFF_RST
    );
  memcontroller_ts_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_7_TFF_RST,
      O => memcontroller_ts(7)
    );
  MD_7_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_7_TFF_RST
    );
  memcontroller_qn_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_8_IFF_RST,
      O => memcontroller_qn(8)
    );
  MD_8_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_8_IFF_RST
    );
  memcontroller_qn_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_9_IFF_RST,
      O => memcontroller_qn(9)
    );
  MD_9_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_9_IFF_RST
    );
  memcontroller_dnout_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_8_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_8_OFF_RST,
      O => memcontroller_dnout(8)
    );
  MD_8_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_8_OFF_RST
    );
  memcontroller_ts_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_8_TFF_RST,
      O => memcontroller_ts(8)
    );
  MD_8_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_8_TFF_RST
    );
  memcontroller_dnout_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_9_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_9_OFF_RST,
      O => memcontroller_dnout(9)
    );
  MD_9_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_9_OFF_RST
    );
  memcontroller_ts_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_9_TFF_RST,
      O => memcontroller_ts(9)
    );
  MD_9_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_9_TFF_RST
    );
  tx_output_addr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(1),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_0_FFY_RST,
      O => addr2ext(1)
    );
  addr2ext_0_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_0_FFY_RST
    );
  tx_output_addr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(3),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_2_FFY_RST,
      O => addr2ext(3)
    );
  addr2ext_2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_2_FFY_RST
    );
  tx_output_addr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(7),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_6_FFY_RST,
      O => addr2ext(7)
    );
  addr2ext_6_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_6_FFY_RST
    );
  tx_output_addr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_Madd_n0000_inst_lut2_0,
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_0_FFX_RST,
      O => addr2ext(0)
    );
  addr2ext_0_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_0_FFX_RST
    );
  tx_output_addr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(2),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_2_FFX_RST,
      O => addr2ext(2)
    );
  addr2ext_2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_2_FFX_RST
    );
  tx_output_addr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(5),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_4_FFY_RST,
      O => addr2ext(5)
    );
  addr2ext_4_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_4_FFY_RST
    );
  memcontroller_dnl1_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(15),
      CE => memcontroller_dnl1_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_15_FFX_RST,
      O => memcontroller_dnl1(15)
    );
  memcontroller_dnl1_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_15_FFX_RST
    );
  memcontroller_dnl1_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(23),
      CE => memcontroller_dnl1_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_23_FFX_RST,
      O => memcontroller_dnl1(23)
    );
  memcontroller_dnl1_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_23_FFX_RST
    );
  memcontroller_dnl1_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(0),
      CE => memcontroller_dnl1_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_0_FFX_RST,
      O => memcontroller_dnl1(0)
    );
  memcontroller_dnl1_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_0_FFX_RST
    );
  memcontroller_dnl1_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(8),
      CE => memcontroller_dnl1_8_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_8_FFX_RST,
      O => memcontroller_dnl1(8)
    );
  memcontroller_dnl1_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_8_FFX_RST
    );
  memcontroller_dnl1_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(16),
      CE => memcontroller_dnl1_16_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_16_FFX_RST,
      O => memcontroller_dnl1(16)
    );
  memcontroller_dnl1_16_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_16_FFX_RST
    );
  rx_output_lenr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(4),
      CE => rx_output_lenr_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_4_FFY_RST,
      O => rx_output_lenr(4)
    );
  rx_output_lenr_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_4_FFY_RST
    );
  rx_output_denl_1754 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_CHOICE1529,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => GSR,
      SSET => rx_output_CHOICE1525,
      SRST => rx_output_denl_LOGIC_ZERO,
      O => rx_output_denl
    );
  rx_output_lenr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(5),
      CE => rx_output_lenr_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_5_FFY_RST,
      O => rx_output_lenr(5)
    );
  rx_output_lenr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_5_FFY_RST
    );
  mac_control_RXBCAST : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lrxbcast,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbcast_FFY_RST,
      O => rxbcast
    );
  rxbcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbcast_FFY_RST
    );
  mac_control_dout_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N77791,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_14_FFY_RST,
      O => mac_control_dout(14)
    );
  mac_control_dout_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_14_FFY_RST
    );
  rx_output_bpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(5),
      CE => rx_output_bpl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_5_FFX_RST,
      O => rx_output_bpl(5)
    );
  rx_output_bpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_5_FFX_RST
    );
  tx_output_datal_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(3),
      CE => tx_output_datal_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_3_FFX_RST,
      O => tx_output_datal(3)
    );
  tx_output_datal_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_3_FFX_RST
    );
  rx_output_bpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(7),
      CE => rx_output_bpl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_7_FFX_RST,
      O => rx_output_bpl(7)
    );
  rx_output_bpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_7_FFX_RST
    );
  tx_output_datal_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(5),
      CE => tx_output_datal_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_5_FFX_RST,
      O => tx_output_datal(5)
    );
  tx_output_datal_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_5_FFX_RST
    );
  rx_output_bpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(9),
      CE => rx_output_bpl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_9_FFX_RST,
      O => rx_output_bpl(9)
    );
  rx_output_bpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_9_FFX_RST
    );
  rx_output_bpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(8),
      CE => rx_output_bpl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_9_FFY_RST,
      O => rx_output_bpl(8)
    );
  rx_output_bpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_9_FFY_RST
    );
  tx_output_datal_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(7),
      CE => tx_output_datal_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_7_FFX_RST,
      O => tx_output_datal(7)
    );
  tx_output_datal_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_7_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(7),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_8_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(8)
    );
  mac_control_PHY_status_MII_Interface_dreg_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_8_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(8),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_10_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(9)
    );
  mac_control_PHY_status_MII_Interface_dreg_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_10_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(9),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_10_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(10)
    );
  mac_control_PHY_status_MII_Interface_dreg_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_10_FFX_RST
    );
  tx_output_crcl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(0),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_0_FFY_RST,
      O => tx_output_crcl(0)
    );
  tx_output_crcl_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_0_FFY_RST
    );
  slowclock_txfl_1755 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_txfl_GROM,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => txf,
      SRST => slowclock_txfl_LOGIC_ZERO,
      O => slowclock_txfl
    );
  slowclock_rxfl_1756 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_rxfl_GROM,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => rxf,
      SRST => slowclock_rxfl_LOGIC_ZERO,
      O => slowclock_rxfl
    );
  tx_input_dh_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(0),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_1_FFY_RST,
      O => tx_input_dh(0)
    );
  tx_input_dh_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_1_FFY_RST
    );
  mac_control_bitcnt_109_1757 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_256,
      CE => mac_control_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_bitcnt_109_FFX_RST,
      O => mac_control_bitcnt_109
    );
  mac_control_bitcnt_109_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_109_FFX_RST
    );
  tx_input_cs_FFd1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd2,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_DONE_FFY_RST,
      O => tx_input_DONE
    );
  tx_input_DONE_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_DONE_FFY_RST
    );
  mac_control_SOUT : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => SOUT_OD,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => SOUT_OFF_RST,
      O => mac_control_SOUT_OBUF
    );
  SOUT_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => SOUT_OFF_RST
    );
  mac_control_sclkl_1758 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_SCLK_IBUF,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => SCLK_IFF_RST,
      O => mac_control_sclkl
    );
  SCLK_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => SCLK_IFF_RST
    );
  mac_control_LEDRX : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDRX_OD,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => LEDRX_OFF_RST,
      O => mac_control_LEDRX_OBUF
    );
  LEDRX_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDRX_OFF_RST
    );
  mac_control_LEDTX : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDTX_OD,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => LEDTX_OFF_RST,
      O => mac_control_LEDTX_OBUF
    );
  LEDTX_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDTX_OFF_RST
    );
  tx_input_dinl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_0_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_0_IFF_RST,
      O => tx_input_dinl(0)
    );
  DIN_0_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_0_IFF_RST
    );
  tx_input_dinl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_1_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_1_IFF_RST,
      O => tx_input_dinl(1)
    );
  DIN_1_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_1_IFF_RST
    );
  tx_input_dinl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_2_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_2_IFF_RST,
      O => tx_input_dinl(2)
    );
  DIN_2_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_2_IFF_RST
    );
  rx_input_memio_addrchk_validucast_1759 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_n0052,
      CE => rx_input_memio_addrchk_validucast_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_validucast_FFY_RST,
      O => rx_input_memio_addrchk_validucast
    );
  rx_input_memio_addrchk_validucast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_validucast_FFY_RST
    );
  mac_control_RXMCAST : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lrxmcast,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxmcast_FFY_RST,
      O => rxmcast
    );
  rxmcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxmcast_FFY_RST
    );
  mac_control_RXUCAST : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lrxucast,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxucast_FFY_RST,
      O => rxucast
    );
  rxucast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxucast_FFY_RST
    );
  rx_input_memio_crcl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(30),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_30_FFY_RST,
      O => rx_input_memio_crcl(30)
    );
  rx_input_memio_crcl_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_30_FFY_RST
    );
  rx_input_memio_addrchk_cs_FFd7_1760 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd7_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_memio_addrchk_cs_FFd7_FFX_SET,
      RST => GND,
      O => rx_input_memio_addrchk_cs_FFd7
    );
  rx_input_memio_addrchk_cs_FFd7_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_RESET_1,
      O => rx_input_memio_addrchk_cs_FFd7_FFX_SET
    );
  rx_input_memio_addrchk_cs_FFd5_1761 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd5_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd5_FFX_RST,
      O => rx_input_memio_addrchk_cs_FFd5
    );
  rx_input_memio_addrchk_cs_FFd5_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd5_FFX_RST
    );
  tx_output_addrl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(10),
      CE => tx_output_addrl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_11_FFY_RST,
      O => tx_output_addrl(10)
    );
  tx_output_addrl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_11_FFY_RST
    );
  tx_output_addrl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(11),
      CE => tx_output_addrl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_11_FFX_RST,
      O => tx_output_addrl(11)
    );
  tx_output_addrl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_11_FFX_RST
    );
  tx_output_addrl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(12),
      CE => tx_output_addrl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_13_FFY_RST,
      O => tx_output_addrl(12)
    );
  tx_output_addrl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_13_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(13),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_13_FFX_RST,
      O => mac_control_PHY_status_dout(13)
    );
  mac_control_PHY_status_dout_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_13_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(15),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_15_FFX_RST,
      O => mac_control_PHY_status_dout(15)
    );
  mac_control_PHY_status_dout_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_15_FFX_RST
    );
  tx_output_ncrcbytel_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(1),
      CE => tx_output_ncrcbytel_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_1_FFY_RST,
      O => tx_output_ncrcbytel(1)
    );
  tx_output_ncrcbytel_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_1_FFY_RST
    );
  tx_output_ncrcbytel_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(2),
      CE => tx_output_ncrcbytel_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_2_FFY_RST,
      O => tx_output_ncrcbytel(2)
    );
  tx_output_ncrcbytel_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_2_FFY_RST
    );
  tx_output_ncrcbytel_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(3),
      CE => tx_output_ncrcbytel_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_3_FFY_RST,
      O => tx_output_ncrcbytel(3)
    );
  tx_output_ncrcbytel_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_3_FFY_RST
    );
  tx_output_addrl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(13),
      CE => tx_output_addrl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_13_FFX_RST,
      O => tx_output_addrl(13)
    );
  tx_output_addrl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_13_FFX_RST
    );
  rx_input_memio_addrchk_bcast_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(3),
      CE => rx_input_memio_addrchk_bcast_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_3_FFY_RST,
      O => rx_input_memio_addrchk_bcast(3)
    );
  rx_input_memio_addrchk_bcast_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_3_FFY_RST
    );
  slowclock_TXFIFOWERRSR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_txfifowerrl,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfifowerrsr_FFY_RST,
      O => txfifowerrsr
    );
  txfifowerrsr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfifowerrsr_FFY_RST
    );
  tx_output_addrl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(14),
      CE => tx_output_addrl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_15_FFY_RST,
      O => tx_output_addrl(14)
    );
  tx_output_addrl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_15_FFY_RST
    );
  tx_output_addrl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(15),
      CE => tx_output_addrl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_15_FFX_RST,
      O => tx_output_addrl(15)
    );
  tx_output_addrl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_15_FFX_RST
    );
  rx_input_memio_addrchk_bcast_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(0),
      CE => rx_input_memio_addrchk_bcast_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_0_FFY_RST,
      O => rx_input_memio_addrchk_bcast(0)
    );
  rx_input_memio_addrchk_bcast_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_0_FFY_RST
    );
  rx_input_memio_addrchk_bcast_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(5),
      CE => rx_input_memio_addrchk_bcast_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_5_FFY_RST,
      O => rx_input_memio_addrchk_bcast(5)
    );
  rx_input_memio_addrchk_bcast_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_5_FFY_RST
    );
  rx_output_lenr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(9),
      CE => rx_output_lenr_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_9_FFY_RST,
      O => rx_output_lenr(9)
    );
  rx_output_lenr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_9_FFY_RST
    );
  rx_input_memio_addrchk_mcast_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmcast(0),
      CE => rx_input_memio_addrchk_mcast_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_mcast_0_FFY_RST,
      O => rx_input_memio_addrchk_mcast(0)
    );
  rx_input_memio_addrchk_mcast_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_mcast_0_FFY_RST
    );
  tx_output_ncrcbytel_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(0),
      CE => tx_output_ncrcbytel_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_0_FFY_RST,
      O => tx_output_ncrcbytel(0)
    );
  tx_output_ncrcbytel_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_0_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(10),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_11_FFY_RST,
      O => mac_control_PHY_status_dout(10)
    );
  mac_control_PHY_status_dout_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_11_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(11),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_11_FFX_RST,
      O => mac_control_PHY_status_dout(11)
    );
  mac_control_PHY_status_dout_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_11_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(12),
      CE => mac_control_PHY_status_MII_Interface_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_13_FFY_RST,
      O => mac_control_PHY_status_dout(12)
    );
  mac_control_PHY_status_dout_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_13_FFY_RST
    );
  tx_output_crcl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(1),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_1_FFY_RST,
      O => tx_output_crcl(1)
    );
  tx_output_crcl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_1_FFY_RST
    );
  rx_output_lenr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(7),
      CE => rx_output_lenr_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_7_FFY_RST,
      O => rx_output_lenr(7)
    );
  rx_output_lenr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_7_FFY_RST
    );
  mac_control_dout_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N74276,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_31_FFY_RST,
      O => mac_control_dout(31)
    );
  mac_control_dout_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_31_FFY_RST
    );
  mac_control_dout_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N74572,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_23_FFY_RST,
      O => mac_control_dout(23)
    );
  mac_control_dout_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_23_FFY_RST
    );
  rx_output_lenr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(8),
      CE => rx_output_lenr_8_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_8_FFY_RST,
      O => rx_output_lenr(8)
    );
  rx_output_lenr_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_8_FFY_RST
    );
  tx_output_bcntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_49,
      CE => tx_output_bcntl_12_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_12_FFY_RST,
      O => tx_output_bcntl(11)
    );
  tx_output_bcntl_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_12_FFY_RST
    );
  tx_output_bcntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_50,
      CE => tx_output_bcntl_12_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_12_FFX_RST,
      O => tx_output_bcntl(12)
    );
  tx_output_bcntl_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_12_FFX_RST
    );
  tx_output_bcntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_52,
      CE => tx_output_bcntl_14_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_14_FFX_RST,
      O => tx_output_bcntl(14)
    );
  tx_output_bcntl_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_14_FFX_RST
    );
  rx_output_bpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(10),
      CE => rx_output_bpl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_11_FFY_RST,
      O => rx_output_bpl(10)
    );
  rx_output_bpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_11_FFY_RST
    );
  rx_output_bpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(11),
      CE => rx_output_bpl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_11_FFX_RST,
      O => rx_output_bpl(11)
    );
  rx_output_bpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_11_FFX_RST
    );
  rx_output_bpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(13),
      CE => rx_output_bpl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_13_FFX_RST,
      O => rx_output_bpl(13)
    );
  rx_output_bpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_13_FFX_RST
    );
  rx_output_bpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(15),
      CE => rx_output_bpl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_15_FFX_RST,
      O => rx_output_bpl(15)
    );
  rx_output_bpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_15_FFX_RST
    );
  tx_output_cs_FFd15_1762 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd16,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd15_FFX_RST,
      O => tx_output_cs_FFd15
    );
  tx_output_cs_FFd15_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd15_FFX_RST
    );
  rx_input_memio_crcl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(1),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_1_FFY_RST,
      O => rx_input_memio_crcl(1)
    );
  rx_input_memio_crcl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_1_FFY_RST
    );
  tx_output_crcl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(30),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_30_FFY_RST,
      O => tx_output_crcl(30)
    );
  tx_output_crcl_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_30_FFY_RST
    );
  rx_input_memio_crcen_1763 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0049,
      CE => rx_input_memio_crcen_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcen_FFX_RST,
      O => rx_input_memio_crcen
    );
  rx_input_memio_crcen_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcen_FFX_RST
    );
  tx_fifocheck_fbbpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_7_FFX_RST,
      O => tx_fifocheck_fbbpl(7)
    );
  tx_fifocheck_fbbpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_7_FFX_RST
    );
  tx_fifocheck_fbbpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_9_FFX_RST,
      O => tx_fifocheck_fbbpl(9)
    );
  tx_fifocheck_fbbpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_9_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(11),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_11_FFX_RST,
      O => mac_control_phydo(11)
    );
  mac_control_phydo_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_11_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(13),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_13_FFX_RST,
      O => mac_control_phydo(13)
    );
  mac_control_phydo_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_13_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(15),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_15_FFX_RST,
      O => mac_control_phydo(15)
    );
  mac_control_phydo_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_15_FFX_RST
    );
  tx_output_ltxen2_1764 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ltxen,
      CE => tx_output_ltxen3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ltxen3_FFY_RST,
      O => tx_output_ltxen2
    );
  tx_output_ltxen3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ltxen3_FFY_RST
    );
  tx_output_ltxen3_1765 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ltxen2,
      CE => tx_output_ltxen3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ltxen3_FFX_RST,
      O => tx_output_ltxen3
    );
  tx_output_ltxen3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ltxen3_FFX_RST
    );
  slowclock_lclken_1766 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_lclken_LOGIC_ONE,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => slowclock_n0005,
      O => slowclock_lclken
    );
  rx_input_memio_crcl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(0),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_0_FFY_RST,
      O => rx_input_memio_crcl(0)
    );
  rx_input_memio_crcl_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_0_FFY_RST
    );
  tx_fifocheck_fbbpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_1_FFX_RST,
      O => tx_fifocheck_fbbpl(1)
    );
  tx_fifocheck_fbbpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_1_FFX_RST
    );
  tx_fifocheck_fbbpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_1_FFY_RST,
      O => tx_fifocheck_fbbpl(0)
    );
  tx_fifocheck_fbbpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_1_FFY_RST
    );
  tx_fifocheck_fbbpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_3_FFX_RST,
      O => tx_fifocheck_fbbpl(3)
    );
  tx_fifocheck_fbbpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_3_FFX_RST
    );
  tx_fifocheck_fbbpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_5_FFX_RST,
      O => tx_fifocheck_fbbpl(5)
    );
  tx_fifocheck_fbbpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_5_FFX_RST
    );
  memcontroller_Q3_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(15),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_15_FFX_RST,
      O => q3(15)
    );
  q3_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_15_FFX_RST
    );
  rx_output_fifo_BU390 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1547,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1579_FFX_RST,
      O => rx_output_fifo_N1579
    );
  rx_output_fifo_N1579_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1579_FFX_RST
    );
  rx_output_fifo_BU384 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1550,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1583_FFY_RST,
      O => rx_output_fifo_N1582
    );
  rx_output_fifo_N1583_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1583_FFY_RST
    );
  rx_output_fifo_BU382 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1551,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1583_FFX_RST,
      O => rx_output_fifo_N1583
    );
  rx_output_fifo_N1583_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1583_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(10),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_27_FFY_RST,
      O => mac_control_phystat(26)
    );
  mac_control_phystat_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_27_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(11),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_27_FFX_RST,
      O => mac_control_phystat(27)
    );
  mac_control_phystat_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_27_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(3),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_19_FFX_RST,
      O => mac_control_phystat(19)
    );
  mac_control_phystat_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_19_FFX_RST
    );
  memcontroller_Q3_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(25),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_25_FFX_RST,
      O => q3(25)
    );
  q3_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_25_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(12),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_29_FFY_RST,
      O => mac_control_phystat(28)
    );
  mac_control_phystat_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_29_FFY_RST
    );
  memcontroller_Q3_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(17),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_17_FFX_RST,
      O => q3(17)
    );
  q3_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_17_FFX_RST
    );
  memcontroller_oe_1767 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_wen,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_oe_FFX_RST,
      O => memcontroller_oe
    );
  memcontroller_oe_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_oe_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_sin,
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MDIO_IFF_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(0)
    );
  MDIO_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MDIO_IFF_RST
    );
  rx_output_DOUT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_10_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_10_OFF_RST,
      O => rx_output_DOUT_10_OBUF
    );
  DOUT_10_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_10_OFF_RST
    );
  slowclock_RXCRCERRSR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_rxcrcerrl,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxcrcerrsr_FFY_RST,
      O => rxcrcerrsr
    );
  rxcrcerrsr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxcrcerrsr_FFY_RST
    );
  mac_control_dout_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N74720,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_27_FFY_RST,
      O => mac_control_dout(27)
    );
  mac_control_dout_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_27_FFY_RST
    );
  mac_control_dout_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N74424,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_19_FFY_RST,
      O => mac_control_dout(19)
    );
  mac_control_dout_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_19_FFY_RST
    );
  mac_control_txf_rst_1768 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0062,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_txf_rst_FFY_RST,
      O => mac_control_txf_rst
    );
  mac_control_txf_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_rst_FFY_RST
    );
  memcontroller_Q2_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(23),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_23_FFX_RST,
      O => q2(23)
    );
  q2_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_23_FFX_RST
    );
  memcontroller_Q2_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(15),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_15_FFX_RST,
      O => q2(15)
    );
  q2_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_15_FFX_RST
    );
  rx_output_fifo_BU325 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1569,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1577_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1577
    );
  rx_output_fifo_N1577_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1577_FFX_SET
    );
  mac_control_PHY_status_PHYSTAT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(11),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_11_FFX_RST,
      O => mac_control_phystat(11)
    );
  mac_control_phystat_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_11_FFX_RST
    );
  rx_output_fifo_BU334 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1567,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1575_FFX_RST,
      O => rx_output_fifo_N1575
    );
  rx_output_fifo_N1575_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1575_FFX_RST
    );
  memcontroller_Q2_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(24),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_25_FFY_RST,
      O => q2(24)
    );
  q2_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_25_FFY_RST
    );
  memcontroller_Q2_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(25),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_25_FFX_RST,
      O => q2(25)
    );
  q2_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_25_FFX_RST
    );
  rx_output_fifo_BU370 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N4,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1605_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1604
    );
  rx_output_fifo_N1605_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1605_FFY_SET
    );
  memcontroller_Q2_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(17),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_17_FFX_RST,
      O => q2(17)
    );
  q2_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_17_FFX_RST
    );
  rx_output_fifo_BU372 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1603_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1603
    );
  rx_output_fifo_N1603_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1603_FFX_SET
    );
  rx_output_fifo_BU364 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N7,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1607_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1607
    );
  rx_output_fifo_N1607_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1607_FFX_SET
    );
  mac_control_PHY_status_PHYSTAT_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(9),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_25_FFX_RST,
      O => mac_control_phystat(25)
    );
  mac_control_phystat_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_25_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(1),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_17_FFX_RST,
      O => mac_control_phystat(17)
    );
  mac_control_phystat_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_17_FFX_RST
    );
  memcontroller_Q3_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(31),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_31_FFX_RST,
      O => q3(31)
    );
  q3_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_31_FFX_RST
    );
  memcontroller_Q3_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(23),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_23_FFX_RST,
      O => q3(23)
    );
  q3_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_23_FFX_RST
    );
  rx_output_fifo_BU140 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N10,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1546_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1546
    );
  rx_output_fifo_N1546_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1546_FFX_SET
    );
  rx_output_fifo_BU301 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N2,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1610_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1610
    );
  rx_output_fifo_N1610_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1610_FFX_SET
    );
  rx_output_fifo_BU318 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1547,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1563_FFX_RST,
      O => rx_output_fifo_N1563
    );
  rx_output_fifo_N1563_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1563_FFX_RST
    );
  rx_output_fifo_BU310 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1551,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1567_FFX_RST,
      O => rx_output_fifo_N1567
    );
  rx_output_fifo_N1567_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1567_FFX_RST
    );
  memcontroller_Q2_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(10),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_11_FFY_RST,
      O => q2(10)
    );
  q2_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_11_FFY_RST
    );
  rx_output_fifo_BU167 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1611,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1627_FFX_RST,
      O => rx_output_fifo_N1627
    );
  rx_output_fifo_N1627_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1627_FFX_RST
    );
  memcontroller_Q2_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(11),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_11_FFX_RST,
      O => q2(11)
    );
  q2_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_11_FFX_RST
    );
  rx_output_fifo_BU308 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1552,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1569_FFY_RST,
      O => rx_output_fifo_N1568
    );
  rx_output_fifo_N1569_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1569_FFY_RST
    );
  rx_output_fifo_BU314 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1549,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1565_FFX_RST,
      O => rx_output_fifo_N1565
    );
  rx_output_fifo_N1565_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1565_FFX_RST
    );
  rx_output_fifo_BU306 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1553,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1569_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1569
    );
  rx_output_fifo_N1569_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1569_FFX_SET
    );
  rx_output_fifo_BU161 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1613,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1629_FFX_RST,
      O => rx_output_fifo_N1629
    );
  rx_output_fifo_N1629_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1629_FFX_RST
    );
  rx_output_fifo_BU146 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1617,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1633_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1633
    );
  rx_output_fifo_N1633_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1633_FFX_SET
    );
  memcontroller_Q2_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(21),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_21_FFX_RST,
      O => q2(21)
    );
  q2_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_21_FFX_RST
    );
  memcontroller_Q2_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(13),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_13_FFX_RST,
      O => q2(13)
    );
  q2_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_13_FFX_RST
    );
  rx_output_fifo_BU155 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1615,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1631_FFX_RST,
      O => rx_output_fifo_N1631
    );
  rx_output_fifo_N1631_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1631_FFX_RST
    );
  rx_output_fifo_BU340 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1565,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1573_FFX_RST,
      O => rx_output_fifo_N1573
    );
  rx_output_fifo_N1573_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1573_FFX_RST
    );
  memcontroller_Q2_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(31),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_31_FFX_RST,
      O => q2(31)
    );
  q2_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_31_FFX_RST
    );
  memcontroller_Q2_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(22),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_23_FFY_RST,
      O => q2(22)
    );
  q2_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_23_FFY_RST
    );
  rx_input_memio_addrchk_maceq_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq_2_rt,
      CE => rx_input_memio_addrchk_maceq_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_2_FFX_RST,
      O => rx_input_memio_addrchk_maceq(2)
    );
  rx_input_memio_addrchk_maceq_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_2_FFX_RST
    );
  rx_input_memio_addrchk_maceq_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq_4_rt,
      CE => rx_input_memio_addrchk_maceq_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_4_FFX_RST,
      O => rx_input_memio_addrchk_maceq(4)
    );
  rx_input_memio_addrchk_maceq_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_4_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd2,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_done_FFY_RST,
      O => mac_control_PHY_status_done
    );
  mac_control_PHY_status_done_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_done_FFY_RST
    );
  tx_output_crcl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(24),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_24_FFY_RST,
      O => tx_output_crcl(24)
    );
  tx_output_crcl_24_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_24_FFY_RST
    );
  tx_output_crcl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(16),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_16_FFY_RST,
      O => tx_output_crcl(16)
    );
  tx_output_crcl_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_16_FFY_RST
    );
  mac_control_dout_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N76959,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_6_FFY_RST,
      O => mac_control_dout(6)
    );
  mac_control_dout_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_6_FFY_RST
    );
  rx_input_memio_crcl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(11),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_11_FFY_RST,
      O => rx_input_memio_crcl(11)
    );
  rx_input_memio_crcl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_11_FFY_RST
    );
  tx_output_addrl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(0),
      CE => tx_output_addrl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_1_FFY_RST,
      O => tx_output_addrl(0)
    );
  tx_output_addrl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_1_FFY_RST
    );
  tx_output_addrl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(1),
      CE => tx_output_addrl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_1_FFX_RST,
      O => tx_output_addrl(1)
    );
  tx_output_addrl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_1_FFX_RST
    );
  tx_output_addrl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(3),
      CE => tx_output_addrl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_3_FFX_RST,
      O => tx_output_addrl(3)
    );
  tx_output_addrl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_3_FFX_RST
    );
  tx_output_addrl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(5),
      CE => tx_output_addrl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_5_FFX_RST,
      O => tx_output_addrl(5)
    );
  tx_output_addrl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_5_FFX_RST
    );
  tx_output_addrl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(7),
      CE => tx_output_addrl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_7_FFX_RST,
      O => tx_output_addrl(7)
    );
  tx_output_addrl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_7_FFX_RST
    );
  rx_output_len_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(11),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_11_FFX_RST,
      O => rx_output_len(11)
    );
  rx_output_len_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_11_FFX_RST
    );
  rx_output_mdl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(11),
      CE => rx_output_mdl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_11_FFX_RST,
      O => rx_output_mdl(11)
    );
  rx_output_mdl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_11_FFX_RST
    );
  tx_output_addrl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(8),
      CE => tx_output_addrl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_9_FFY_RST,
      O => tx_output_addrl(8)
    );
  tx_output_addrl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_9_FFY_RST
    );
  rx_output_DOUT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_5_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_5_OFF_RST,
      O => rx_output_DOUT_5_OBUF
    );
  DOUT_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_5_OFF_RST
    );
  rx_output_DOUT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_6_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_6_OFF_RST,
      O => rx_output_DOUT_6_OBUF
    );
  DOUT_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_6_OFF_RST
    );
  rx_output_DOUT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_7_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_7_OFF_RST,
      O => rx_output_DOUT_7_OBUF
    );
  DOUT_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_7_OFF_RST
    );
  rx_output_DOUT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_8_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_8_OFF_RST,
      O => rx_output_DOUT_8_OBUF
    );
  DOUT_8_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_8_OFF_RST
    );
  rx_output_DOUT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_9_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_9_OFF_RST,
      O => rx_output_DOUT_9_OBUF
    );
  DOUT_9_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_9_OFF_RST
    );
  rx_output_len_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(7),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_7_FFX_RST,
      O => rx_output_len(7)
    );
  rx_output_len_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_7_FFX_RST
    );
  rx_output_mdl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(7),
      CE => rx_output_mdl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_7_FFX_RST,
      O => rx_output_mdl(7)
    );
  rx_output_mdl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_7_FFX_RST
    );
  rx_output_len_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(8),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_9_FFY_RST,
      O => rx_output_len(8)
    );
  rx_output_len_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_9_FFY_RST
    );
  rx_output_len_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(9),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_9_FFX_RST,
      O => rx_output_len(9)
    );
  rx_output_len_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_9_FFX_RST
    );
  rx_output_mdl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(9),
      CE => rx_output_mdl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_9_FFX_RST,
      O => rx_output_mdl(9)
    );
  rx_output_mdl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_9_FFX_RST
    );
  rx_input_GMII_ro_1769 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_ro_LOGIC_ONE,
      CE => rx_input_GMII_dvdelta,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_endf,
      O => rx_input_GMII_ro
    );
  tx_output_outselll_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => tx_output_outsell(0),
      CE => tx_output_outselll_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => tx_output_outselll_1_FFY_SET,
      RST => GND,
      O => tx_output_outselll(0)
    );
  tx_output_outselll_1_FFY_SETOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outselll_1_FFY_SET
    );
  tx_output_outselll_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_outsell(1),
      CE => tx_output_outselll_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outselll_1_FFX_RST,
      O => tx_output_outselll(1)
    );
  tx_output_outselll_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outselll_1_FFX_RST
    );
  tx_output_outselll_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_outsell(2),
      CE => tx_output_outselll_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outselll_3_FFY_RST,
      O => tx_output_outselll(2)
    );
  tx_output_outselll_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outselll_3_FFY_RST
    );
  tx_output_outselll_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_outsell(3),
      CE => tx_output_outselll_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outselll_3_FFX_RST,
      O => tx_output_outselll(3)
    );
  tx_output_outselll_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outselll_3_FFX_RST
    );
  tx_output_data_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(0),
      CE => tx_output_data_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_0_FFY_RST,
      O => tx_output_data(0)
    );
  tx_output_data_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_0_FFY_RST
    );
  tx_output_data_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(1),
      CE => tx_output_data_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_1_FFY_RST,
      O => tx_output_data(1)
    );
  tx_output_data_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_1_FFY_RST
    );
  tx_output_crcl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(12),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_12_FFY_RST,
      O => tx_output_crcl(12)
    );
  tx_output_crcl_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_12_FFY_RST
    );
  tx_output_data_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(2),
      CE => tx_output_data_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_2_FFY_RST,
      O => tx_output_data(2)
    );
  tx_output_data_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_2_FFY_RST
    );
  tx_output_data_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(3),
      CE => tx_output_data_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_3_FFY_RST,
      O => tx_output_data(3)
    );
  tx_output_data_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_3_FFY_RST
    );
  mac_control_dout_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N76751,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_2_FFY_RST,
      O => mac_control_dout(2)
    );
  mac_control_dout_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_2_FFY_RST
    );
  tx_output_cs_FFd2_1770 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd3,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd2_FFX_RST,
      O => tx_output_cs_FFd2
    );
  tx_output_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd2_FFX_RST
    );
  tx_output_cs_FFd3_1771 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd7,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd3_FFX_RST,
      O => tx_output_cs_FFd3
    );
  tx_output_cs_FFd3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd3_FFX_RST
    );
  tx_output_cs_FFd9_1772 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd10,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd10_FFY_RST,
      O => tx_output_cs_FFd9
    );
  tx_output_cs_FFd10_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd10_FFY_RST
    );
  tx_output_cs_FFd10_1773 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd11,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd10_FFX_RST,
      O => tx_output_cs_FFd10
    );
  tx_output_cs_FFd10_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd10_FFX_RST
    );
  tx_input_enable_1774 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_enable_LOGIC_ONE,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => tx_input_enable,
      O => tx_input_enable
    );
  rx_input_memio_crcl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(3),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_3_FFY_RST,
      O => rx_input_memio_crcl(3)
    );
  rx_input_memio_crcl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_3_FFY_RST
    );
  tx_fifocheck_FIFOFULL : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfifofull_LOGIC_ONE,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => tx_fifocheck_N73964,
      O => txfifofull
    );
  tx_output_bcntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_39,
      CE => tx_output_bcntl_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_2_FFY_RST,
      O => tx_output_bcntl(1)
    );
  tx_output_bcntl_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_2_FFY_RST
    );
  tx_output_bcntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_40,
      CE => tx_output_bcntl_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_2_FFX_RST,
      O => tx_output_bcntl(2)
    );
  tx_output_bcntl_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_2_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(13),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_29_FFX_RST,
      O => mac_control_phystat(29)
    );
  mac_control_phystat_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_29_FFX_RST
    );
  memcontroller_Q3_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(27),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_27_FFX_RST,
      O => q3(27)
    );
  q3_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_27_FFX_RST
    );
  memcontroller_Q3_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(19),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_19_FFX_RST,
      O => q3(19)
    );
  q3_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_19_FFX_RST
    );
  rx_output_fifo_BU386 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1549,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1581_FFX_RST,
      O => rx_output_fifo_N1581
    );
  rx_output_fifo_N1581_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1581_FFX_RST
    );
  memcontroller_Q3_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(29),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_29_FFX_RST,
      O => q3(29)
    );
  q3_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_29_FFX_RST
    );
  rx_output_ceinll_1775 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_ceinl,
      CE => rx_output_ceinll_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_ceinll_FFY_RST,
      O => rx_output_ceinll
    );
  rx_output_ceinll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_ceinll_FFY_RST
    );
  tx_output_crcl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(10),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_10_FFY_RST,
      O => tx_output_crcl(10)
    );
  tx_output_crcl_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_10_FFY_RST
    );
  memcontroller_dnout_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_28_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_28_OFF_RST,
      O => memcontroller_dnout(28)
    );
  MD_28_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_28_OFF_RST
    );
  memcontroller_ts_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_28_TFF_RST,
      O => memcontroller_ts(28)
    );
  MD_28_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_28_TFF_RST
    );
  memcontroller_qn_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(29),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_29_IFF_RST,
      O => memcontroller_qn(29)
    );
  MD_29_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_29_IFF_RST
    );
  memcontroller_dnout_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_29_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_29_OFF_RST,
      O => memcontroller_dnout(29)
    );
  MD_29_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_29_OFF_RST
    );
  memcontroller_ts_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_29_TFF_RST,
      O => memcontroller_ts(29)
    );
  MD_29_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_29_TFF_RST
    );
  memcontroller_addr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_0_OD,
      CE => MA_0_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_0_OFF_RST,
      O => memcontroller_ADDREXT(0)
    );
  MA_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_0_OFF_RST
    );
  rx_input_GMII_rxdl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_3_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_3_IFF_RST,
      O => rx_input_GMII_rxdl(3)
    );
  RXD_3_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_3_IFF_RST
    );
  rx_input_GMII_rxdl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_4_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_4_IFF_RST,
      O => rx_input_GMII_rxdl(4)
    );
  RXD_4_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_4_IFF_RST
    );
  rx_input_GMII_rxdl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_5_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_5_IFF_RST,
      O => rx_input_GMII_rxdl(5)
    );
  RXD_5_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_5_IFF_RST
    );
  rx_input_GMII_rxdl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_6_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_6_IFF_RST,
      O => rx_input_GMII_rxdl(6)
    );
  RXD_6_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_6_IFF_RST
    );
  rx_input_GMII_rxdl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_7_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_7_IFF_RST,
      O => rx_input_GMII_rxdl(7)
    );
  RXD_7_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_7_IFF_RST
    );
  tx_input_dinl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_10_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_10_IFF_RST,
      O => tx_input_dinl(10)
    );
  DIN_10_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_10_IFF_RST
    );
  tx_input_dinl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_11_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_11_IFF_RST,
      O => tx_input_dinl(11)
    );
  DIN_11_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_11_IFF_RST
    );
  tx_input_dinl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_12_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_12_IFF_RST,
      O => tx_input_dinl(12)
    );
  DIN_12_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_12_IFF_RST
    );
  tx_input_dinl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_13_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_13_IFF_RST,
      O => tx_input_dinl(13)
    );
  DIN_13_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_13_IFF_RST
    );
  tx_input_dinl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_14_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_14_IFF_RST,
      O => tx_input_dinl(14)
    );
  DIN_14_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_14_IFF_RST
    );
  tx_output_data_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(4),
      CE => tx_output_data_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_4_FFY_RST,
      O => tx_output_data(4)
    );
  tx_output_data_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_4_FFY_RST
    );
  tx_output_data_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(5),
      CE => tx_output_data_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_5_FFY_RST,
      O => tx_output_data(5)
    );
  tx_output_data_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_5_FFY_RST
    );
  tx_output_data_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(6),
      CE => tx_output_data_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_6_FFY_RST,
      O => tx_output_data(6)
    );
  tx_output_data_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_6_FFY_RST
    );
  tx_output_data_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(7),
      CE => tx_output_data_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_7_FFY_RST,
      O => tx_output_data(7)
    );
  tx_output_data_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_7_FFY_RST
    );
  rx_output_denll_1776 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_denl,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => rx_output_denll_FFY_RST,
      O => rx_output_denll
    );
  rx_output_denll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_denll_FFY_RST
    );
  rx_output_len_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(0),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_1_FFY_RST,
      O => rx_output_len(0)
    );
  rx_output_len_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_1_FFY_RST
    );
  rx_output_len_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(1),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_1_FFX_RST,
      O => rx_output_len(1)
    );
  rx_output_len_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_1_FFX_RST
    );
  rx_output_mdl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(1),
      CE => rx_output_mdl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_1_FFX_RST,
      O => rx_output_mdl(1)
    );
  rx_output_mdl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_1_FFX_RST
    );
  rx_output_len_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(2),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_3_FFY_RST,
      O => rx_output_len(2)
    );
  rx_output_len_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_3_FFY_RST
    );
  rx_output_len_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(3),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_3_FFX_RST,
      O => rx_output_len(3)
    );
  rx_output_len_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_3_FFX_RST
    );
  rx_output_mdl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(3),
      CE => rx_output_mdl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_3_FFX_RST,
      O => rx_output_mdl(3)
    );
  rx_output_mdl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_3_FFX_RST
    );
  rx_output_len_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(4),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_5_FFY_RST,
      O => rx_output_len(4)
    );
  rx_output_len_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_5_FFY_RST
    );
  rx_output_len_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(5),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_5_FFX_RST,
      O => rx_output_len(5)
    );
  rx_output_len_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_5_FFX_RST
    );
  rx_output_len_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(6),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_7_FFY_RST,
      O => rx_output_len(6)
    );
  rx_output_len_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_7_FFY_RST
    );
  rx_output_mdl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(5),
      CE => rx_output_mdl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_5_FFX_RST,
      O => rx_output_mdl(5)
    );
  rx_output_mdl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_5_FFX_RST
    );
  tx_output_addrl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(9),
      CE => tx_output_addrl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_addrl_9_FFX_RST,
      O => tx_output_addrl(9)
    );
  tx_output_addrl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_addrl_9_FFX_RST
    );
  rx_output_len_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(13),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_13_FFX_RST,
      O => rx_output_len(13)
    );
  rx_output_len_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_13_FFX_RST
    );
  rx_output_mdl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(21),
      CE => rx_output_mdl_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_21_FFX_RST,
      O => rx_output_mdl(21)
    );
  rx_output_mdl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_21_FFX_RST
    );
  rx_output_mdl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(13),
      CE => rx_output_mdl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_13_FFX_RST,
      O => rx_output_mdl(13)
    );
  rx_output_mdl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_13_FFX_RST
    );
  rx_output_len_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(14),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_15_FFY_RST,
      O => rx_output_len(14)
    );
  rx_output_len_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_15_FFY_RST
    );
  rx_output_len_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(15),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_15_FFX_RST,
      O => rx_output_len(15)
    );
  rx_output_len_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_15_FFX_RST
    );
  rx_output_mdl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(31),
      CE => rx_output_mdl_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_31_FFX_RST,
      O => rx_output_mdl(31)
    );
  rx_output_mdl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_31_FFX_RST
    );
  rx_output_mdl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(23),
      CE => rx_output_mdl_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_23_FFX_RST,
      O => rx_output_mdl(23)
    );
  rx_output_mdl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_23_FFX_RST
    );
  rx_output_mdl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(24),
      CE => rx_output_mdl_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_25_FFY_RST,
      O => rx_output_mdl(24)
    );
  rx_output_mdl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_25_FFY_RST
    );
  rx_output_mdl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(15),
      CE => rx_output_mdl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_15_FFX_RST,
      O => rx_output_mdl(15)
    );
  rx_output_mdl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_15_FFX_RST
    );
  rx_output_DOUTEN : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUTEN_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUTEN_OFF_RST,
      O => rx_output_DOUTEN_OBUF
    );
  DOUTEN_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUTEN_OFF_RST
    );
  memcontroller_we : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => MWE_OD,
      CE => MWE_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => MWE_OFF_SET,
      RST => GND,
      O => memcontroller_WEEXT
    );
  MWE_OFF_SETOR : X_BUF
    port map (
      I => GSR,
      O => MWE_OFF_SET
    );
  rx_output_nf_1777 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_NEXTFRAME_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => NEXTFRAME_IFF_RST,
      O => rx_output_nf
    );
  NEXTFRAME_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => NEXTFRAME_IFF_RST
    );
  mac_control_LEDACT : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDACT_OD,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => LEDACT_OFF_RST,
      O => mac_control_LEDACT_OBUF
    );
  LEDACT_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDACT_OFF_RST
    );
  tx_output_TXD_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_0_OD,
      CE => TXD_0_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_0_OFF_RST,
      O => tx_output_TXD_0_OBUF
    );
  TXD_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_0_OFF_RST
    );
  tx_output_bcntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_42,
      CE => tx_output_bcntl_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_4_FFX_RST,
      O => tx_output_bcntl(4)
    );
  tx_output_bcntl_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_4_FFX_RST
    );
  tx_output_bcntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_44,
      CE => tx_output_bcntl_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_6_FFX_RST,
      O => tx_output_bcntl(6)
    );
  tx_output_bcntl_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_6_FFX_RST
    );
  rx_output_bpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(1),
      CE => rx_output_bpl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_1_FFX_RST,
      O => rx_output_bpl(1)
    );
  rx_output_bpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_1_FFX_RST
    );
  tx_output_bcntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_46,
      CE => tx_output_bcntl_8_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_8_FFX_RST,
      O => tx_output_bcntl(8)
    );
  tx_output_bcntl_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_8_FFX_RST
    );
  rx_output_bpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(3),
      CE => rx_output_bpl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bpl_3_FFX_RST,
      O => rx_output_bpl(3)
    );
  rx_output_bpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bpl_3_FFX_RST
    );
  tx_output_datal_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(1),
      CE => tx_output_datal_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_1_FFX_RST,
      O => tx_output_datal(1)
    );
  tx_output_datal_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_1_FFX_RST
    );
  tx_output_bcntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_48,
      CE => tx_output_bcntl_10_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_10_FFX_RST,
      O => tx_output_bcntl(10)
    );
  tx_output_bcntl_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_10_FFX_RST
    );
  mac_control_LED100 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LED100_OD,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => LED100_OFF_RST,
      O => mac_control_LED100_OBUF
    );
  LED100_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LED100_OFF_RST
    );
  tx_input_newframel_1778 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_NEWFRAME_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => NEWFRAME_IFF_RST,
      O => tx_input_newframel
    );
  NEWFRAME_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => NEWFRAME_IFF_RST
    );
  mac_control_LED1000 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LED1000_OD,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => LED1000_OFF_RST,
      O => mac_control_LED1000_OBUF
    );
  LED1000_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LED1000_OFF_RST
    );
  tx_output_TXEN_1779 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TX_EN_OD,
      CE => TX_EN_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TX_EN_OFF_RST,
      O => tx_output_TXEN
    );
  TX_EN_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TX_EN_OFF_RST
    );
  memcontroller_dnout_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_13_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_13_OFF_RST,
      O => memcontroller_dnout(13)
    );
  MD_13_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_13_OFF_RST
    );
  memcontroller_ts_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_13_TFF_RST,
      O => memcontroller_ts(13)
    );
  MD_13_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_13_TFF_RST
    );
  memcontroller_qn_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(22),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_22_IFF_RST,
      O => memcontroller_qn(22)
    );
  MD_22_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_22_IFF_RST
    );
  memcontroller_dnout_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_22_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_22_OFF_RST,
      O => memcontroller_dnout(22)
    );
  MD_22_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_22_OFF_RST
    );
  memcontroller_ts_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_22_TFF_RST,
      O => memcontroller_ts(22)
    );
  MD_22_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_22_TFF_RST
    );
  memcontroller_qn_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_14_IFF_RST,
      O => memcontroller_qn(14)
    );
  MD_14_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_14_IFF_RST
    );
  memcontroller_qn_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(30),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_30_IFF_RST,
      O => memcontroller_qn(30)
    );
  MD_30_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_30_IFF_RST
    );
  memcontroller_dnout_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_14_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_14_OFF_RST,
      O => memcontroller_dnout(14)
    );
  MD_14_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_14_OFF_RST
    );
  memcontroller_ts_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_14_TFF_RST,
      O => memcontroller_ts(14)
    );
  MD_14_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_14_TFF_RST
    );
  rx_output_DOUT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_11_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_11_OFF_RST,
      O => rx_output_DOUT_11_OBUF
    );
  DOUT_11_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_11_OFF_RST
    );
  rx_output_DOUT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_12_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_12_OFF_RST,
      O => rx_output_DOUT_12_OBUF
    );
  DOUT_12_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_12_OFF_RST
    );
  rx_output_DOUT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_13_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_13_OFF_RST,
      O => rx_output_DOUT_13_OBUF
    );
  DOUT_13_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_13_OFF_RST
    );
  rx_output_DOUT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_14_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_14_OFF_RST,
      O => rx_output_DOUT_14_OBUF
    );
  DOUT_14_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_14_OFF_RST
    );
  rx_output_DOUT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_15_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_15_OFF_RST,
      O => rx_output_DOUT_15_OBUF
    );
  DOUT_15_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_15_OFF_RST
    );
  tx_input_dinl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_15_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_15_IFF_RST,
      O => tx_input_dinl(15)
    );
  DIN_15_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_15_IFF_RST
    );
  rx_output_DOUT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_0_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_0_OFF_RST,
      O => rx_output_DOUT_0_OBUF
    );
  DOUT_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_0_OFF_RST
    );
  rx_output_DOUT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_1_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_1_OFF_RST,
      O => rx_output_DOUT_1_OBUF
    );
  DOUT_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_1_OFF_RST
    );
  rx_output_DOUT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_2_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_2_OFF_RST,
      O => rx_output_DOUT_2_OBUF
    );
  DOUT_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_2_OFF_RST
    );
  rx_output_DOUT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_3_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_3_OFF_RST,
      O => rx_output_DOUT_3_OBUF
    );
  DOUT_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_3_OFF_RST
    );
  rx_output_DOUT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_4_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_4_OFF_RST,
      O => rx_output_DOUT_4_OBUF
    );
  DOUT_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_4_OFF_RST
    );
  memcontroller_addr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_15_OD,
      CE => MA_15_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_15_OFF_RST,
      O => memcontroller_ADDREXT(15)
    );
  MA_15_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_15_OFF_RST
    );
  memcontroller_addr_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_16_OD,
      CE => MA_16_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_16_OFF_RST,
      O => memcontroller_ADDREXT(16)
    );
  MA_16_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_16_OFF_RST
    );
  memcontroller_qn_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_10_IFF_RST,
      O => memcontroller_qn(10)
    );
  MD_10_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_10_IFF_RST
    );
  memcontroller_dnout_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_10_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_10_OFF_RST,
      O => memcontroller_dnout(10)
    );
  MD_10_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_10_OFF_RST
    );
  memcontroller_ts_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_10_TFF_RST,
      O => memcontroller_ts(10)
    );
  MD_10_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_10_TFF_RST
    );
  memcontroller_qn_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_11_IFF_RST,
      O => memcontroller_qn(11)
    );
  MD_11_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_11_IFF_RST
    );
  memcontroller_qn_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(20),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_20_IFF_RST,
      O => memcontroller_qn(20)
    );
  MD_20_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_20_IFF_RST
    );
  memcontroller_dnout_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_11_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_11_OFF_RST,
      O => memcontroller_dnout(11)
    );
  MD_11_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_11_OFF_RST
    );
  memcontroller_ts_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_11_TFF_RST,
      O => memcontroller_ts(11)
    );
  MD_11_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_11_TFF_RST
    );
  tx_output_TXD_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_1_OD,
      CE => TXD_1_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_1_OFF_RST,
      O => tx_output_TXD_1_OBUF
    );
  TXD_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_1_OFF_RST
    );
  tx_output_TXD_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_2_OD,
      CE => TXD_2_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_2_OFF_RST,
      O => tx_output_TXD_2_OBUF
    );
  TXD_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_2_OFF_RST
    );
  tx_output_TXD_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_3_OD,
      CE => TXD_3_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_3_OFF_RST,
      O => tx_output_TXD_3_OBUF
    );
  TXD_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_3_OFF_RST
    );
  tx_output_TXD_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_4_OD,
      CE => TXD_4_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_4_OFF_RST,
      O => tx_output_TXD_4_OBUF
    );
  TXD_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_4_OFF_RST
    );
  tx_output_TXD_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_5_OD,
      CE => TXD_5_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_5_OFF_RST,
      O => tx_output_TXD_5_OBUF
    );
  TXD_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_5_OFF_RST
    );
  tx_output_TXD_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_6_OD,
      CE => TXD_6_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_6_OFF_RST,
      O => tx_output_TXD_6_OBUF
    );
  TXD_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_6_OFF_RST
    );
  tx_output_TXD_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_7_OD,
      CE => TXD_7_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_7_OFF_RST,
      O => tx_output_TXD_7_OBUF
    );
  TXD_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_7_OFF_RST
    );
  mac_control_LEDDPX : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDDPX_OD,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => LEDDPX_OFF_RST,
      O => mac_control_LEDDPX_OBUF
    );
  LEDDPX_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDDPX_OFF_RST
    );
  rx_input_GMII_rxdl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_0_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_0_IFF_RST,
      O => rx_input_GMII_rxdl(0)
    );
  RXD_0_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_0_IFF_RST
    );
  rx_input_GMII_rxdl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_1_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_1_IFF_RST,
      O => rx_input_GMII_rxdl(1)
    );
  RXD_1_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_1_IFF_RST
    );
  rx_input_GMII_rxdl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_2_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_2_IFF_RST,
      O => rx_input_GMII_rxdl(2)
    );
  RXD_2_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_2_IFF_RST
    );
  memcontroller_addr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_11_OD,
      CE => MA_11_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_11_OFF_RST,
      O => memcontroller_ADDREXT(11)
    );
  MA_11_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_11_OFF_RST
    );
  memcontroller_addr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_12_OD,
      CE => MA_12_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_12_OFF_RST,
      O => memcontroller_ADDREXT(12)
    );
  MA_12_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_12_OFF_RST
    );
  memcontroller_addr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_13_OD,
      CE => MA_13_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_13_OFF_RST,
      O => memcontroller_ADDREXT(13)
    );
  MA_13_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_13_OFF_RST
    );
  memcontroller_addr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_14_OD,
      CE => MA_14_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_14_OFF_RST,
      O => memcontroller_ADDREXT(14)
    );
  MA_14_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_14_OFF_RST
    );
  memcontroller_addr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_5_OD,
      CE => MA_5_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_5_OFF_RST,
      O => memcontroller_ADDREXT(5)
    );
  MA_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_5_OFF_RST
    );
  memcontroller_addr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_6_OD,
      CE => MA_6_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_6_OFF_RST,
      O => memcontroller_ADDREXT(6)
    );
  MA_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_6_OFF_RST
    );
  memcontroller_addr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_7_OD,
      CE => MA_7_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_7_OFF_RST,
      O => memcontroller_ADDREXT(7)
    );
  MA_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_7_OFF_RST
    );
  memcontroller_addr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_8_OD,
      CE => MA_8_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_8_OFF_RST,
      O => memcontroller_ADDREXT(8)
    );
  MA_8_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_8_OFF_RST
    );
  memcontroller_addr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_9_OD,
      CE => MA_9_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_9_OFF_RST,
      O => memcontroller_ADDREXT(9)
    );
  MA_9_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_9_OFF_RST
    );
  mac_control_PHYRESET : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => PHYRESET_OD,
      CE => mac_control_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => PHYRESET_OFF_RST,
      O => mac_control_PHYRESET_OBUF
    );
  PHYRESET_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => PHYRESET_OFF_RST
    );
  memcontroller_dnl1_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(3),
      CE => memcontroller_dnl1_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_3_FFX_RST,
      O => memcontroller_dnl1(3)
    );
  memcontroller_dnl1_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_3_FFX_RST
    );
  memcontroller_dnl1_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(4),
      CE => memcontroller_dnl1_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_4_FFX_RST,
      O => memcontroller_dnl1(4)
    );
  memcontroller_dnl1_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_4_FFX_RST
    );
  memcontroller_qn_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_0_IFF_RST,
      O => memcontroller_qn(0)
    );
  MD_0_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_0_IFF_RST
    );
  memcontroller_dnout_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_0_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_0_OFF_RST,
      O => memcontroller_dnout(0)
    );
  MD_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_0_OFF_RST
    );
  memcontroller_ts_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_0_TFF_RST,
      O => memcontroller_ts(0)
    );
  MD_0_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_0_TFF_RST
    );
  memcontroller_qn_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_1_IFF_RST,
      O => memcontroller_qn(1)
    );
  MD_1_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_1_IFF_RST
    );
  memcontroller_dnout_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_1_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_1_OFF_RST,
      O => memcontroller_dnout(1)
    );
  MD_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_1_OFF_RST
    );
  memcontroller_ts_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_1_TFF_RST,
      O => memcontroller_ts(1)
    );
  MD_1_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_1_TFF_RST
    );
  memcontroller_qn_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_2_IFF_RST,
      O => memcontroller_qn(2)
    );
  MD_2_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_2_IFF_RST
    );
  memcontroller_qn_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_3_IFF_RST,
      O => memcontroller_qn(3)
    );
  MD_3_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_3_IFF_RST
    );
  memcontroller_dnout_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_2_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_2_OFF_RST,
      O => memcontroller_dnout(2)
    );
  MD_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_2_OFF_RST
    );
  memcontroller_ts_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_2_TFF_RST,
      O => memcontroller_ts(2)
    );
  MD_2_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_2_TFF_RST
    );
  memcontroller_dnout_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_3_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_3_OFF_RST,
      O => memcontroller_dnout(3)
    );
  MD_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_3_OFF_RST
    );
  memcontroller_ts_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_3_TFF_RST,
      O => memcontroller_ts(3)
    );
  MD_3_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_3_TFF_RST
    );
  memcontroller_qn_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_4_IFF_RST,
      O => memcontroller_qn(4)
    );
  MD_4_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_4_IFF_RST
    );
  memcontroller_dnout_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_4_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_4_OFF_RST,
      O => memcontroller_dnout(4)
    );
  MD_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_4_OFF_RST
    );
  memcontroller_ts_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_4_TFF_RST,
      O => memcontroller_ts(4)
    );
  MD_4_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_4_TFF_RST
    );
  memcontroller_qn_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_5_IFF_RST,
      O => memcontroller_qn(5)
    );
  MD_5_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_5_IFF_RST
    );
  memcontroller_qn_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_6_IFF_RST,
      O => memcontroller_qn(6)
    );
  MD_6_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_6_IFF_RST
    );
  memcontroller_dnout_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_20_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_20_OFF_RST,
      O => memcontroller_dnout(20)
    );
  MD_20_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_20_OFF_RST
    );
  memcontroller_ts_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_20_TFF_RST,
      O => memcontroller_ts(20)
    );
  MD_20_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_20_TFF_RST
    );
  memcontroller_qn_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_12_IFF_RST,
      O => memcontroller_qn(12)
    );
  MD_12_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_12_IFF_RST
    );
  memcontroller_dnout_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_12_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_12_OFF_RST,
      O => memcontroller_dnout(12)
    );
  MD_12_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_12_OFF_RST
    );
  memcontroller_ts_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_12_TFF_RST,
      O => memcontroller_ts(12)
    );
  MD_12_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_12_TFF_RST
    );
  memcontroller_qn_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(21),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_21_IFF_RST,
      O => memcontroller_qn(21)
    );
  MD_21_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_21_IFF_RST
    );
  memcontroller_qn_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_13_IFF_RST,
      O => memcontroller_qn(13)
    );
  MD_13_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_13_IFF_RST
    );
  memcontroller_dnout_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_21_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_21_OFF_RST,
      O => memcontroller_dnout(21)
    );
  MD_21_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_21_OFF_RST
    );
  memcontroller_ts_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_21_TFF_RST,
      O => memcontroller_ts(21)
    );
  MD_21_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_21_TFF_RST
    );
  memcontroller_addr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_1_OD,
      CE => MA_1_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_1_OFF_RST,
      O => memcontroller_ADDREXT(1)
    );
  MA_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_1_OFF_RST
    );
  memcontroller_addr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_2_OD,
      CE => MA_2_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_2_OFF_RST,
      O => memcontroller_ADDREXT(2)
    );
  MA_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_2_OFF_RST
    );
  memcontroller_addr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_3_OD,
      CE => MA_3_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_3_OFF_RST,
      O => memcontroller_ADDREXT(3)
    );
  MA_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_3_OFF_RST
    );
  memcontroller_addr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_4_OD,
      CE => MA_4_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_4_OFF_RST,
      O => memcontroller_ADDREXT(4)
    );
  MA_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_4_OFF_RST
    );
  mac_control_dout_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N75420,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_28_FFY_RST,
      O => mac_control_dout(28)
    );
  mac_control_dout_28_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_28_FFY_RST
    );
  mac_control_dout_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N75654,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_29_FFY_RST,
      O => mac_control_dout(29)
    );
  mac_control_dout_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_29_FFY_RST
    );
  memcontroller_dnl2_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(31),
      CE => memcontroller_dnl2_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_31_FFX_RST,
      O => memcontroller_dnl2(31)
    );
  memcontroller_dnl2_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_31_FFX_RST
    );
  memcontroller_dnl2_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(23),
      CE => memcontroller_dnl2_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_23_FFX_RST,
      O => memcontroller_dnl2(23)
    );
  memcontroller_dnl2_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_23_FFX_RST
    );
  memcontroller_dnl2_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(14),
      CE => memcontroller_dnl2_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_15_FFY_RST,
      O => memcontroller_dnl2(14)
    );
  memcontroller_dnl2_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_15_FFY_RST
    );
  memcontroller_dnl2_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(15),
      CE => memcontroller_dnl2_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_15_FFX_RST,
      O => memcontroller_dnl2(15)
    );
  memcontroller_dnl2_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_15_FFX_RST
    );
  memcontroller_dnl2_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(24),
      CE => memcontroller_dnl2_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_25_FFY_RST,
      O => memcontroller_dnl2(24)
    );
  memcontroller_dnl2_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_25_FFY_RST
    );
  memcontroller_dnl2_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(25),
      CE => memcontroller_dnl2_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_25_FFX_RST,
      O => memcontroller_dnl2(25)
    );
  memcontroller_dnl2_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_25_FFX_RST
    );
  memcontroller_dnl2_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(16),
      CE => memcontroller_dnl2_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_17_FFY_RST,
      O => memcontroller_dnl2(16)
    );
  memcontroller_dnl2_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_17_FFY_RST
    );
  memcontroller_dnl2_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(17),
      CE => memcontroller_dnl2_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_17_FFX_RST,
      O => memcontroller_dnl2(17)
    );
  memcontroller_dnl2_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_17_FFX_RST
    );
  memcontroller_dnl2_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(26),
      CE => memcontroller_dnl2_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_27_FFY_RST,
      O => memcontroller_dnl2(26)
    );
  memcontroller_dnl2_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_27_FFY_RST
    );
  memcontroller_dnl2_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(27),
      CE => memcontroller_dnl2_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_27_FFX_RST,
      O => memcontroller_dnl2(27)
    );
  memcontroller_dnl2_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_27_FFX_RST
    );
  memcontroller_dnl2_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(18),
      CE => memcontroller_dnl2_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_19_FFY_RST,
      O => memcontroller_dnl2(18)
    );
  memcontroller_dnl2_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_19_FFY_RST
    );
  memcontroller_dnl2_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(19),
      CE => memcontroller_dnl2_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_19_FFX_RST,
      O => memcontroller_dnl2(19)
    );
  memcontroller_dnl2_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_19_FFX_RST
    );
  memcontroller_dnl2_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(28),
      CE => memcontroller_dnl2_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_29_FFY_RST,
      O => memcontroller_dnl2(28)
    );
  memcontroller_dnl2_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_29_FFY_RST
    );
  rx_input_memio_datal_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_datal_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_1_FFY_RST,
      O => rx_input_memio_datal(0)
    );
  rx_input_memio_datal_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_1_FFY_RST
    );
  memcontroller_dnl2_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(0),
      CE => memcontroller_dnl2_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_1_FFY_RST,
      O => memcontroller_dnl2(0)
    );
  memcontroller_dnl2_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_1_FFY_RST
    );
  slowclock_RXPHYERRSR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_rxphyerrl,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxphyerrsr_FFY_RST,
      O => rxphyerrsr
    );
  rxphyerrsr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxphyerrsr_FFY_RST
    );
  memcontroller_dnl2_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(1),
      CE => memcontroller_dnl2_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_1_FFX_RST,
      O => memcontroller_dnl2(1)
    );
  memcontroller_dnl2_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_1_FFX_RST
    );
  memcontroller_dnl2_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(2),
      CE => memcontroller_dnl2_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_3_FFY_RST,
      O => memcontroller_dnl2(2)
    );
  memcontroller_dnl2_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_3_FFY_RST
    );
  memcontroller_dnl2_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(3),
      CE => memcontroller_dnl2_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_3_FFX_RST,
      O => memcontroller_dnl2(3)
    );
  memcontroller_dnl2_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_3_FFX_RST
    );
  memcontroller_dnl2_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(4),
      CE => memcontroller_dnl2_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_5_FFY_RST,
      O => memcontroller_dnl2(4)
    );
  memcontroller_dnl2_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_5_FFY_RST
    );
  memcontroller_dnl2_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(5),
      CE => memcontroller_dnl2_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_5_FFX_RST,
      O => memcontroller_dnl2(5)
    );
  memcontroller_dnl2_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_5_FFX_RST
    );
  memcontroller_dnl2_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(6),
      CE => memcontroller_dnl2_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_7_FFY_RST,
      O => memcontroller_dnl2(6)
    );
  memcontroller_dnl2_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_7_FFY_RST
    );
  memcontroller_dnl2_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(7),
      CE => memcontroller_dnl2_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_7_FFX_RST,
      O => memcontroller_dnl2(7)
    );
  memcontroller_dnl2_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_7_FFX_RST
    );
  memcontroller_dnl2_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(8),
      CE => memcontroller_dnl2_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_9_FFY_RST,
      O => memcontroller_dnl2(8)
    );
  memcontroller_dnl2_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_9_FFY_RST
    );
  mac_control_sclkdeltal_1780 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_sclkdelta,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_sclkdeltal_FFY_RST,
      O => mac_control_sclkdeltal
    );
  mac_control_sclkdeltal_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_sclkdeltal_FFY_RST
    );
  mac_control_rxcrcerr_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_lut2_16,
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(0)
    );
  mac_control_rxcrcerr_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(2),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(2)
    );
  mac_control_rxcrcerr_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(4),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(4)
    );
  mac_control_rxcrcerr_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(7),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(7)
    );
  mac_control_rxcrcerr_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(11),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(11)
    );
  mac_control_rxcrcerr_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(6),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(6)
    );
  mac_control_rxcrcerr_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(9),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(9)
    );
  tx_output_addr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(14),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_14_FFX_RST,
      O => addr2ext(14)
    );
  addr2ext_14_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => addr2ext_14_FFX_RST
    );
  rx_input_memio_bcnt_88_1781 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_237,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_87_FFY_RST,
      O => rx_input_memio_bcnt_88
    );
  rx_input_memio_bcnt_87_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_87_FFY_RST
    );
  rx_input_memio_bcnt_87_1782 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_236,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_87_FFX_RST,
      O => rx_input_memio_bcnt_87
    );
  rx_input_memio_bcnt_87_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_87_FFX_RST
    );
  rx_input_memio_bcnt_90_1783 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_239,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_89_FFY_RST,
      O => rx_input_memio_bcnt_90
    );
  rx_input_memio_bcnt_89_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_89_FFY_RST
    );
  rx_input_memio_bcnt_92_1784 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_241,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_91_FFY_RST,
      O => rx_input_memio_bcnt_92
    );
  rx_input_memio_bcnt_91_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_91_FFY_RST
    );
  mac_control_rxcrcerr_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(14),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(14)
    );
  mac_control_rxcrcerr_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(16),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(16)
    );
  mac_control_rxcrcerr_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(19),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(19)
    );
  mac_control_rxcrcerr_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(23),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(23)
    );
  mac_control_rxcrcerr_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(18),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(18)
    );
  mac_control_rxcrcerr_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(21),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(21)
    );
  memcontroller_dnl1_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(2),
      CE => memcontroller_dnl1_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_2_FFX_RST,
      O => memcontroller_dnl1(2)
    );
  memcontroller_dnl1_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_2_FFX_RST
    );
  memcontroller_dnl1_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(10),
      CE => memcontroller_dnl1_10_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_10_FFX_RST,
      O => memcontroller_dnl1(10)
    );
  memcontroller_dnl1_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_10_FFX_RST
    );
  memcontroller_dnl1_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(18),
      CE => memcontroller_dnl1_18_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_18_FFX_RST,
      O => memcontroller_dnl1(18)
    );
  memcontroller_dnl1_18_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_18_FFX_RST
    );
  memcontroller_dnl1_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(26),
      CE => memcontroller_dnl1_26_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_26_FFX_RST,
      O => memcontroller_dnl1(26)
    );
  memcontroller_dnl1_26_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_26_FFX_RST
    );
  memcontroller_dnl1_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(11),
      CE => memcontroller_dnl1_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_11_FFX_RST,
      O => memcontroller_dnl1(11)
    );
  memcontroller_dnl1_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_11_FFX_RST
    );
  memcontroller_dnl1_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(24),
      CE => memcontroller_dnl1_24_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_24_FFX_RST,
      O => memcontroller_dnl1(24)
    );
  memcontroller_dnl1_24_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_24_FFX_RST
    );
  memcontroller_dnl1_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(1),
      CE => memcontroller_dnl1_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_1_FFX_RST,
      O => memcontroller_dnl1(1)
    );
  memcontroller_dnl1_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_1_FFX_RST
    );
  memcontroller_dnl1_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(9),
      CE => memcontroller_dnl1_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_9_FFX_RST,
      O => memcontroller_dnl1(9)
    );
  memcontroller_dnl1_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_9_FFX_RST
    );
  memcontroller_dnl1_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(17),
      CE => memcontroller_dnl1_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_17_FFX_RST,
      O => memcontroller_dnl1(17)
    );
  memcontroller_dnl1_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_17_FFX_RST
    );
  memcontroller_dnl1_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(25),
      CE => memcontroller_dnl1_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_25_FFX_RST,
      O => memcontroller_dnl1(25)
    );
  memcontroller_dnl1_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_25_FFX_RST
    );
  rx_input_memio_bcnt_89_1785 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_238,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_89_FFX_RST,
      O => rx_input_memio_bcnt_89
    );
  rx_input_memio_bcnt_89_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_89_FFX_RST
    );
  rx_input_memio_bcnt_91_1786 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_240,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_91_FFX_RST,
      O => rx_input_memio_bcnt_91
    );
  rx_input_memio_bcnt_91_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_91_FFX_RST
    );
  rx_input_memio_bcnt_94_1787 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_243,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_93_FFY_RST,
      O => rx_input_memio_bcnt_94
    );
  rx_input_memio_bcnt_93_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_93_FFY_RST
    );
  rx_input_memio_bcnt_93_1788 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_242,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_93_FFX_RST,
      O => rx_input_memio_bcnt_93
    );
  rx_input_memio_bcnt_93_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_93_FFX_RST
    );
  rx_input_memio_bcnt_96_1789 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_245,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_95_FFY_RST,
      O => rx_input_memio_bcnt_96
    );
  rx_input_memio_bcnt_95_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_95_FFY_RST
    );
  rx_input_memio_bcnt_98_1790 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_247,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_97_FFY_RST,
      O => rx_input_memio_bcnt_98
    );
  rx_input_memio_bcnt_97_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_97_FFY_RST
    );
  memcontroller_dnl1_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(21),
      CE => memcontroller_dnl1_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_21_FFX_RST,
      O => memcontroller_dnl1(21)
    );
  memcontroller_dnl1_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_21_FFX_RST
    );
  memcontroller_dnl1_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(29),
      CE => memcontroller_dnl1_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_29_FFX_RST,
      O => memcontroller_dnl1(29)
    );
  memcontroller_dnl1_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_29_FFX_RST
    );
  memcontroller_dnl1_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(22),
      CE => memcontroller_dnl1_22_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_22_FFX_RST,
      O => memcontroller_dnl1(22)
    );
  memcontroller_dnl1_22_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_22_FFX_RST
    );
  memcontroller_dnl1_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(30),
      CE => memcontroller_dnl1_30_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_30_FFX_RST,
      O => memcontroller_dnl1(30)
    );
  memcontroller_dnl1_30_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_30_FFX_RST
    );
  memcontroller_dnl1_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(31),
      CE => memcontroller_dnl1_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_31_FFX_RST,
      O => memcontroller_dnl1(31)
    );
  memcontroller_dnl1_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_31_FFX_RST
    );
  rx_input_memio_bp_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(0),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_0_FFX_RST,
      O => rx_input_memio_bp(0)
    );
  rx_input_memio_bp_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_0_FFX_RST
    );
  rx_input_memio_bp_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(2),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_2_FFX_RST,
      O => rx_input_memio_bp(2)
    );
  rx_input_memio_bp_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_2_FFX_RST
    );
  rx_input_memio_bp_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(4),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_4_FFX_RST,
      O => rx_input_memio_bp(4)
    );
  rx_input_memio_bp_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_4_FFX_RST
    );
  memcontroller_dnl1_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(19),
      CE => memcontroller_dnl1_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_19_FFX_RST,
      O => memcontroller_dnl1(19)
    );
  memcontroller_dnl1_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_19_FFX_RST
    );
  memcontroller_dnl1_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(27),
      CE => memcontroller_dnl1_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_27_FFX_RST,
      O => memcontroller_dnl1(27)
    );
  memcontroller_dnl1_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_27_FFX_RST
    );
  memcontroller_dnl1_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(12),
      CE => memcontroller_dnl1_12_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_12_FFX_RST,
      O => memcontroller_dnl1(12)
    );
  memcontroller_dnl1_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_12_FFX_RST
    );
  memcontroller_dnl1_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(20),
      CE => memcontroller_dnl1_20_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_20_FFX_RST,
      O => memcontroller_dnl1(20)
    );
  memcontroller_dnl1_20_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_20_FFX_RST
    );
  memcontroller_dnl1_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(28),
      CE => memcontroller_dnl1_28_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_28_FFX_RST,
      O => memcontroller_dnl1(28)
    );
  memcontroller_dnl1_28_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_28_FFX_RST
    );
  mac_control_rxoferr_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(6),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(6)
    );
  mac_control_rxoferr_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(8),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(8)
    );
  mac_control_rxoferr_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(15),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(15)
    );
  mac_control_rxoferr_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(10),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(10)
    );
  mac_control_rxoferr_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(13),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(13)
    );
  mac_control_rxoferr_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(17),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(17)
    );
  mac_control_rxcrcerr_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(26),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(26)
    );
  mac_control_rxcrcerr_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(28),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(28)
    );
  mac_control_rxcrcerr_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(31),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(31)
    );
  mac_control_rxcrcerr_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(30),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(30)
    );
  rx_input_memio_bp_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(1),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_0_FFY_RST,
      O => rx_input_memio_bp(1)
    );
  rx_input_memio_bp_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_0_FFY_RST
    );
  mac_control_rxoferr_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_lut2_16,
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(0)
    );
  mac_control_rxoferr_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(5),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(5)
    );
  mac_control_rxoferr_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(2),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(2)
    );
  mac_control_rxoferr_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(9),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(9)
    );
  mac_control_rxoferr_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(4),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(4)
    );
  mac_control_rxoferr_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(7),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(7)
    );
  mac_control_rxoferr_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(11),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(11)
    );
  mac_control_rxphyerr_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(22),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(22)
    );
  mac_control_rxphyerr_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(24),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(24)
    );
  mac_control_rxphyerr_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(27),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(27)
    );
  mac_control_rxphyerr_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(31),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(31)
    );
  mac_control_rxphyerr_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(26),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(26)
    );
  mac_control_rxphyerr_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(29),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(29)
    );
  mac_control_rxcrcerr_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(20),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(20)
    );
  mac_control_rxcrcerr_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(22),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(22)
    );
  mac_control_rxcrcerr_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(25),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(25)
    );
  mac_control_rxcrcerr_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(29),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(29)
    );
  mac_control_rxcrcerr_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(24),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(24)
    );
  mac_control_rxcrcerr_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(27),
      CE => mac_control_n0055,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0054,
      O => mac_control_rxcrcerr_cnt(27)
    );
  rx_input_memio_bp_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(10),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_10_FFX_RST,
      O => rx_input_memio_bp(10)
    );
  rx_input_memio_bp_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_10_FFX_RST
    );
  rx_input_memio_bp_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(12),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_12_FFX_RST,
      O => rx_input_memio_bp(12)
    );
  rx_input_memio_bp_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_12_FFX_RST
    );
  rx_input_memio_bp_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(15),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_14_FFY_RST,
      O => rx_input_memio_bp(15)
    );
  rx_input_memio_bp_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_14_FFY_RST
    );
  rx_input_memio_bp_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(14),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_14_FFX_RST,
      O => rx_input_memio_bp(14)
    );
  rx_input_memio_bp_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_14_FFX_RST
    );
  mac_control_rxoferr_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(1),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(1)
    );
  mac_control_rxoferr_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(3),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(3)
    );
  mac_control_rxphyerr_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(4),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(4)
    );
  mac_control_rxphyerr_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(6),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(6)
    );
  mac_control_rxphyerr_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(9),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(9)
    );
  mac_control_rxphyerr_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(13),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(13)
    );
  mac_control_rxphyerr_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(8),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(8)
    );
  mac_control_rxphyerr_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(11),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(11)
    );
  mac_control_ledrx_cnt_159_1791 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_306,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_159_FFX_RST,
      O => mac_control_ledrx_cnt_159
    );
  mac_control_ledrx_cnt_159_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_159_FFX_RST
    );
  mac_control_ledrx_cnt_162_1792 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_309,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_161_FFY_RST,
      O => mac_control_ledrx_cnt_162
    );
  mac_control_ledrx_cnt_161_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_161_FFY_RST
    );
  mac_control_ledrx_cnt_161_1793 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_308,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_161_FFX_RST,
      O => mac_control_ledrx_cnt_161
    );
  mac_control_ledrx_cnt_161_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_161_FFX_RST
    );
  mac_control_ledrx_cnt_164_1794 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_311,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_163_FFY_RST,
      O => mac_control_ledrx_cnt_164
    );
  mac_control_ledrx_cnt_163_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_163_FFY_RST
    );
  mac_control_ledrx_cnt_165_1795 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_312,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_165_FFX_RST,
      O => mac_control_ledrx_cnt_165
    );
  mac_control_ledrx_cnt_165_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_165_FFX_RST
    );
  rx_input_memio_bp_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(6),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_6_FFX_RST,
      O => rx_input_memio_bp(6)
    );
  rx_input_memio_bp_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_6_FFX_RST
    );
  rx_input_memio_bp_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(13),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_12_FFY_RST,
      O => rx_input_memio_bp(13)
    );
  rx_input_memio_bp_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_12_FFY_RST
    );
  rx_input_memio_bp_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(8),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_8_FFX_RST,
      O => rx_input_memio_bp(8)
    );
  rx_input_memio_bp_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_8_FFX_RST
    );
  mac_control_rxoferr_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(24),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(24)
    );
  mac_control_rxoferr_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(26),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(26)
    );
  mac_control_ledrx_cnt_154_1796 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_301,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_154_FFY_RST,
      O => mac_control_ledrx_cnt_154
    );
  mac_control_ledrx_cnt_154_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_154_FFY_RST
    );
  mac_control_rxoferr_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(28),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(28)
    );
  mac_control_rxoferr_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(31),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(31)
    );
  mac_control_rxoferr_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(30),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(30)
    );
  mac_control_ledrx_cnt_163_1797 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_310,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_163_FFX_RST,
      O => mac_control_ledrx_cnt_163
    );
  mac_control_ledrx_cnt_163_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_163_FFX_RST
    );
  mac_control_txfifowerr_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(24),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(24)
    );
  mac_control_txfifowerr_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(26),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(26)
    );
  mac_control_txfifowerr_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(28),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(28)
    );
  mac_control_txfifowerr_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(31),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(31)
    );
  mac_control_txfifowerr_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(30),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(30)
    );
  mac_control_rxoferr_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(18),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(18)
    );
  mac_control_rxoferr_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(20),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(20)
    );
  mac_control_rxoferr_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(27),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(27)
    );
  mac_control_rxoferr_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(22),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(22)
    );
  mac_control_rxoferr_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(25),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(25)
    );
  mac_control_rxoferr_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(29),
      CE => mac_control_n0053,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0052,
      O => mac_control_rxoferr_cnt(29)
    );
  mac_control_txfifowerr_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(12),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(12)
    );
  mac_control_txfifowerr_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(14),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(14)
    );
  mac_control_txfifowerr_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(21),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(21)
    );
  mac_control_txfifowerr_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(16),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(16)
    );
  mac_control_txfifowerr_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(19),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(19)
    );
  mac_control_txfifowerr_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(23),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(23)
    );
  rx_output_bp_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(8),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_8_FFX_RST,
      O => rx_output_bp(8)
    );
  rx_output_bp_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_8_FFX_RST
    );
  rx_output_bp_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(10),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_10_FFX_RST,
      O => rx_output_bp(10)
    );
  rx_output_bp_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_10_FFX_RST
    );
  rx_output_bp_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(13),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_12_FFY_RST,
      O => rx_output_bp(13)
    );
  rx_output_bp_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_12_FFY_RST
    );
  rx_output_bp_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(12),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_12_FFX_RST,
      O => rx_output_bp(12)
    );
  rx_output_bp_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_12_FFX_RST
    );
  rx_output_bp_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(15),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_14_FFY_RST,
      O => rx_output_bp(15)
    );
  rx_output_bp_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_14_FFY_RST
    );
  rx_output_bp_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(14),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_14_FFX_RST,
      O => rx_output_bp(14)
    );
  rx_output_bp_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_14_FFX_RST
    );
  tx_output_bcnt_38_1798 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_171,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_38_FFY_RST,
      O => tx_output_bcnt_38
    );
  tx_output_bcnt_38_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_38_FFY_RST
    );
  mac_control_txfifowerr_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_lut2_16,
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(0)
    );
  mac_control_txfifowerr_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(5),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(5)
    );
  mac_control_txfifowerr_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(2),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(2)
    );
  mac_control_txfifowerr_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(9),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(9)
    );
  mac_control_txfifowerr_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(4),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(4)
    );
  mac_control_txfifowerr_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(7),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(7)
    );
  mac_control_txfifowerr_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(11),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(11)
    );
  mac_control_rxphyerr_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(1),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(1)
    );
  mac_control_rxphyerr_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_lut2_16,
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(0)
    );
  mac_control_rxphyerr_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(7),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(7)
    );
  mac_control_rxphyerr_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(2),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(2)
    );
  mac_control_rxphyerr_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(5),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(5)
    );
  mac_control_ledrx_cnt_156_1799 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_303,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_155_FFY_RST,
      O => mac_control_ledrx_cnt_156
    );
  mac_control_ledrx_cnt_155_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_155_FFY_RST
    );
  mac_control_ledrx_cnt_160_1800 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_307,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_159_FFY_RST,
      O => mac_control_ledrx_cnt_160
    );
  mac_control_ledrx_cnt_159_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_159_FFY_RST
    );
  mac_control_ledrx_cnt_155_1801 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_302,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_155_FFX_RST,
      O => mac_control_ledrx_cnt_155
    );
  mac_control_ledrx_cnt_155_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_155_FFX_RST
    );
  mac_control_ledrx_cnt_158_1802 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_305,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_157_FFY_RST,
      O => mac_control_ledrx_cnt_158
    );
  mac_control_ledrx_cnt_157_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_157_FFY_RST
    );
  mac_control_ledrx_cnt_157_1803 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_304,
      CE => mac_control_n0040,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_cnt_157_FFX_RST,
      O => mac_control_ledrx_cnt_157
    );
  mac_control_ledrx_cnt_157_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_157_FFX_RST
    );
  mac_control_rxphyerr_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(28),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(28)
    );
  mac_control_rxphyerr_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(30),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(30)
    );
  mac_control_rxfifowerr_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(1),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(1)
    );
  mac_control_rxfifowerr_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(7),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(7)
    );
  mac_control_rxfifowerr_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_lut2_16,
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(0)
    );
  mac_control_rxfifowerr_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(5),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(5)
    );
  mac_control_rxphyerr_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(10),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(10)
    );
  mac_control_rxphyerr_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(12),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(12)
    );
  mac_control_rxphyerr_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(15),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(15)
    );
  mac_control_rxphyerr_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(19),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(19)
    );
  mac_control_rxphyerr_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(14),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(14)
    );
  mac_control_rxphyerr_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(17),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(17)
    );
  tx_fifocheck_diff_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_2_FFX_RST,
      O => tx_fifocheck_diff(2)
    );
  tx_fifocheck_diff_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_2_FFX_RST
    );
  tx_fifocheck_diff_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_4_FFX_RST,
      O => tx_fifocheck_diff(4)
    );
  tx_fifocheck_diff_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_4_FFX_RST
    );
  tx_fifocheck_diff_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_6_FFX_RST,
      O => tx_fifocheck_diff(6)
    );
  tx_fifocheck_diff_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_6_FFX_RST
    );
  mac_control_rxfifowerr_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(2),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(2)
    );
  mac_control_rxfifowerr_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(4),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(4)
    );
  mac_control_rxfifowerr_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(11),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(11)
    );
  mac_control_rxfifowerr_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(6),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(6)
    );
  mac_control_rxfifowerr_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(9),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(9)
    );
  mac_control_rxfifowerr_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(13),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(13)
    );
  mac_control_rxphyerr_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(16),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(16)
    );
  mac_control_rxphyerr_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(18),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(18)
    );
  mac_control_rxphyerr_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(21),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(21)
    );
  mac_control_rxphyerr_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(25),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(25)
    );
  mac_control_rxphyerr_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(20),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(20)
    );
  mac_control_rxphyerr_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(23),
      CE => mac_control_n0051,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0050,
      O => mac_control_rxphyerr_cnt(23)
    );
  mac_control_rxfifowerr_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(20),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(20)
    );
  mac_control_rxfifowerr_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(22),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(22)
    );
  mac_control_rxfifowerr_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(29),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(29)
    );
  mac_control_rxfifowerr_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(24),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(24)
    );
  mac_control_rxfifowerr_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(27),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(27)
    );
  mac_control_rxfifowerr_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(31),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(31)
    );
  mac_control_rxfifowerr_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(14),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(14)
    );
  mac_control_rxfifowerr_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(16),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(16)
    );
  mac_control_rxfifowerr_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(23),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(23)
    );
  mac_control_rxfifowerr_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(18),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(18)
    );
  mac_control_rxfifowerr_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(21),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(21)
    );
  mac_control_rxfifowerr_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(25),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(25)
    );
  mac_control_rxfifowerr_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(8),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(8)
    );
  mac_control_rxfifowerr_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(10),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(10)
    );
  mac_control_rxfifowerr_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(17),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(17)
    );
  mac_control_rxfifowerr_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(12),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(12)
    );
  mac_control_rxfifowerr_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(15),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(15)
    );
  mac_control_rxfifowerr_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(19),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(19)
    );
  mac_control_rxfifowerr_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(26),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(26)
    );
  mac_control_rxfifowerr_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(28),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(28)
    );
  mac_control_rxfifowerr_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(30),
      CE => mac_control_n0049,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0048,
      O => mac_control_rxfifowerr_cnt(30)
    );
  mac_control_txfifowerr_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(3),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(3)
    );
  mac_control_txfifowerr_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(1),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(1)
    );
  rx_output_fifo_BU65 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1908,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N13_FFX_RST,
      O => rx_output_fifo_N13
    );
  rx_output_fifo_N13_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N13_FFX_RST
    );
  rx_output_fifo_BU77 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1910,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N11_FFX_RST,
      O => rx_output_fifo_N11
    );
  rx_output_fifo_N11_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N11_FFX_RST
    );
  mac_control_txfifowerr_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(6),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(6)
    );
  mac_control_txfifowerr_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(8),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(8)
    );
  mac_control_txfifowerr_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(15),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(15)
    );
  mac_control_txfifowerr_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(10),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(10)
    );
  mac_control_txfifowerr_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(13),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(13)
    );
  mac_control_txfifowerr_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(17),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(17)
    );
  rx_output_bp_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(1),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_0_FFY_RST,
      O => rx_output_bp(1)
    );
  rx_output_bp_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_0_FFY_RST
    );
  rx_output_bp_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(3),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_2_FFY_RST,
      O => rx_output_bp(3)
    );
  rx_output_bp_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_2_FFY_RST
    );
  rx_output_bp_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(0),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_0_FFX_RST,
      O => rx_output_bp(0)
    );
  rx_output_bp_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_0_FFX_RST
    );
  rx_output_bp_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(5),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_4_FFY_RST,
      O => rx_output_bp(5)
    );
  rx_output_bp_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_4_FFY_RST
    );
  tx_output_bcnt_49_1804 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_182,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_49_FFX_RST,
      O => tx_output_bcnt_49
    );
  tx_output_bcnt_49_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_49_FFX_RST
    );
  tx_output_bcnt_52_1805 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_185,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_51_FFY_RST,
      O => tx_output_bcnt_52
    );
  tx_output_bcnt_51_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_51_FFY_RST
    );
  tx_output_bcnt_51_1806 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_184,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_51_FFX_RST,
      O => tx_output_bcnt_51
    );
  tx_output_bcnt_51_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_51_FFX_RST
    );
  tx_output_bcnt_53_1807 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_186,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_53_FFX_RST,
      O => tx_output_bcnt_53
    );
  tx_output_bcnt_53_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_53_FFX_RST
    );
  tx_fifocheck_diff_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_14_FFX_RST,
      O => tx_fifocheck_diff(14)
    );
  tx_fifocheck_diff_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_14_FFX_RST
    );
  mac_control_ledtx_cnt_144_1808 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_291,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_143_FFY_RST,
      O => mac_control_ledtx_cnt_144
    );
  mac_control_ledtx_cnt_143_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_143_FFY_RST
    );
  mac_control_ledtx_cnt_148_1809 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_295,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_147_FFY_RST,
      O => mac_control_ledtx_cnt_148
    );
  mac_control_ledtx_cnt_147_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_147_FFY_RST
    );
  mac_control_ledtx_cnt_143_1810 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_290,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_143_FFX_RST,
      O => mac_control_ledtx_cnt_143
    );
  mac_control_ledtx_cnt_143_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_143_FFX_RST
    );
  mac_control_ledtx_cnt_146_1811 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_293,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_145_FFY_RST,
      O => mac_control_ledtx_cnt_146
    );
  mac_control_ledtx_cnt_145_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_145_FFY_RST
    );
  mac_control_ledtx_cnt_145_1812 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_292,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_145_FFX_RST,
      O => mac_control_ledtx_cnt_145
    );
  mac_control_ledtx_cnt_145_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_145_FFX_RST
    );
  mac_control_txfifowerr_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(18),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(18)
    );
  mac_control_txfifowerr_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(20),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(20)
    );
  mac_control_txfifowerr_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(27),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(27)
    );
  mac_control_txfifowerr_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(22),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(22)
    );
  mac_control_txfifowerr_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(25),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(25)
    );
  mac_control_txfifowerr_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(29),
      CE => mac_control_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0046,
      O => mac_control_txfifowerr_cnt(29)
    );
  mac_control_ledtx_cnt_151_1813 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_298,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_151_FFX_RST,
      O => mac_control_ledtx_cnt_151
    );
  mac_control_ledtx_cnt_151_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_151_FFX_RST
    );
  rx_output_fifo_BU47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1905,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N17_FFY_RST,
      O => rx_output_fifo_N16
    );
  rx_output_fifo_N17_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N17_FFY_RST
    );
  rx_output_fifo_BU41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1904,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N17_FFX_RST,
      O => rx_output_fifo_N17
    );
  rx_output_fifo_N17_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N17_FFX_RST
    );
  rx_output_fifo_BU59 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1907,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N15_FFY_RST,
      O => rx_output_fifo_N14
    );
  rx_output_fifo_N15_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N15_FFY_RST
    );
  rx_output_fifo_BU82 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1911,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N11_FFY_RST,
      O => rx_output_fifo_N10
    );
  rx_output_fifo_N11_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N11_FFY_RST
    );
  rx_output_fifo_BU53 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1906,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N15_FFX_RST,
      O => rx_output_fifo_N15
    );
  rx_output_fifo_N15_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N15_FFX_RST
    );
  rx_output_fifo_BU71 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1909,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N13_FFY_RST,
      O => rx_output_fifo_N12
    );
  rx_output_fifo_N13_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N13_FFY_RST
    );
  rx_fifocheck_diff_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_0_FFX_RST,
      O => rx_fifocheck_diff(0)
    );
  rx_fifocheck_diff_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_0_FFX_RST
    );
  rx_fifocheck_diff_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_2_FFX_RST,
      O => rx_fifocheck_diff(2)
    );
  rx_fifocheck_diff_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_2_FFX_RST
    );
  rx_fifocheck_diff_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_4_FFY_RST,
      O => rx_fifocheck_diff(5)
    );
  rx_fifocheck_diff_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_4_FFY_RST
    );
  rx_fifocheck_diff_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_8_FFY_RST,
      O => rx_fifocheck_diff(9)
    );
  rx_fifocheck_diff_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_8_FFY_RST
    );
  rx_fifocheck_diff_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_4_FFX_RST,
      O => rx_fifocheck_diff(4)
    );
  rx_fifocheck_diff_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_4_FFX_RST
    );
  rx_fifocheck_diff_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_6_FFY_RST,
      O => rx_fifocheck_diff(7)
    );
  rx_fifocheck_diff_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_6_FFY_RST
    );
  rx_output_bp_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(2),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_2_FFX_RST,
      O => rx_output_bp(2)
    );
  rx_output_bp_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_2_FFX_RST
    );
  rx_output_bp_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(4),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_4_FFX_RST,
      O => rx_output_bp(4)
    );
  rx_output_bp_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_4_FFX_RST
    );
  rx_output_bp_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(7),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_6_FFY_RST,
      O => rx_output_bp(7)
    );
  rx_output_bp_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_6_FFY_RST
    );
  rx_output_bp_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(11),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_10_FFY_RST,
      O => rx_output_bp(11)
    );
  rx_output_bp_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_10_FFY_RST
    );
  rx_output_bp_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(6),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_6_FFX_RST,
      O => rx_output_bp(6)
    );
  rx_output_bp_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_6_FFX_RST
    );
  rx_output_bp_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(9),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_8_FFY_RST,
      O => rx_output_bp(9)
    );
  rx_output_bp_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_8_FFY_RST
    );
  mac_control_phyrstcnt_111_1814 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_258,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_111_FFX_RST,
      O => mac_control_phyrstcnt_111
    );
  mac_control_phyrstcnt_111_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_111_FFX_RST
    );
  mac_control_phyrstcnt_114_1815 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_261,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_113_FFY_RST,
      O => mac_control_phyrstcnt_114
    );
  mac_control_phyrstcnt_113_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_113_FFY_RST
    );
  mac_control_phyrstcnt_118_1816 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_265,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_117_FFY_RST,
      O => mac_control_phyrstcnt_118
    );
  mac_control_phyrstcnt_117_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_117_FFY_RST
    );
  mac_control_phyrstcnt_113_1817 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_260,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_113_FFX_RST,
      O => mac_control_phyrstcnt_113
    );
  mac_control_phyrstcnt_113_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_113_FFX_RST
    );
  mac_control_phyrstcnt_116_1818 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_263,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_115_FFY_RST,
      O => mac_control_phyrstcnt_116
    );
  mac_control_phyrstcnt_115_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_115_FFY_RST
    );
  mac_control_txf_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(24),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(24)
    );
  mac_control_txf_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(26),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(26)
    );
  mac_control_txf_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(29),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(29)
    );
  rx_output_macnt_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_95,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_0_FFY_RST,
      O => addr3ext(0)
    );
  addr3ext_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_0_FFY_RST
    );
  mac_control_txf_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(28),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(28)
    );
  mac_control_txf_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(31),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(31)
    );
  tx_output_bcnt_39_1819 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_172,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_39_FFX_RST,
      O => tx_output_bcnt_39
    );
  tx_output_bcnt_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_39_FFX_RST
    );
  tx_output_bcnt_42_1820 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_175,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_41_FFY_RST,
      O => tx_output_bcnt_42
    );
  tx_output_bcnt_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_41_FFY_RST
    );
  tx_output_bcnt_41_1821 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_174,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_41_FFX_RST,
      O => tx_output_bcnt_41
    );
  tx_output_bcnt_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_41_FFX_RST
    );
  tx_output_bcnt_44_1822 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_177,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_43_FFY_RST,
      O => tx_output_bcnt_44
    );
  tx_output_bcnt_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_43_FFY_RST
    );
  tx_output_bcnt_43_1823 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_176,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_43_FFX_RST,
      O => tx_output_bcnt_43
    );
  tx_output_bcnt_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_43_FFX_RST
    );
  tx_output_bcnt_46_1824 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_179,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_45_FFY_RST,
      O => tx_output_bcnt_46
    );
  tx_output_bcnt_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_45_FFY_RST
    );
  tx_output_bcnt_45_1825 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_178,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_45_FFX_RST,
      O => tx_output_bcnt_45
    );
  tx_output_bcnt_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_45_FFX_RST
    );
  tx_output_bcnt_48_1826 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_181,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_47_FFY_RST,
      O => tx_output_bcnt_48
    );
  tx_output_bcnt_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_47_FFY_RST
    );
  tx_output_bcnt_47_1827 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_180,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_47_FFX_RST,
      O => tx_output_bcnt_47
    );
  tx_output_bcnt_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_47_FFX_RST
    );
  tx_output_bcnt_50_1828 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_183,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_49_FFY_RST,
      O => tx_output_bcnt_50
    );
  tx_output_bcnt_49_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_49_FFY_RST
    );
  rx_fifocheck_diff_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_0_FFY_RST,
      O => rx_fifocheck_diff(1)
    );
  rx_fifocheck_diff_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_0_FFY_RST
    );
  rx_fifocheck_diff_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_2_FFY_RST,
      O => rx_fifocheck_diff(3)
    );
  rx_fifocheck_diff_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_2_FFY_RST
    );
  rx_fifocheck_diff_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_12_FFX_RST,
      O => rx_fifocheck_diff(12)
    );
  rx_fifocheck_diff_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_12_FFX_RST
    );
  rx_fifocheck_diff_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_14_FFX_RST,
      O => rx_fifocheck_diff(14)
    );
  rx_fifocheck_diff_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_14_FFX_RST
    );
  tx_fifocheck_diff_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_0_FFY_RST,
      O => tx_fifocheck_diff(1)
    );
  tx_fifocheck_diff_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_0_FFY_RST
    );
  tx_fifocheck_diff_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_0_FFX_RST,
      O => tx_fifocheck_diff(0)
    );
  tx_fifocheck_diff_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_0_FFX_RST
    );
  mac_control_ledtx_cnt_147_1829 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_294,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_147_FFX_RST,
      O => mac_control_ledtx_cnt_147
    );
  mac_control_ledtx_cnt_147_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_147_FFX_RST
    );
  mac_control_ledtx_cnt_150_1830 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_297,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_149_FFY_RST,
      O => mac_control_ledtx_cnt_150
    );
  mac_control_ledtx_cnt_149_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_149_FFY_RST
    );
  mac_control_ledtx_cnt_149_1831 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_296,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_149_FFX_RST,
      O => mac_control_ledtx_cnt_149
    );
  mac_control_ledtx_cnt_149_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_149_FFX_RST
    );
  mac_control_ledtx_cnt_152_1832 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_299,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_151_FFY_RST,
      O => mac_control_ledtx_cnt_152
    );
  mac_control_ledtx_cnt_151_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_151_FFY_RST
    );
  mac_control_ledtx_cnt_153_1833 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_300,
      CE => mac_control_n0038,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_cnt_153_FFX_RST,
      O => mac_control_ledtx_cnt_153
    );
  mac_control_ledtx_cnt_153_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_153_FFX_RST
    );
  mac_control_phyrstcnt_127_1834 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_274,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_127_FFX_RST,
      O => mac_control_phyrstcnt_127
    );
  mac_control_phyrstcnt_127_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_127_FFX_RST
    );
  mac_control_phyrstcnt_130_1835 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_277,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_129_FFY_RST,
      O => mac_control_phyrstcnt_130
    );
  mac_control_phyrstcnt_129_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_129_FFY_RST
    );
  mac_control_phyrstcnt_134_1836 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_281,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_133_FFY_RST,
      O => mac_control_phyrstcnt_134
    );
  mac_control_phyrstcnt_133_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_133_FFY_RST
    );
  mac_control_phyrstcnt_129_1837 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_276,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_129_FFX_RST,
      O => mac_control_phyrstcnt_129
    );
  mac_control_phyrstcnt_129_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_129_FFX_RST
    );
  mac_control_phyrstcnt_132_1838 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_279,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_131_FFY_RST,
      O => mac_control_phyrstcnt_132
    );
  mac_control_phyrstcnt_131_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_131_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_32_1839 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_165,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_32_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_32
    );
  mac_control_PHY_status_MII_Interface_mdccnt_32_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_32_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_34_1840 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_167,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_33_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_34
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_33_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_1841 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_166,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_33_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_33
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_33_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_36_1842 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_169,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_35_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_36
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_35_FFY_RST
    );
  mac_control_phyrstcnt_110_1843 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_257,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_110_FFY_RST,
      O => mac_control_phyrstcnt_110
    );
  mac_control_phyrstcnt_110_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_110_FFY_RST
    );
  rx_fifocheck_diff_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_6_FFX_RST,
      O => rx_fifocheck_diff(6)
    );
  rx_fifocheck_diff_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_6_FFX_RST
    );
  rx_fifocheck_diff_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_8_FFX_RST,
      O => rx_fifocheck_diff(8)
    );
  rx_fifocheck_diff_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_8_FFX_RST
    );
  rx_fifocheck_diff_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_10_FFY_RST,
      O => rx_fifocheck_diff(11)
    );
  rx_fifocheck_diff_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_10_FFY_RST
    );
  rx_fifocheck_diff_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_14_FFY_RST,
      O => rx_fifocheck_diff(15)
    );
  rx_fifocheck_diff_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_14_FFY_RST
    );
  rx_fifocheck_diff_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_10_FFX_RST,
      O => rx_fifocheck_diff(10)
    );
  rx_fifocheck_diff_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_10_FFX_RST
    );
  rx_fifocheck_diff_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_12_FFY_RST,
      O => rx_fifocheck_diff(13)
    );
  rx_fifocheck_diff_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_12_FFY_RST
    );
  mac_control_phyrstcnt_137_1844 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_284,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_137_FFX_RST,
      O => mac_control_phyrstcnt_137
    );
  mac_control_phyrstcnt_137_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_137_FFX_RST
    );
  rx_input_memio_macnt_72_1845 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_221,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_71_FFY_RST,
      O => rx_input_memio_macnt_72
    );
  rx_input_memio_macnt_71_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_71_FFY_RST
    );
  rx_input_memio_macnt_70_1846 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_219,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_70_FFY_RST,
      O => rx_input_memio_macnt_70
    );
  rx_input_memio_macnt_70_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_70_FFY_RST
    );
  mac_control_phyrstcnt_139_1847 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_286,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_139_FFX_RST,
      O => mac_control_phyrstcnt_139
    );
  mac_control_phyrstcnt_139_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_139_FFX_RST
    );
  mac_control_phyrstcnt_141_1848 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_288,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_141_FFX_RST,
      O => mac_control_phyrstcnt_141
    );
  mac_control_phyrstcnt_141_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_141_FFX_RST
    );
  rx_input_memio_macnt_74_1849 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_223,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_73_FFY_RST,
      O => rx_input_memio_macnt_74
    );
  rx_input_memio_macnt_73_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_73_FFY_RST
    );
  tx_fifocheck_diff_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_8_FFX_RST,
      O => tx_fifocheck_diff(8)
    );
  tx_fifocheck_diff_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_8_FFX_RST
    );
  tx_fifocheck_diff_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_10_FFX_RST,
      O => tx_fifocheck_diff(10)
    );
  tx_fifocheck_diff_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_10_FFX_RST
    );
  tx_fifocheck_diff_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_12_FFX_RST,
      O => tx_fifocheck_diff(12)
    );
  tx_fifocheck_diff_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_12_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_1850 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_168,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_35_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_35
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_35_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_37_1851 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_170,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_37_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_37
    );
  mac_control_PHY_status_MII_Interface_mdccnt_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_37_FFX_RST
    );
  mac_control_txf_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(1),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(1)
    );
  tx_input_addr_19_1852 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_130,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_19_FFX_RST,
      O => tx_input_addr_19
    );
  tx_input_addr_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_19_FFX_RST
    );
  tx_input_addr_21_1853 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_132,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_21_FFX_RST,
      O => tx_input_addr_21
    );
  tx_input_addr_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_21_FFX_RST
    );
  tx_input_addr_24_1854 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_135,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_23_FFY_RST,
      O => tx_input_addr_24
    );
  tx_input_addr_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_23_FFY_RST
    );
  tx_input_addr_28_1855 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_139,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_27_FFY_RST,
      O => tx_input_addr_28
    );
  tx_input_addr_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_27_FFY_RST
    );
  tx_input_addr_23_1856 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_134,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_23_FFX_RST,
      O => tx_input_addr_23
    );
  tx_input_addr_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_23_FFX_RST
    );
  tx_input_addr_26_1857 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_137,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_25_FFY_RST,
      O => tx_input_addr_26
    );
  tx_input_addr_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_25_FFY_RST
    );
  mac_control_txf_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(12),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(12)
    );
  mac_control_txf_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(14),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(14)
    );
  mac_control_txf_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(17),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(17)
    );
  mac_control_txf_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(21),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(21)
    );
  mac_control_txf_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(16),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(16)
    );
  mac_control_txf_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(19),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(19)
    );
  rx_output_macnt_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_98,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_3_FFX_RST,
      O => addr3ext(3)
    );
  addr3ext_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_3_FFX_RST
    );
  rx_output_macnt_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_100,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_5_FFX_RST,
      O => addr3ext(5)
    );
  addr3ext_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_5_FFX_RST
    );
  rx_output_macnt_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_103,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_7_FFY_RST,
      O => addr3ext(8)
    );
  addr3ext_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_7_FFY_RST
    );
  rx_output_macnt_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_102,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_7_FFX_RST,
      O => addr3ext(7)
    );
  addr3ext_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_7_FFX_RST
    );
  rx_output_macnt_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_105,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_9_FFY_RST,
      O => addr3ext(10)
    );
  addr3ext_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_9_FFY_RST
    );
  rx_output_macnt_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_107,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_11_FFY_RST,
      O => addr3ext(12)
    );
  addr3ext_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_11_FFY_RST
    );
  mac_control_txf_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(18),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(18)
    );
  mac_control_txf_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(20),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(20)
    );
  mac_control_txf_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(23),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(23)
    );
  mac_control_txf_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(27),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(27)
    );
  mac_control_txf_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(22),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(22)
    );
  mac_control_txf_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(25),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(25)
    );
  mac_control_txf_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_lut2_16,
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(0)
    );
  mac_control_txf_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(2),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(2)
    );
  mac_control_txf_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(5),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(5)
    );
  mac_control_txf_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(9),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(9)
    );
  mac_control_txf_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(4),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(4)
    );
  mac_control_txf_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(7),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(7)
    );
  mac_control_txf_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(6),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(6)
    );
  mac_control_txf_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(8),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(8)
    );
  mac_control_txf_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(11),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(11)
    );
  mac_control_txf_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(15),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(15)
    );
  mac_control_txf_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(10),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(10)
    );
  mac_control_txf_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(13),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(13)
    );
  rx_output_macnt_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_97,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_1_FFY_RST,
      O => addr3ext(2)
    );
  addr3ext_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_1_FFY_RST
    );
  mac_control_txf_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(30),
      CE => mac_control_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0042,
      O => mac_control_txf_cnt(30)
    );
  rx_output_macnt_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_96,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_1_FFX_RST,
      O => addr3ext(1)
    );
  addr3ext_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_1_FFX_RST
    );
  rx_output_macnt_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_99,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_3_FFY_RST,
      O => addr3ext(4)
    );
  addr3ext_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_3_FFY_RST
    );
  rx_output_macnt_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_101,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_5_FFY_RST,
      O => addr3ext(6)
    );
  addr3ext_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_5_FFY_RST
    );
  rx_input_memio_crcl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(6),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_6_FFY_RST,
      O => rx_input_memio_crcl(6)
    );
  rx_input_memio_crcl_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_6_FFY_RST
    );
  rx_fifocheck_bpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_11_FFY_RST,
      O => rx_fifocheck_bpl(10)
    );
  rx_fifocheck_bpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_11_FFY_RST
    );
  rx_fifocheck_bpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_11_FFX_RST,
      O => rx_fifocheck_bpl(11)
    );
  rx_fifocheck_bpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_11_FFX_RST
    );
  rx_fifocheck_bpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_13_FFY_RST,
      O => rx_fifocheck_bpl(12)
    );
  rx_fifocheck_bpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_13_FFY_RST
    );
  rx_fifocheck_bpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_13_FFX_RST,
      O => rx_fifocheck_bpl(13)
    );
  rx_fifocheck_bpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_13_FFX_RST
    );
  rx_fifocheck_bpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_15_FFY_RST,
      O => rx_fifocheck_bpl(14)
    );
  rx_fifocheck_bpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_15_FFY_RST
    );
  rx_fifocheck_bpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_15_FFX_RST,
      O => rx_fifocheck_bpl(15)
    );
  rx_fifocheck_bpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_15_FFX_RST
    );
  tx_output_crcsell_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd3,
      CE => tx_output_crcsell_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcsell_3_FFY_RST,
      O => tx_output_crcsell(2)
    );
  tx_output_crcsell_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcsell_3_FFY_RST
    );
  tx_output_crcsell_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd7,
      CE => tx_output_crcsell_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcsell_3_FFX_RST,
      O => tx_output_crcsell(3)
    );
  tx_output_crcsell_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcsell_3_FFX_RST
    );
  tx_input_cs_FFd5_1858 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd5_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd5_FFY_RST,
      O => tx_input_cs_FFd5
    );
  tx_input_cs_FFd5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd5_FFY_RST
    );
  rx_output_macnt_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_104,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_9_FFX_RST,
      O => addr3ext(9)
    );
  addr3ext_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_9_FFX_RST
    );
  rx_output_macnt_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_106,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_11_FFX_RST,
      O => addr3ext(11)
    );
  addr3ext_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_11_FFX_RST
    );
  rx_output_macnt_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_109,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_13_FFY_RST,
      O => addr3ext(14)
    );
  addr3ext_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_13_FFY_RST
    );
  rx_output_macnt_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_108,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_13_FFX_RST,
      O => addr3ext(13)
    );
  addr3ext_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_13_FFX_RST
    );
  rx_output_macnt_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_110,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_15_FFX_RST,
      O => addr3ext(15)
    );
  addr3ext_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_15_FFX_RST
    );
  rx_output_fifo_BU214 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2834,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N7_FFX_RST,
      O => rx_output_fifo_N7
    );
  rx_output_fifo_N7_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N7_FFX_RST
    );
  rx_output_fifo_BU226 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2836,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N5_FFX_RST,
      O => rx_output_fifo_N5
    );
  rx_output_fifo_N5_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N5_FFX_RST
    );
  rx_output_fifo_BU238 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2838,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N3_FFX_RST,
      O => rx_output_fifo_N3
    );
  rx_output_fifo_N3_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N3_FFX_RST
    );
  memcontroller_dnl2_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(9),
      CE => memcontroller_dnl2_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_9_FFX_RST,
      O => memcontroller_dnl2(9)
    );
  memcontroller_dnl2_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_9_FFX_RST
    );
  rx_input_memio_crcl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(7),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_7_FFY_RST,
      O => rx_input_memio_crcl(7)
    );
  rx_input_memio_crcl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_7_FFY_RST
    );
  rx_input_memio_addrchk_datal_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_1_FFX_RST,
      O => rx_input_memio_addrchk_datal(1)
    );
  rx_input_memio_addrchk_datal_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_1_FFX_RST
    );
  rx_input_memio_addrchk_datal_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_1_FFY_RST,
      O => rx_input_memio_addrchk_datal(0)
    );
  rx_input_memio_addrchk_datal_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_1_FFY_RST
    );
  rx_input_memio_addrchk_datal_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_3_FFY_RST,
      O => rx_input_memio_addrchk_datal(2)
    );
  rx_input_memio_addrchk_datal_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_3_FFY_RST
    );
  rx_input_memio_addrchk_datal_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_3_FFX_RST,
      O => rx_input_memio_addrchk_datal(3)
    );
  rx_input_memio_addrchk_datal_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_3_FFX_RST
    );
  rx_input_memio_addrchk_datal_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_5_FFY_RST,
      O => rx_input_memio_addrchk_datal(4)
    );
  rx_input_memio_addrchk_datal_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_5_FFY_RST
    );
  rx_input_memio_addrchk_datal_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_5_FFX_RST,
      O => rx_input_memio_addrchk_datal(5)
    );
  rx_input_memio_addrchk_datal_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_5_FFX_RST
    );
  rx_input_memio_addrchk_datal_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_7_FFY_RST,
      O => rx_input_memio_addrchk_datal(6)
    );
  rx_input_memio_addrchk_datal_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_7_FFY_RST
    );
  rx_input_memio_addrchk_datal_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_7_FFX_RST,
      O => rx_input_memio_addrchk_datal(7)
    );
  rx_input_memio_addrchk_datal_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_7_FFX_RST
    );
  rx_fifocheck_fbbpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_1_FFY_RST,
      O => rx_fifocheck_fbbpl(0)
    );
  rx_fifocheck_fbbpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_1_FFY_RST
    );
  rx_input_memio_addrchk_datal_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_9_FFY_RST,
      O => rx_input_memio_addrchk_datal(8)
    );
  rx_input_memio_addrchk_datal_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_9_FFY_RST
    );
  rx_input_memio_addrchk_datal_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_9_FFX_RST,
      O => rx_input_memio_addrchk_datal(9)
    );
  rx_input_memio_addrchk_datal_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_9_FFX_RST
    );
  rx_fifocheck_fbbpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_1_FFX_RST,
      O => rx_fifocheck_fbbpl(1)
    );
  rx_fifocheck_fbbpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_1_FFX_RST
    );
  slowclock_rxcrcerrl_1859 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_rxcrcerrl_GROM,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => rxcrcerr,
      SRST => slowclock_rxcrcerrl_LOGIC_ZERO,
      O => slowclock_rxcrcerrl
    );
  mac_control_phyrstcnt_115_1860 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_262,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_115_FFX_RST,
      O => mac_control_phyrstcnt_115
    );
  mac_control_phyrstcnt_115_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_115_FFX_RST
    );
  mac_control_phyrstcnt_117_1861 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_264,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_117_FFX_RST,
      O => mac_control_phyrstcnt_117
    );
  mac_control_phyrstcnt_117_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_117_FFX_RST
    );
  mac_control_phyrstcnt_120_1862 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_267,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_119_FFY_RST,
      O => mac_control_phyrstcnt_120
    );
  mac_control_phyrstcnt_119_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_119_FFY_RST
    );
  mac_control_phyrstcnt_119_1863 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_266,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_119_FFX_RST,
      O => mac_control_phyrstcnt_119
    );
  mac_control_phyrstcnt_119_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_119_FFX_RST
    );
  mac_control_phyrstcnt_122_1864 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_269,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_121_FFY_RST,
      O => mac_control_phyrstcnt_122
    );
  mac_control_phyrstcnt_121_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_121_FFY_RST
    );
  mac_control_phyrstcnt_131_1865 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_278,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_131_FFX_RST,
      O => mac_control_phyrstcnt_131
    );
  mac_control_phyrstcnt_131_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_131_FFX_RST
    );
  mac_control_phyrstcnt_133_1866 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_280,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_133_FFX_RST,
      O => mac_control_phyrstcnt_133
    );
  mac_control_phyrstcnt_133_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_133_FFX_RST
    );
  mac_control_phyrstcnt_136_1867 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_283,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_135_FFY_RST,
      O => mac_control_phyrstcnt_136
    );
  mac_control_phyrstcnt_135_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_135_FFY_RST
    );
  mac_control_phyrstcnt_140_1868 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_287,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_139_FFY_RST,
      O => mac_control_phyrstcnt_140
    );
  mac_control_phyrstcnt_139_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_139_FFY_RST
    );
  mac_control_phyrstcnt_135_1869 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_282,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_135_FFX_RST,
      O => mac_control_phyrstcnt_135
    );
  mac_control_phyrstcnt_135_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_135_FFX_RST
    );
  mac_control_phyrstcnt_138_1870 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_285,
      CE => mac_control_N80441,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyrstcnt_137_FFY_RST,
      O => mac_control_phyrstcnt_138
    );
  mac_control_phyrstcnt_137_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_137_FFY_RST
    );
  rx_input_memio_bcntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(1),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_0_FFY_RST,
      O => rx_input_memio_bcntl(1)
    );
  rx_input_memio_bcntl_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_0_FFY_RST
    );
  rx_input_memio_bcntl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(0),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_0_FFX_RST,
      O => rx_input_memio_bcntl(0)
    );
  rx_input_memio_bcntl_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_0_FFX_RST
    );
  rx_input_memio_macnt_71_1871 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_220,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_71_FFX_RST,
      O => rx_input_memio_macnt_71
    );
  rx_input_memio_macnt_71_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_71_FFX_RST
    );
  rx_input_memio_macnt_73_1872 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_222,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_73_FFX_RST,
      O => rx_input_memio_macnt_73
    );
  rx_input_memio_macnt_73_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_73_FFX_RST
    );
  rx_input_memio_macnt_76_1873 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_225,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_75_FFY_RST,
      O => rx_input_memio_macnt_76
    );
  rx_input_memio_macnt_75_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_75_FFY_RST
    );
  rx_input_memio_macnt_80_1874 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_229,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_79_FFY_RST,
      O => rx_input_memio_macnt_80
    );
  rx_input_memio_macnt_79_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_79_FFY_RST
    );
  rx_input_memio_macnt_75_1875 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_224,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_75_FFX_RST,
      O => rx_input_memio_macnt_75
    );
  rx_input_memio_macnt_75_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_75_FFX_RST
    );
  rx_input_memio_macnt_78_1876 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_227,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_77_FFY_RST,
      O => rx_input_memio_macnt_78
    );
  rx_input_memio_macnt_77_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_77_FFY_RST
    );
  rx_input_memio_bcntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(2),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_2_FFX_RST,
      O => rx_input_memio_bcntl(2)
    );
  rx_input_memio_bcntl_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_2_FFX_RST
    );
  rx_input_memio_bcntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(4),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_4_FFX_RST,
      O => rx_input_memio_bcntl(4)
    );
  rx_input_memio_bcntl_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_4_FFX_RST
    );
  rx_input_memio_bcntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(6),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_6_FFX_RST,
      O => rx_input_memio_bcntl(6)
    );
  rx_input_memio_bcntl_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_6_FFX_RST
    );
  rx_input_memio_macnt_83_1877 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_232,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_83_FFX_RST,
      O => rx_input_memio_macnt_83
    );
  rx_input_memio_macnt_83_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_83_FFX_RST
    );
  rx_input_memio_macnt_85_1878 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_234,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_85_FFX_RST,
      O => rx_input_memio_macnt_85
    );
  rx_input_memio_macnt_85_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_85_FFX_RST
    );
  tx_input_addr_25_1879 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_136,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_25_FFX_RST,
      O => tx_input_addr_25
    );
  tx_input_addr_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_25_FFX_RST
    );
  tx_input_addr_27_1880 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_138,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_27_FFX_RST,
      O => tx_input_addr_27
    );
  tx_input_addr_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_27_FFX_RST
    );
  tx_input_addr_30_1881 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_141,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_29_FFY_RST,
      O => tx_input_addr_30
    );
  tx_input_addr_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_29_FFY_RST
    );
  mac_control_rxf_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(1),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(1)
    );
  tx_input_addr_29_1882 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_140,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_29_FFX_RST,
      O => tx_input_addr_29
    );
  tx_input_addr_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_29_FFX_RST
    );
  tx_input_addr_31_1883 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_142,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_31_FFX_RST,
      O => tx_input_addr_31
    );
  tx_input_addr_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_31_FFX_RST
    );
  rx_input_memio_macnt_77_1884 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_226,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_77_FFX_RST,
      O => rx_input_memio_macnt_77
    );
  rx_input_memio_macnt_77_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_77_FFX_RST
    );
  rx_input_memio_macnt_79_1885 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_228,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_79_FFX_RST,
      O => rx_input_memio_macnt_79
    );
  rx_input_memio_macnt_79_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_79_FFX_RST
    );
  rx_input_memio_macnt_82_1886 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_231,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_81_FFY_RST,
      O => rx_input_memio_macnt_82
    );
  rx_input_memio_macnt_81_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_81_FFY_RST
    );
  rx_input_memio_macnt_81_1887 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_230,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_81_FFX_RST,
      O => rx_input_memio_macnt_81
    );
  rx_input_memio_macnt_81_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_81_FFX_RST
    );
  rx_input_memio_macnt_84_1888 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_233,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_83_FFY_RST,
      O => rx_input_memio_macnt_84
    );
  rx_input_memio_macnt_83_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_83_FFY_RST
    );
  mac_control_rxf_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(18),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(18)
    );
  mac_control_rxf_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(20),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(20)
    );
  mac_control_rxf_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(23),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(23)
    );
  mac_control_rxf_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(27),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(27)
    );
  mac_control_rxf_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(22),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(22)
    );
  mac_control_rxf_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(25),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(25)
    );
  mac_control_rxf_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(6),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(6)
    );
  mac_control_rxf_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(8),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(8)
    );
  mac_control_rxf_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(11),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(11)
    );
  mac_control_rxf_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(15),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(15)
    );
  mac_control_rxf_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(10),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(10)
    );
  mac_control_rxf_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(13),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(13)
    );
  mac_control_rxf_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(12),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(12)
    );
  mac_control_rxf_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(14),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(14)
    );
  mac_control_rxf_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(17),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(17)
    );
  mac_control_rxf_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(21),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(21)
    );
  mac_control_rxf_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(16),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(16)
    );
  mac_control_rxf_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(19),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(19)
    );
  rx_input_memio_bcntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(8),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_8_FFX_RST,
      O => rx_input_memio_bcntl(8)
    );
  rx_input_memio_bcntl_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_8_FFX_RST
    );
  rx_input_memio_bcntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(10),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_10_FFX_RST,
      O => rx_input_memio_bcntl(10)
    );
  rx_input_memio_bcntl_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_10_FFX_RST
    );
  rx_input_memio_bcntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(12),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_12_FFX_RST,
      O => rx_input_memio_bcntl(12)
    );
  rx_input_memio_bcntl_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_12_FFX_RST
    );
  tx_input_CNT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(9),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_9_FFX_RST,
      O => tx_input_CNT(9)
    );
  tx_input_CNT_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_9_FFX_RST
    );
  rx_input_GMII_ENDFIN : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_endfin_GROM,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_endfin_FFY_RST,
      O => rx_input_endfin
    );
  rx_input_endfin_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_endfin_FFY_RST
    );
  rx_output_fifo_BU98 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2299,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1553_FFY_RST,
      O => rx_output_fifo_N1552
    );
  rx_output_fifo_N1553_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1553_FFY_RST
    );
  rx_output_fifo_BU91 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2259,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1553_FFX_RST,
      O => rx_output_fifo_N1553
    );
  rx_output_fifo_N1553_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1553_FFX_RST
    );
  tx_output_crcl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(2),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_31_FFY_RST,
      O => tx_output_crcl(2)
    );
  tx_output_crcl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_31_FFY_RST
    );
  tx_output_crcl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(31),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_31_FFX_RST,
      O => tx_output_crcl(31)
    );
  tx_output_crcl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_31_FFX_RST
    );
  mac_control_sclkdelta_1889 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lsclkdelta,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_sclkdelta_FFY_RST,
      O => mac_control_sclkdelta
    );
  mac_control_sclkdelta_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_sclkdelta_FFY_RST
    );
  tx_output_crcenl_1890 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_crcenl_FROM,
      CE => tx_output_crcenl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcenl_FFX_RST,
      O => tx_output_crcenl
    );
  tx_output_crcenl_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcenl_FFX_RST
    );
  rx_input_memio_crcl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(2),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_2_FFY_RST,
      O => rx_input_memio_crcl(2)
    );
  rx_input_memio_crcl_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_2_FFY_RST
    );
  mac_control_rxf_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(30),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(30)
    );
  mac_control_rxf_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_lut2_16,
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(0)
    );
  mac_control_rxf_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(2),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(2)
    );
  mac_control_rxf_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(5),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(5)
    );
  mac_control_rxf_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(9),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(9)
    );
  mac_control_rxf_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(4),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(4)
    );
  mac_control_rxf_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(7),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(7)
    );
  tx_input_addr_18_1891 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_129,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_17_FFY_RST,
      O => tx_input_addr_18
    );
  tx_input_addr_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_17_FFY_RST
    );
  rx_input_memio_bcntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(14),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_14_FFX_RST,
      O => rx_input_memio_bcntl(14)
    );
  rx_input_memio_bcntl_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_14_FFX_RST
    );
  tx_input_addr_22_1892 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_133,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_21_FFY_RST,
      O => tx_input_addr_22
    );
  tx_input_addr_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_21_FFY_RST
    );
  tx_input_addr_17_1893 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_128,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_17_FFX_RST,
      O => tx_input_addr_17
    );
  tx_input_addr_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_17_FFX_RST
    );
  tx_input_addr_20_1894 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_131,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_19_FFY_RST,
      O => tx_input_addr_20
    );
  tx_input_addr_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_19_FFY_RST
    );
  mac_control_rxf_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(24),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(24)
    );
  mac_control_rxf_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(26),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(26)
    );
  mac_control_rxf_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(29),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(29)
    );
  mac_control_rxf_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(28),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(28)
    );
  mac_control_rxf_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(31),
      CE => mac_control_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_n0044,
      O => mac_control_rxf_cnt(31)
    );
  rx_output_fifo_BU176 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N2580,
      CE => rx_output_fifo_N2579,
      CLK => clkio,
      SET => rx_output_fifo_empty_FFX_SET,
      RST => GND,
      O => rx_output_fifo_empty
    );
  rx_output_fifo_empty_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_empty_FFX_SET
    );
  mac_control_PHY_status_MII_Interface_cs_FFd5_1895 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd5_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_cs_FFd5_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_cs_FFd5
    );
  mac_control_PHY_status_MII_Interface_cs_FFd5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_MII_Interface_cs_FFd5_FFX_RST
    );
  rx_input_memio_MA_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_7_FFX_RST,
      O => addr1ext(7)
    );
  addr1ext_7_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_7_FFX_RST
    );
  rx_input_memio_MA_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_5_FFX_RST,
      O => addr1ext(5)
    );
  addr1ext_5_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_5_FFX_RST
    );
  rx_input_memio_MA_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_7_FFY_RST,
      O => addr1ext(6)
    );
  addr1ext_7_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_7_FFY_RST
    );
  rx_input_memio_MA_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_9_FFX_RST,
      O => addr1ext(9)
    );
  addr1ext_9_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_9_FFX_RST
    );
  rx_input_memio_MA_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_9_FFY_RST,
      O => addr1ext(8)
    );
  addr1ext_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_9_FFY_RST
    );
  rx_input_memio_MD_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_1_FFX_RST,
      O => d1(1)
    );
  d1_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_1_FFX_RST
    );
  rx_input_memio_MD_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_1_FFY_RST,
      O => d1(0)
    );
  d1_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_1_FFY_RST
    );
  rx_input_memio_MD_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_3_FFX_RST,
      O => d1(3)
    );
  d1_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_3_FFX_RST
    );
  rx_input_memio_MD_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_3_FFY_RST,
      O => d1(2)
    );
  d1_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_3_FFY_RST
    );
  rx_input_memio_MD_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_5_FFY_RST,
      O => d1(4)
    );
  d1_5_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_5_FFY_RST
    );
  rx_output_fifo_BU208 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2833,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N9_FFY_RST,
      O => rx_output_fifo_N8
    );
  rx_output_fifo_N9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N9_FFY_RST
    );
  rx_output_fifo_BU202 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2832,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N9_FFX_RST,
      O => rx_output_fifo_N9
    );
  rx_output_fifo_N9_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N9_FFX_RST
    );
  rx_output_fifo_BU220 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2835,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N7_FFY_RST,
      O => rx_output_fifo_N6
    );
  rx_output_fifo_N7_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N7_FFY_RST
    );
  rx_output_fifo_BU232 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2837,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N5_FFY_RST,
      O => rx_output_fifo_N4
    );
  rx_output_fifo_N5_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N5_FFY_RST
    );
  rx_output_fifo_BU243 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2839,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N3_FFY_RST,
      O => rx_output_fifo_N2
    );
  rx_output_fifo_N3_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N3_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(3),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_3_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(3)
    );
  mac_control_PHY_status_MII_Interface_statecnt_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_3_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(4),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_5_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(4)
    );
  mac_control_PHY_status_MII_Interface_statecnt_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_5_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(5),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_5_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(5)
    );
  mac_control_PHY_status_MII_Interface_statecnt_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_5_FFX_RST
    );
  rx_input_memio_MA_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_1_FFY_RST,
      O => addr1ext(0)
    );
  addr1ext_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_1_FFY_RST
    );
  rx_input_memio_MA_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_1_FFX_RST,
      O => addr1ext(1)
    );
  addr1ext_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_1_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd3_1896 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd3_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_cs_FFd3_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_cs_FFd3
    );
  mac_control_PHY_status_MII_Interface_cs_FFd3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_MII_Interface_cs_FFd3_FFY_RST
    );
  rx_input_memio_MA_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_3_FFY_RST,
      O => addr1ext(2)
    );
  addr1ext_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_3_FFY_RST
    );
  rx_input_memio_MA_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_3_FFX_RST,
      O => addr1ext(3)
    );
  addr1ext_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_3_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd4_1897 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd4_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_cs_FFd5_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_cs_FFd4
    );
  mac_control_PHY_status_MII_Interface_cs_FFd5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_MII_Interface_cs_FFd5_FFY_RST
    );
  rx_input_memio_MA_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_5_FFY_RST,
      O => addr1ext(4)
    );
  addr1ext_5_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_5_FFY_RST
    );
  rx_output_fifo_BU355 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3618,
      CE => rx_output_fifo_N3617,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_full_FFX_SET,
      RST => GND,
      O => rx_output_fifo_full_0
    );
  rx_output_fifo_full_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_full_FFX_SET
    );
  rx_output_fifo_BU504 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N4755,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_wrcount_0_FFY_RST,
      O => rx_output_fifo_wrcount(1)
    );
  rx_output_fifo_wrcount_0_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_wrcount_0_FFY_RST
    );
  mac_control_bitcnt_104_1898 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_251,
      CE => mac_control_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_bitcnt_104_FFY_RST,
      O => mac_control_bitcnt_104
    );
  mac_control_bitcnt_104_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_104_FFY_RST
    );
  rx_output_fifo_BU498 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N4754,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_wrcount_0_FFX_RST,
      O => rx_output_fifo_wrcount(0)
    );
  rx_output_fifo_wrcount_0_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_wrcount_0_FFX_RST
    );
  mac_control_bitcnt_106_1899 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_253,
      CE => mac_control_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_bitcnt_105_FFY_RST,
      O => mac_control_bitcnt_106
    );
  mac_control_bitcnt_105_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_105_FFY_RST
    );
  tx_output_crcsell_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => tx_output_crcsel(0),
      CE => tx_output_crcsell_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => tx_output_crcsell_1_FFY_SET,
      RST => GND,
      O => tx_output_crcsell(0)
    );
  tx_output_crcsell_1_FFY_SETOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcsell_1_FFY_SET
    );
  mac_control_bitcnt_105_1900 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_252,
      CE => mac_control_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_bitcnt_105_FFX_RST,
      O => mac_control_bitcnt_105
    );
  mac_control_bitcnt_105_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_105_FFX_RST
    );
  mac_control_bitcnt_108_1901 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_255,
      CE => mac_control_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_bitcnt_107_FFY_RST,
      O => mac_control_bitcnt_108
    );
  mac_control_bitcnt_107_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_107_FFY_RST
    );
  rx_input_memio_MD_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(23),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_23_FFX_RST,
      O => d1(23)
    );
  d1_23_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_23_FFX_RST
    );
  rx_input_memio_MD_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_15_FFX_RST,
      O => d1(15)
    );
  d1_15_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_15_FFX_RST
    );
  rx_input_memio_MD_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(25),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_25_FFX_RST,
      O => d1(25)
    );
  d1_25_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_25_FFX_RST
    );
  rx_input_memio_MD_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(24),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_25_FFY_RST,
      O => d1(24)
    );
  d1_25_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_25_FFY_RST
    );
  rx_input_memio_MD_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(16),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_17_FFY_RST,
      O => d1(16)
    );
  d1_17_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_17_FFY_RST
    );
  rx_input_memio_MD_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(17),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_17_FFX_RST,
      O => d1(17)
    );
  d1_17_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_17_FFX_RST
    );
  rx_input_memio_MD_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(26),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_27_FFY_RST,
      O => d1(26)
    );
  d1_27_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_27_FFY_RST
    );
  rx_input_memio_MD_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(27),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_27_FFX_RST,
      O => d1(27)
    );
  d1_27_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_27_FFX_RST
    );
  rx_input_memio_MD_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(18),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_19_FFY_RST,
      O => d1(18)
    );
  d1_19_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_19_FFY_RST
    );
  rx_input_memio_cs_FFd12_1902 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd12_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd12_FFX_RST,
      O => rx_input_memio_cs_FFd12
    );
  rx_input_memio_cs_FFd12_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd12_FFX_RST
    );
  rx_input_memio_cs_FFd14_1903 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd14_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd14_FFX_RST,
      O => rx_input_memio_cs_FFd14
    );
  rx_input_memio_cs_FFd14_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd14_FFX_RST
    );
  mac_control_rxoferr_rst_1904 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0067,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_rxfifowerr_rst_FFY_RST,
      O => mac_control_rxoferr_rst
    );
  mac_control_rxfifowerr_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_rst_FFY_RST
    );
  mac_control_rxfifowerr_rst_1905 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0065,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_rxfifowerr_rst_FFX_RST,
      O => mac_control_rxfifowerr_rst
    );
  mac_control_rxfifowerr_rst_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_rst_FFX_RST
    );
  rx_input_memio_MA_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_11_FFY_RST,
      O => addr1ext(10)
    );
  addr1ext_11_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_11_FFY_RST
    );
  rx_input_memio_menl_1906 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_menl_FROM,
      CE => rx_input_memio_menl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_menl_FFX_RST,
      O => rx_input_memio_menl
    );
  rx_input_memio_menl_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_menl_FFX_RST
    );
  rx_input_memio_MA_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_11_FFX_RST,
      O => addr1ext(11)
    );
  addr1ext_11_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_11_FFX_RST
    );
  rx_input_memio_MA_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_13_FFX_RST,
      O => addr1ext(13)
    );
  addr1ext_13_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_13_FFX_RST
    );
  rx_input_memio_MA_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_13_FFY_RST,
      O => addr1ext(12)
    );
  addr1ext_13_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_13_FFY_RST
    );
  rx_input_memio_MA_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_15_FFY_RST,
      O => addr1ext(14)
    );
  addr1ext_15_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_15_FFY_RST
    );
  mac_control_PHY_status_cs_FFd1_1907 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd1_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd2_FFY_RST,
      O => mac_control_PHY_status_cs_FFd1
    );
  mac_control_PHY_status_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd2_FFY_RST
    );
  mac_control_PHY_status_cs_FFd2_1908 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd2_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd2_FFX_RST,
      O => mac_control_PHY_status_cs_FFd2
    );
  mac_control_PHY_status_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd2_FFX_RST
    );
  mac_control_PHY_status_cs_FFd3_1909 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd3_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd4_FFY_RST,
      O => mac_control_PHY_status_cs_FFd3
    );
  mac_control_PHY_status_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd4_FFY_RST
    );
  mac_control_PHY_status_cs_FFd4_1910 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd4_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd4_FFX_RST,
      O => mac_control_PHY_status_cs_FFd4
    );
  mac_control_PHY_status_cs_FFd4_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd4_FFX_RST
    );
  mac_control_PHY_status_cs_FFd5_1911 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd5_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd6_FFY_RST,
      O => mac_control_PHY_status_cs_FFd5
    );
  mac_control_PHY_status_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd6_FFY_RST
    );
  mac_control_PHY_status_cs_FFd6_1912 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd6_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd6_FFX_RST,
      O => mac_control_PHY_status_cs_FFd6
    );
  mac_control_PHY_status_cs_FFd6_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd6_FFX_RST
    );
  mac_control_PHY_status_cs_FFd7_1913 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd7_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd8_FFY_RST,
      O => mac_control_PHY_status_cs_FFd7
    );
  mac_control_PHY_status_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd8_FFY_RST
    );
  slowclock_clkcnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_clkcnt_n0000(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => slowclock_n0002,
      O => slowclock_clkcnt(2)
    );
  mac_control_PHY_status_cs_FFd8_1914 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd8_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => mac_control_PHY_status_cs_FFd8_FFX_SET,
      RST => GND,
      O => mac_control_PHY_status_cs_FFd8
    );
  mac_control_PHY_status_cs_FFd8_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => mac_control_PHY_status_cs_FFd8_FFX_SET
    );
  tx_output_crcsell_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd2,
      CE => tx_output_crcsell_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcsell_1_FFX_RST,
      O => tx_output_crcsell(1)
    );
  tx_output_crcsell_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcsell_1_FFX_RST
    );
  mac_control_bitcnt_107_1915 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_254,
      CE => mac_control_n0016,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_bitcnt_107_FFX_RST,
      O => mac_control_bitcnt_107
    );
  mac_control_bitcnt_107_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_107_FFX_RST
    );
  mac_control_txfifowerr_rst_1916 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0064,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_rxf_rst_FFY_RST,
      O => mac_control_txfifowerr_rst
    );
  mac_control_rxf_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_rst_FFY_RST
    );
  mac_control_rxf_rst_1917 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0063,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_rxf_rst_FFX_RST,
      O => mac_control_rxf_rst
    );
  mac_control_rxf_rst_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_rst_FFX_RST
    );
  rx_input_memio_addrchk_cs_FFd3_1918 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd4_FFY_RST,
      O => rx_input_memio_addrchk_cs_FFd3
    );
  rx_input_memio_addrchk_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd4_FFY_RST
    );
  rx_input_memio_addrchk_cs_FFd4_1919 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd4_FFX_RST,
      O => rx_input_memio_addrchk_cs_FFd4
    );
  rx_input_memio_addrchk_cs_FFd4_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd4_FFX_RST
    );
  rx_input_memio_cs_FFd9_1920 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd9_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd10_FFY_RST,
      O => rx_input_memio_cs_FFd9
    );
  rx_input_memio_cs_FFd10_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd10_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(2),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_3_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(2)
    );
  mac_control_PHY_status_MII_Interface_statecnt_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_3_FFY_RST
    );
  rx_input_memio_cs_FFd10_1921 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd10_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd10_FFX_RST,
      O => rx_input_memio_cs_FFd10
    );
  rx_input_memio_cs_FFd10_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd10_FFX_RST
    );
  tx_input_den_1922 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_lden,
      CE => tx_input_den_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_den_FFY_RST,
      O => tx_input_den
    );
  tx_input_den_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_den_FFY_RST
    );
  tx_input_CNT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(0),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_1_FFY_RST,
      O => tx_input_CNT(0)
    );
  tx_input_CNT_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_1_FFY_RST
    );
  tx_input_CNT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(1),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_1_FFX_RST,
      O => tx_input_CNT(1)
    );
  tx_input_CNT_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_1_FFX_RST
    );
  tx_input_CNT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(3),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_3_FFX_RST,
      O => tx_input_CNT(3)
    );
  tx_input_CNT_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_3_FFX_RST
    );
  tx_input_CNT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(2),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_3_FFY_RST,
      O => tx_input_CNT(2)
    );
  tx_input_CNT_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_3_FFY_RST
    );
  tx_input_CNT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(5),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_5_FFX_RST,
      O => tx_input_CNT(5)
    );
  tx_input_CNT_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_5_FFX_RST
    );
  tx_input_CNT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(4),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_5_FFY_RST,
      O => tx_input_CNT(4)
    );
  tx_input_CNT_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_5_FFY_RST
    );
  tx_input_CNT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(7),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_7_FFX_RST,
      O => tx_input_CNT(7)
    );
  tx_input_CNT_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_7_FFX_RST
    );
  tx_input_CNT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(6),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_7_FFY_RST,
      O => tx_input_CNT(6)
    );
  tx_input_CNT_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_7_FFY_RST
    );
  tx_input_CNT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(8),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_9_FFY_RST,
      O => tx_input_CNT(8)
    );
  tx_input_CNT_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_9_FFY_RST
    );
  rx_input_memio_MD_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_5_FFX_RST,
      O => d1(5)
    );
  d1_5_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_5_FFX_RST
    );
  rx_input_memio_MD_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_7_FFX_RST,
      O => d1(7)
    );
  d1_7_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_7_FFX_RST
    );
  rx_input_memio_MD_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_7_FFY_RST,
      O => d1(6)
    );
  d1_7_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_7_FFY_RST
    );
  rx_input_memio_MD_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_9_FFX_RST,
      O => d1(9)
    );
  d1_9_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_9_FFX_RST
    );
  rx_input_memio_MD_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_9_FFY_RST,
      O => d1(8)
    );
  d1_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_9_FFY_RST
    );
  rx_input_memio_crcl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(21),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_21_FFX_RST,
      O => rx_input_memio_crcl(21)
    );
  rx_input_memio_crcl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_21_FFX_RST
    );
  rx_input_memio_crcl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(20),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_21_FFY_RST,
      O => rx_input_memio_crcl(20)
    );
  rx_input_memio_crcl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_21_FFY_RST
    );
  rx_input_memio_crcl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(31),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_31_FFX_RST,
      O => rx_input_memio_crcl(31)
    );
  rx_input_memio_crcl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_31_FFX_RST
    );
  rx_input_memio_cs_FFd13_1923 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd13_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd14_FFY_RST,
      O => rx_input_memio_cs_FFd13
    );
  rx_input_memio_cs_FFd14_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd14_FFY_RST
    );
  rx_input_memio_cs_FFd11_1924 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd11_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd12_FFY_RST,
      O => rx_input_memio_cs_FFd11
    );
  rx_input_memio_cs_FFd12_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd12_FFY_RST
    );
  rx_input_memio_MD_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(19),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_19_FFX_RST,
      O => d1(19)
    );
  d1_19_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_19_FFX_RST
    );
  rx_input_memio_MD_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(28),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_29_FFY_RST,
      O => d1(28)
    );
  d1_29_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_29_FFY_RST
    );
  rx_input_memio_MD_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(29),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_29_FFX_RST,
      O => d1(29)
    );
  d1_29_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_29_FFX_RST
    );
  rx_output_fifodin_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(10),
      CE => rx_output_fifodin_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_11_FFY_RST,
      O => rx_output_fifodin(10)
    );
  rx_output_fifodin_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_11_FFY_RST
    );
  rx_output_fifodin_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(11),
      CE => rx_output_fifodin_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_11_FFX_RST,
      O => rx_output_fifodin(11)
    );
  rx_output_fifodin_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_11_FFX_RST
    );
  rx_output_fifodin_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(12),
      CE => rx_output_fifodin_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_13_FFY_RST,
      O => rx_output_fifodin(12)
    );
  rx_output_fifodin_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_13_FFY_RST
    );
  rx_output_fifodin_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(13),
      CE => rx_output_fifodin_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_13_FFX_RST,
      O => rx_output_fifodin(13)
    );
  rx_output_fifodin_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_13_FFX_RST
    );
  rx_output_fifodin_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(14),
      CE => rx_output_fifodin_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_15_FFY_RST,
      O => rx_output_fifodin(14)
    );
  rx_output_fifodin_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_15_FFY_RST
    );
  rx_output_fifodin_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(15),
      CE => rx_output_fifodin_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_15_FFX_RST,
      O => rx_output_fifodin(15)
    );
  rx_output_fifodin_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_15_FFX_RST
    );
  tx_input_enableintl_1925 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_enableintl_GSHIFT,
      CE => tx_input_enableintl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_enableintl_FFY_RST,
      O => tx_input_enableintl
    );
  tx_input_enableintl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_enableintl_FFY_RST
    );
  rx_input_memio_MA_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_15_FFX_RST,
      O => addr1ext(15)
    );
  addr1ext_15_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_15_FFX_RST
    );
  rx_input_memio_MD_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_11_FFX_RST,
      O => d1(11)
    );
  d1_11_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_11_FFX_RST
    );
  rx_input_memio_MD_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_11_FFY_RST,
      O => d1(10)
    );
  d1_11_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_11_FFY_RST
    );
  rx_input_memio_MD_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(21),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_21_FFX_RST,
      O => d1(21)
    );
  d1_21_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_21_FFX_RST
    );
  rx_input_memio_MD_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(20),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_21_FFY_RST,
      O => d1(20)
    );
  d1_21_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_21_FFY_RST
    );
  rx_input_memio_MD_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_13_FFY_RST,
      O => d1(12)
    );
  d1_13_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_13_FFY_RST
    );
  rx_input_memio_MD_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_13_FFX_RST,
      O => d1(13)
    );
  d1_13_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_13_FFX_RST
    );
  rx_input_memio_MD_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(31),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_31_FFX_RST,
      O => d1(31)
    );
  d1_31_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_31_FFX_RST
    );
  rx_input_memio_MD_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(30),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_31_FFY_RST,
      O => d1(30)
    );
  d1_31_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_31_FFY_RST
    );
  rx_input_memio_MD_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_15_FFY_RST,
      O => d1(14)
    );
  d1_15_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_15_FFY_RST
    );
  rx_input_memio_MD_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(22),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_23_FFY_RST,
      O => d1(22)
    );
  d1_23_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_23_FFY_RST
    );
  mac_control_rxcrcerr_rst_1926 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0068,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_rxcrcerr_rst_FFX_RST,
      O => mac_control_rxcrcerr_rst
    );
  mac_control_rxcrcerr_rst_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_rst_FFX_RST
    );
  mac_control_rxphyerr_rst_1927 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0066,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_rxcrcerr_rst_FFY_RST,
      O => mac_control_rxphyerr_rst
    );
  mac_control_rxcrcerr_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_rst_FFY_RST
    );
  rx_output_fifodin_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(0),
      CE => rx_output_fifodin_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_1_FFY_RST,
      O => rx_output_fifodin(0)
    );
  rx_output_fifodin_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_1_FFY_RST
    );
  rx_output_fifodin_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(1),
      CE => rx_output_fifodin_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_1_FFX_RST,
      O => rx_output_fifodin(1)
    );
  rx_output_fifodin_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_1_FFX_RST
    );
  rx_output_fifodin_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(2),
      CE => rx_output_fifodin_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_3_FFY_RST,
      O => rx_output_fifodin(2)
    );
  rx_output_fifodin_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_3_FFY_RST
    );
  rx_output_fifodin_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(3),
      CE => rx_output_fifodin_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_3_FFX_RST,
      O => rx_output_fifodin(3)
    );
  rx_output_fifodin_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_3_FFX_RST
    );
  rx_output_fifodin_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(4),
      CE => rx_output_fifodin_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_5_FFY_RST,
      O => rx_output_fifodin(4)
    );
  rx_output_fifodin_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_5_FFY_RST
    );
  rx_output_fifodin_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(5),
      CE => rx_output_fifodin_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_5_FFX_RST,
      O => rx_output_fifodin(5)
    );
  rx_output_fifodin_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_5_FFX_RST
    );
  rx_output_fifodin_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(6),
      CE => rx_output_fifodin_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_7_FFY_RST,
      O => rx_output_fifodin(6)
    );
  rx_output_fifodin_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_7_FFY_RST
    );
  rx_output_fifodin_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(7),
      CE => rx_output_fifodin_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_7_FFX_RST,
      O => rx_output_fifodin(7)
    );
  rx_output_fifodin_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_7_FFX_RST
    );
  rx_output_fifodin_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(8),
      CE => rx_output_fifodin_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_9_FFY_RST,
      O => rx_output_fifodin(8)
    );
  rx_output_fifodin_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_9_FFY_RST
    );
  tx_input_dinint_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(11),
      CE => tx_input_dinint_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_11_FFX_RST,
      O => tx_input_dinint(11)
    );
  tx_input_dinint_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_11_FFX_RST
    );
  tx_input_dinint_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(12),
      CE => tx_input_dinint_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_13_FFY_RST,
      O => tx_input_dinint(12)
    );
  tx_input_dinint_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_13_FFY_RST
    );
  tx_input_dinint_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(13),
      CE => tx_input_dinint_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_13_FFX_RST,
      O => tx_input_dinint(13)
    );
  tx_input_dinint_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_13_FFX_RST
    );
  tx_input_dinint_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(14),
      CE => tx_input_dinint_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_15_FFY_RST,
      O => tx_input_dinint(14)
    );
  tx_input_dinint_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_15_FFY_RST
    );
  tx_input_dinint_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(15),
      CE => tx_input_dinint_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_15_FFX_RST,
      O => tx_input_dinint(15)
    );
  tx_input_dinint_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_15_FFX_RST
    );
  rx_input_memio_RXCRCERR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0060,
      CE => rxfifowerr_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfifowerr_FFY_RST,
      O => rxcrcerr
    );
  rxfifowerr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfifowerr_FFY_RST
    );
  rx_input_memio_RXFIFOWERR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0061,
      CE => rxfifowerr_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfifowerr_FFX_RST,
      O => rxfifowerr
    );
  rxfifowerr_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfifowerr_FFX_RST
    );
  rx_output_cs_FFd19_1928 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_cs_FFd19_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_cs_FFd5_FFY_SET,
      RST => GND,
      O => rx_output_cs_FFd19
    );
  rx_output_cs_FFd5_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => rx_output_cs_FFd5_FFY_SET
    );
  tx_input_dinint_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(1),
      CE => tx_input_dinint_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_1_FFX_RST,
      O => tx_input_dinint(1)
    );
  tx_input_dinint_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_1_FFX_RST
    );
  tx_input_dinint_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(2),
      CE => tx_input_dinint_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_3_FFY_RST,
      O => tx_input_dinint(2)
    );
  tx_input_dinint_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_3_FFY_RST
    );
  tx_input_dinint_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(3),
      CE => tx_input_dinint_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_3_FFX_RST,
      O => tx_input_dinint(3)
    );
  tx_input_dinint_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_3_FFX_RST
    );
  tx_input_dinint_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(4),
      CE => tx_input_dinint_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_5_FFY_RST,
      O => tx_input_dinint(4)
    );
  tx_input_dinint_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_5_FFY_RST
    );
  tx_input_dinint_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(5),
      CE => tx_input_dinint_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_5_FFX_RST,
      O => tx_input_dinint(5)
    );
  tx_input_dinint_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_5_FFX_RST
    );
  tx_input_dinint_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(6),
      CE => tx_input_dinint_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_7_FFY_RST,
      O => tx_input_dinint(6)
    );
  tx_input_dinint_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_7_FFY_RST
    );
  tx_input_dinint_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(7),
      CE => tx_input_dinint_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_7_FFX_RST,
      O => tx_input_dinint(7)
    );
  tx_input_dinint_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_7_FFX_RST
    );
  tx_input_dinint_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(8),
      CE => tx_input_dinint_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_9_FFY_RST,
      O => tx_input_dinint(8)
    );
  tx_input_dinint_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_9_FFY_RST
    );
  tx_input_dinint_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(9),
      CE => tx_input_dinint_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_9_FFX_RST,
      O => tx_input_dinint(9)
    );
  tx_input_dinint_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_9_FFX_RST
    );
  mac_control_Mshreg_scslll_103_1929 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_Mshreg_scslll_net187,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_Mshreg_scslll_103_FFY_RST,
      O => mac_control_Mshreg_scslll_103
    );
  mac_control_Mshreg_scslll_103_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_Mshreg_scslll_103_FFY_RST
    );
  memcontroller_dnl2_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(10),
      CE => memcontroller_dnl2_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_11_FFY_RST,
      O => memcontroller_dnl2(10)
    );
  memcontroller_dnl2_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_11_FFY_RST
    );
  memcontroller_dnl2_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(11),
      CE => memcontroller_dnl2_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_11_FFX_RST,
      O => memcontroller_dnl2(11)
    );
  memcontroller_dnl2_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_11_FFX_RST
    );
  memcontroller_dnl2_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(20),
      CE => memcontroller_dnl2_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_21_FFY_RST,
      O => memcontroller_dnl2(20)
    );
  memcontroller_dnl2_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_21_FFY_RST
    );
  memcontroller_dnl2_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(21),
      CE => memcontroller_dnl2_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_21_FFX_RST,
      O => memcontroller_dnl2(21)
    );
  memcontroller_dnl2_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_21_FFX_RST
    );
  memcontroller_dnl2_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(12),
      CE => memcontroller_dnl2_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_13_FFY_RST,
      O => memcontroller_dnl2(12)
    );
  memcontroller_dnl2_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_13_FFY_RST
    );
  memcontroller_dnl2_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(13),
      CE => memcontroller_dnl2_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_13_FFX_RST,
      O => memcontroller_dnl2(13)
    );
  memcontroller_dnl2_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_13_FFX_RST
    );
  memcontroller_dnl2_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(30),
      CE => memcontroller_dnl2_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_31_FFY_RST,
      O => memcontroller_dnl2(30)
    );
  memcontroller_dnl2_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_31_FFY_RST
    );
  memcontroller_dnl2_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(22),
      CE => memcontroller_dnl2_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_23_FFY_RST,
      O => memcontroller_dnl2(22)
    );
  memcontroller_dnl2_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_23_FFY_RST
    );
  rx_output_fifodin_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(9),
      CE => rx_output_fifodin_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_9_FFX_RST,
      O => rx_output_fifodin(9)
    );
  rx_output_fifodin_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_9_FFX_RST
    );
  rx_output_fifo_full_1930 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0051,
      CE => rx_output_fifo_full_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_full_FFY_RST,
      O => rx_output_fifo_full
    );
  rx_output_fifo_full_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifo_full_FFY_RST
    );
  rx_input_GMII_FIFOIN_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_GMII_N80573,
      CE => VCC,
      CLK => clkrx,
      SET => GSR,
      RST => GND,
      SSET => rx_input_GMII_rx_erl,
      SRST => GND,
      O => rx_input_fifoin(0)
    );
  rx_input_GMII_FIFOIN_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_GMII_N80576,
      CE => VCC,
      CLK => clkrx,
      SET => GSR,
      RST => GND,
      SSET => rx_input_GMII_rx_of,
      SRST => GND,
      O => rx_input_fifoin(1)
    );
  rx_input_GMII_FIFOIN_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_GMII_N80579,
      CE => VCC,
      CLK => clkrx,
      SET => GSR,
      RST => GND,
      SSET => rx_input_GMII_rx_of,
      SRST => GND,
      O => rx_input_fifoin(2)
    );
  rx_input_GMII_FIFOIN_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_N80582,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_rx_of,
      O => rx_input_fifoin(3)
    );
  rx_input_GMII_FIFOIN_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_N80570,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_rx_of,
      O => rx_input_fifoin(4)
    );
  rx_input_GMII_FIFOIN_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_N80561,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_rx_of,
      O => rx_input_fifoin(5)
    );
  tx_input_dinint_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(10),
      CE => tx_input_dinint_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_11_FFY_RST,
      O => tx_input_dinint(10)
    );
  tx_input_dinint_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_11_FFY_RST
    );
  rx_input_GMII_FIFOIN_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_N80564,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_rx_of,
      O => rx_input_fifoin(6)
    );
  rx_input_GMII_FIFOIN_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_N80567,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_rx_of,
      O => rx_input_fifoin(7)
    );
  rx_input_memio_RXPHYERR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0057,
      CE => rxoferr_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxoferr_FFY_RST,
      O => rxphyerr
    );
  rxoferr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxoferr_FFY_RST
    );
  rx_output_cs_FFd5_1931 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd5_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd5_FFX_RST,
      O => rx_output_cs_FFd5
    );
  rx_output_cs_FFd5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd5_FFX_RST
    );
  rx_input_memio_RXOFERR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0058,
      CE => rxoferr_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxoferr_FFX_RST,
      O => rxoferr
    );
  rxoferr_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxoferr_FFX_RST
    );
  tx_input_cs_FFd11_1932 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd11_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd11_FFY_RST,
      O => tx_input_cs_FFd11
    );
  tx_input_cs_FFd11_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd11_FFY_RST
    );
  tx_input_CNT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(10),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_11_FFY_RST,
      O => tx_input_CNT(10)
    );
  tx_input_CNT_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_11_FFY_RST
    );
  tx_input_CNT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(11),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_11_FFX_RST,
      O => tx_input_CNT(11)
    );
  tx_input_CNT_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_11_FFX_RST
    );
  tx_input_CNT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(13),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_13_FFX_RST,
      O => tx_input_CNT(13)
    );
  tx_input_CNT_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_13_FFX_RST
    );
  tx_input_CNT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(12),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_13_FFY_RST,
      O => tx_input_CNT(12)
    );
  tx_input_CNT_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_13_FFY_RST
    );
  tx_input_CNT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(15),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_15_FFX_RST,
      O => tx_input_CNT(15)
    );
  tx_input_CNT_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_15_FFX_RST
    );
  tx_input_CNT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(14),
      CE => tx_input_N34493,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_15_FFY_RST,
      O => tx_input_CNT(14)
    );
  tx_input_CNT_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_15_FFY_RST
    );
  tx_input_dinint_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(0),
      CE => tx_input_dinint_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_1_FFY_RST,
      O => tx_input_dinint(0)
    );
  tx_input_dinint_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_1_FFY_RST
    );
  tx_output_crcl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(19),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_19_FFY_RST,
      O => tx_output_crcl(19)
    );
  tx_output_crcl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_19_FFY_RST
    );
  mac_control_dout_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N76337,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_0_FFY_RST,
      O => mac_control_dout(0)
    );
  mac_control_dout_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_0_FFY_RST
    );
  rx_input_fifo_control_cs_FFd1_1933 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_cs_FFd1_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_cs_FFd2_FFY_RST,
      O => rx_input_fifo_control_cs_FFd1
    );
  rx_input_fifo_control_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_cs_FFd2_FFY_RST
    );
  rx_input_fifo_control_cs_FFd2_1934 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_cs_FFd2_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_cs_FFd2_FFX_RST,
      O => rx_input_fifo_control_cs_FFd2
    );
  rx_input_fifo_control_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_cs_FFd2_FFX_RST
    );
  rx_input_fifo_control_cs_FFd3_1935 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_cs_FFd4_FFY_RST,
      O => rx_input_fifo_control_cs_FFd3
    );
  rx_input_fifo_control_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_cs_FFd4_FFY_RST
    );
  rx_input_fifo_control_cs_FFd4_1936 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_control_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_control_cs_FFd4_FFX_SET,
      RST => GND,
      O => rx_input_fifo_control_cs_FFd4
    );
  rx_input_fifo_control_cs_FFd4_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF_2,
      O => rx_input_fifo_control_cs_FFd4_FFX_SET
    );
  rx_output_cs_FFd1_1937 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd1_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd2_FFY_RST,
      O => rx_output_cs_FFd1
    );
  rx_output_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd2_FFY_RST
    );
  rx_output_cs_FFd2_1938 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd2_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd2_FFX_RST,
      O => rx_output_cs_FFd2
    );
  rx_output_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd2_FFX_RST
    );
  rx_output_cs_FFd3_1939 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd4_FFY_RST,
      O => rx_output_cs_FFd3
    );
  rx_output_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd4_FFY_RST
    );
  rx_output_cs_FFd4_1940 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd4_FFX_RST,
      O => rx_output_cs_FFd4
    );
  rx_output_cs_FFd4_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd4_FFX_RST
    );
  rx_output_cs_FFd7_1941 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd7_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd8_FFY_RST,
      O => rx_output_cs_FFd7
    );
  rx_output_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd8_FFY_RST
    );
  rx_output_fifo_BU458 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3969,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1593_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1592
    );
  rx_output_fifo_N1593_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1593_FFY_SET
    );
  rx_output_fifo_BU456 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3968,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1593_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1593
    );
  rx_output_fifo_N1593_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1593_FFX_SET
    );
  tx_output_cs_FFd6_1942 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd6_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd6_FFX_RST,
      O => tx_output_cs_FFd6
    );
  tx_output_cs_FFd6_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd6_FFX_RST
    );
  tx_output_cs_FFd5_1943 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd5_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd6_FFY_RST,
      O => tx_output_cs_FFd5
    );
  tx_output_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd6_FFY_RST
    );
  tx_output_cs_FFd7_1944 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd7_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd8_FFY_RST,
      O => tx_output_cs_FFd7
    );
  tx_output_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd8_FFY_RST
    );
  tx_output_cs_FFd8_1945 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd8_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd8_FFX_RST,
      O => tx_output_cs_FFd8
    );
  tx_output_cs_FFd8_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => tx_output_cs_FFd8_FFX_RST
    );
  rx_input_memio_Mshreg_lbpout4_0_69_1946 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_0_net34,
      CE => rx_input_memio_Mshreg_lbpout4_0_69_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_0_69_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_0_69
    );
  rx_input_memio_Mshreg_lbpout4_0_69_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_0_69_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_1_68_1947 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_1_net32,
      CE => rx_input_memio_Mshreg_lbpout4_1_68_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_1_68_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_1_68
    );
  rx_input_memio_Mshreg_lbpout4_1_68_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_1_68_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_2_67_1948 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_2_net30,
      CE => rx_input_memio_Mshreg_lbpout4_2_67_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_2_67_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_2_67
    );
  rx_input_memio_Mshreg_lbpout4_2_67_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_2_67_FFY_RST
    );
  rx_input_memio_crcl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(9),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_9_FFY_RST,
      O => rx_input_memio_crcl(9)
    );
  rx_input_memio_crcl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_9_FFY_RST
    );
  mac_control_sclkdeltall_1949 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_sclkdeltal,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_sclkdeltall_FFY_RST,
      O => mac_control_sclkdeltall
    );
  mac_control_sclkdeltall_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_sclkdeltall_FFY_RST
    );
  mac_control_phyaddr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_11_FFY_RST,
      O => mac_control_phyaddr(10)
    );
  mac_control_phyaddr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_11_FFY_RST
    );
  mac_control_phyaddr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_11_FFX_RST,
      O => mac_control_phyaddr(11)
    );
  mac_control_phyaddr_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_11_FFX_RST
    );
  mac_control_phyaddr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_13_FFY_RST,
      O => mac_control_phyaddr(12)
    );
  mac_control_phyaddr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_13_FFY_RST
    );
  mac_control_phyaddr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_13_FFX_RST,
      O => mac_control_phyaddr(13)
    );
  mac_control_phyaddr_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_13_FFX_RST
    );
  mac_control_phyaddr_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(20),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_21_FFY_RST,
      O => mac_control_phyaddr(20)
    );
  mac_control_phyaddr_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_21_FFY_RST
    );
  mac_control_phyaddr_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(21),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_21_FFX_RST,
      O => mac_control_phyaddr(21)
    );
  mac_control_phyaddr_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_21_FFX_RST
    );
  mac_control_phyaddr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_15_FFY_RST,
      O => mac_control_phyaddr(14)
    );
  mac_control_phyaddr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_15_FFY_RST
    );
  mac_control_phyaddr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_15_FFX_RST,
      O => mac_control_phyaddr(15)
    );
  mac_control_phyaddr_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_15_FFX_RST
    );
  mac_control_phyaddr_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(22),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_23_FFY_RST,
      O => mac_control_phyaddr(22)
    );
  mac_control_phyaddr_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_23_FFY_RST
    );
  mac_control_phyaddr_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(23),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_23_FFX_RST,
      O => mac_control_phyaddr(23)
    );
  mac_control_phyaddr_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_23_FFX_RST
    );
  mac_control_phyaddr_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(30),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_30_FFY_RST,
      O => mac_control_phyaddr(30)
    );
  mac_control_phyaddr_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_30_FFY_RST
    );
  mac_control_phyaddr_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(16),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_17_FFY_RST,
      O => mac_control_phyaddr(16)
    );
  mac_control_phyaddr_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_17_FFY_RST
    );
  rx_output_cs_FFd8_1950 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd8_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd8_FFX_RST,
      O => rx_output_cs_FFd8
    );
  rx_output_cs_FFd8_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd8_FFX_RST
    );
  tx_input_cs_FFd2_1951 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd2_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd4_FFY_RST,
      O => tx_input_cs_FFd2
    );
  tx_input_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd4_FFY_RST
    );
  tx_input_cs_FFd3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfifowerr_FFY_RST,
      O => txfifowerr
    );
  txfifowerr_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => txfifowerr_FFY_RST
    );
  tx_input_cs_FFd4_1952 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd8,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd4_FFX_RST,
      O => tx_input_cs_FFd4
    );
  tx_input_cs_FFd4_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd4_FFX_RST
    );
  tx_input_cs_FFd7_1953 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd7_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd8_FFY_RST,
      O => tx_input_cs_FFd7
    );
  tx_input_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd8_FFY_RST
    );
  tx_input_cs_FFd8_1954 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd8_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd8_FFX_RST,
      O => tx_input_cs_FFd8
    );
  tx_input_cs_FFd8_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd8_FFX_RST
    );
  tx_input_cs_FFd9_1955 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd9_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd9_FFY_RST,
      O => tx_input_cs_FFd9
    );
  tx_input_cs_FFd9_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd9_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_10_59_1956 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_10_net14,
      CE => rx_input_memio_Mshreg_lbpout4_10_59_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_10_59_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_10_59
    );
  rx_input_memio_Mshreg_lbpout4_10_59_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_10_59_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_12_57_1957 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_12_net10,
      CE => rx_input_memio_Mshreg_lbpout4_12_57_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_12_57_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_12_57
    );
  rx_input_memio_Mshreg_lbpout4_12_57_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_12_57_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_11_58_1958 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_11_net12,
      CE => rx_input_memio_Mshreg_lbpout4_11_58_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_11_58_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_11_58
    );
  rx_input_memio_Mshreg_lbpout4_11_58_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_11_58_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_13_56_1959 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_13_net8,
      CE => rx_input_memio_Mshreg_lbpout4_13_56_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_13_56_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_13_56
    );
  rx_input_memio_Mshreg_lbpout4_13_56_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_13_56_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_14_55_1960 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_14_net6,
      CE => rx_input_memio_Mshreg_lbpout4_14_55_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_14_55_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_14_55
    );
  rx_input_memio_Mshreg_lbpout4_14_55_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_14_55_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_15_54_1961 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_15_net4,
      CE => rx_input_memio_Mshreg_lbpout4_15_54_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_15_54_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_15_54
    );
  rx_input_memio_Mshreg_lbpout4_15_54_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_15_54_FFY_RST
    );
  mac_control_Mshreg_sinlll_102_1962 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_Mshreg_sinlll_net185,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_Mshreg_sinlll_102_FFY_RST,
      O => mac_control_Mshreg_sinlll_102
    );
  mac_control_Mshreg_sinlll_102_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_Mshreg_sinlll_102_FFY_RST
    );
  mac_control_PHY_status_PHYADDRSTATUS : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr_31_FROM,
      CE => mac_control_PHY_status_n0017,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_31_FFX_RST,
      O => mac_control_phyaddr(31)
    );
  mac_control_phyaddr_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_31_FFX_RST
    );
  rx_output_fifo_BU105 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2339,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1551_FFX_RST,
      O => rx_output_fifo_N1551
    );
  rx_output_fifo_N1551_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1551_FFX_RST
    );
  rx_output_fifo_BU273 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3307,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1615_FFY_RST,
      O => rx_output_fifo_N1614
    );
  rx_output_fifo_N1615_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1615_FFY_RST
    );
  rx_output_fifo_BU126 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2459,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1549_FFY_RST,
      O => rx_output_fifo_N1548
    );
  rx_output_fifo_N1549_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1549_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_3_66_1963 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_3_net28,
      CE => rx_input_memio_Mshreg_lbpout4_3_66_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_3_66_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_3_66
    );
  rx_input_memio_Mshreg_lbpout4_3_66_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_3_66_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_4_65_1964 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_4_net26,
      CE => rx_input_memio_Mshreg_lbpout4_4_65_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_4_65_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_4_65
    );
  rx_input_memio_Mshreg_lbpout4_4_65_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_4_65_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_5_64_1965 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_5_net24,
      CE => rx_input_memio_Mshreg_lbpout4_5_64_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_5_64_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_5_64
    );
  rx_input_memio_Mshreg_lbpout4_5_64_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_5_64_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_6_63_1966 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_6_net22,
      CE => rx_input_memio_Mshreg_lbpout4_6_63_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_6_63_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_6_63
    );
  rx_input_memio_Mshreg_lbpout4_6_63_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_6_63_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_7_62_1967 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_7_net20,
      CE => rx_input_memio_Mshreg_lbpout4_7_62_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_7_62_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_7_62
    );
  rx_input_memio_Mshreg_lbpout4_7_62_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_7_62_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_8_61_1968 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_8_net18,
      CE => rx_input_memio_Mshreg_lbpout4_8_61_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_8_61_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_8_61
    );
  rx_input_memio_Mshreg_lbpout4_8_61_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_8_61_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_9_60_1969 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_9_net16,
      CE => rx_input_memio_Mshreg_lbpout4_9_60_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_9_60_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_9_60
    );
  rx_input_memio_Mshreg_lbpout4_9_60_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_9_60_FFY_RST
    );
  rx_output_fifo_BU119 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2419,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1549_FFX_RST,
      O => rx_output_fifo_N1549
    );
  rx_output_fifo_N1549_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1549_FFX_RST
    );
  rx_output_fifo_BU266 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3267,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1615_FFX_RST,
      O => rx_output_fifo_N1615
    );
  rx_output_fifo_N1615_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1615_FFX_RST
    );
  rx_output_fifo_BU259 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3227,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1617_FFY_RST,
      O => rx_output_fifo_N1616
    );
  rx_output_fifo_N1617_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1617_FFY_RST
    );
  rx_output_fifo_BU252 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3187,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1617_FFX_RST,
      O => rx_output_fifo_N1617
    );
  rx_output_fifo_N1617_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1617_FFX_RST
    );
  rx_output_fifo_BU287 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3387,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1613_FFY_RST,
      O => rx_output_fifo_N1612
    );
  rx_output_fifo_N1613_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1613_FFY_RST
    );
  rx_output_fifo_BU280 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3347,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1613_FFX_RST,
      O => rx_output_fifo_N1613
    );
  rx_output_fifo_N1613_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1613_FFX_RST
    );
  rx_output_fifo_BU462 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3971,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1589_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1590
    );
  rx_output_fifo_N1589_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1589_FFY_SET
    );
  rx_output_fifo_BU466 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3973,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1588_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1588
    );
  rx_output_fifo_N1588_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1588_FFY_SET
    );
  rx_output_fifo_BU464 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1589_FROM,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1589_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1589
    );
  rx_output_fifo_N1589_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1589_FFX_SET
    );
  tx_output_crcl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(20),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_21_FFY_RST,
      O => tx_output_crcl(20)
    );
  tx_output_crcl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_21_FFY_RST
    );
  tx_input_newfint_1970 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_lnewfint,
      CE => tx_input_newfint_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_newfint_FFY_RST,
      O => tx_input_newfint
    );
  tx_input_newfint_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_newfint_FFY_RST
    );
  tx_output_crcl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(21),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_21_FFX_RST,
      O => tx_output_crcl(21)
    );
  tx_output_crcl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_21_FFX_RST
    );
  tx_output_crcl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(22),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_22_FFY_RST,
      O => tx_output_crcl(22)
    );
  tx_output_crcl_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_22_FFY_RST
    );
  mac_control_dout_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N79864,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_11_FFY_RST,
      O => mac_control_dout(11)
    );
  mac_control_dout_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_11_FFY_RST
    );
  mac_control_phyaddr_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(17),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_17_FFX_RST,
      O => mac_control_phyaddr(17)
    );
  mac_control_phyaddr_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_17_FFX_RST
    );
  mac_control_phyaddr_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(24),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_25_FFY_RST,
      O => mac_control_phyaddr(24)
    );
  mac_control_phyaddr_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_25_FFY_RST
    );
  mac_control_phyaddr_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(25),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_25_FFX_RST,
      O => mac_control_phyaddr(25)
    );
  mac_control_phyaddr_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_25_FFX_RST
    );
  mac_control_phyaddr_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(18),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_19_FFY_RST,
      O => mac_control_phyaddr(18)
    );
  mac_control_phyaddr_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_19_FFY_RST
    );
  mac_control_phyaddr_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(19),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_19_FFX_RST,
      O => mac_control_phyaddr(19)
    );
  mac_control_phyaddr_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_19_FFX_RST
    );
  mac_control_phyaddr_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(26),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_27_FFY_RST,
      O => mac_control_phyaddr(26)
    );
  mac_control_phyaddr_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_27_FFY_RST
    );
  mac_control_phyaddr_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(27),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_27_FFX_RST,
      O => mac_control_phyaddr(27)
    );
  mac_control_phyaddr_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_27_FFX_RST
    );
  mac_control_phyaddr_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(28),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_29_FFY_RST,
      O => mac_control_phyaddr(28)
    );
  mac_control_phyaddr_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_29_FFY_RST
    );
  mac_control_phyaddr_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(29),
      CE => mac_control_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_29_FFX_RST,
      O => mac_control_phyaddr(29)
    );
  mac_control_phyaddr_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_29_FFX_RST
    );
  rx_input_memio_addrchk_datal_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_11_FFY_RST,
      O => rx_input_memio_addrchk_datal(10)
    );
  rx_input_memio_addrchk_datal_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_11_FFY_RST
    );
  rx_input_memio_addrchk_datal_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_11_FFX_RST,
      O => rx_input_memio_addrchk_datal(11)
    );
  rx_input_memio_addrchk_datal_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_11_FFX_RST
    );
  rx_input_memio_addrchk_datal_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_13_FFY_RST,
      O => rx_input_memio_addrchk_datal(12)
    );
  rx_input_memio_addrchk_datal_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_13_FFY_RST
    );
  rx_input_memio_addrchk_datal_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_21_FFY_RST,
      O => rx_input_memio_addrchk_datal(20)
    );
  rx_input_memio_addrchk_datal_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_21_FFY_RST
    );
  rx_input_memio_addrchk_datal_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_21_FFX_RST,
      O => rx_input_memio_addrchk_datal(21)
    );
  rx_input_memio_addrchk_datal_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_21_FFX_RST
    );
  rx_input_memio_addrchk_datal_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_31_FFY_RST,
      O => rx_input_memio_addrchk_datal(30)
    );
  rx_input_memio_addrchk_datal_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_31_FFY_RST
    );
  rx_fifocheck_fbbpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_15_FFX_RST,
      O => rx_fifocheck_fbbpl(15)
    );
  rx_fifocheck_fbbpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_15_FFX_RST
    );
  rx_input_memio_dout_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_11_FFY_RST,
      O => rx_input_memio_dout(10)
    );
  rx_input_memio_dout_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_11_FFY_RST
    );
  rx_input_memio_dout_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_11_FFX_RST,
      O => rx_input_memio_dout(11)
    );
  rx_input_memio_dout_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_11_FFX_RST
    );
  rx_input_memio_dout_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_21_FFX_RST,
      O => rx_input_memio_dout(21)
    );
  rx_input_memio_dout_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_21_FFX_RST
    );
  rx_input_memio_dout_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_13_FFX_RST,
      O => rx_input_memio_dout(13)
    );
  rx_input_memio_dout_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_13_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(11),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_12_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(12)
    );
  mac_control_PHY_status_MII_Interface_dreg_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_12_FFX_RST
    );
  rx_input_memio_dout_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_31_FFY_RST,
      O => rx_input_memio_dout(30)
    );
  rx_input_memio_dout_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_31_FFY_RST
    );
  rx_input_memio_dout_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_31_FFX_RST,
      O => rx_input_memio_dout(31)
    );
  rx_input_memio_dout_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_31_FFX_RST
    );
  rx_input_memio_dout_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_23_FFX_RST,
      O => rx_input_memio_dout(23)
    );
  rx_input_memio_dout_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_23_FFX_RST
    );
  rx_input_memio_dout_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_15_FFX_RST,
      O => rx_input_memio_dout(15)
    );
  rx_input_memio_dout_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_15_FFX_RST
    );
  rx_fifocheck_bpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_9_FFX_RST,
      O => rx_fifocheck_bpl(9)
    );
  rx_fifocheck_bpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_9_FFX_RST
    );
  mac_control_dout_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N78899,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_12_FFY_RST,
      O => mac_control_dout(12)
    );
  mac_control_dout_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_12_FFY_RST
    );
  rx_fifocheck_bpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_1_FFY_RST,
      O => rx_fifocheck_bpl(0)
    );
  rx_fifocheck_bpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_1_FFY_RST
    );
  rx_fifocheck_bpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_1_FFX_RST,
      O => rx_fifocheck_bpl(1)
    );
  rx_fifocheck_bpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_1_FFX_RST
    );
  rx_fifocheck_bpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_3_FFY_RST,
      O => rx_fifocheck_bpl(2)
    );
  rx_fifocheck_bpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_3_FFY_RST
    );
  rx_fifocheck_bpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_3_FFX_RST,
      O => rx_fifocheck_bpl(3)
    );
  rx_fifocheck_bpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_3_FFX_RST
    );
  rx_input_memio_crcll_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(1),
      CE => rx_input_memio_crcll_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_1_FFX_RST,
      O => rx_input_memio_crcll(1)
    );
  rx_input_memio_crcll_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_1_FFX_RST
    );
  rx_input_memio_crcll_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(2),
      CE => rx_input_memio_crcll_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_3_FFY_RST,
      O => rx_input_memio_crcll(2)
    );
  rx_input_memio_crcll_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_3_FFY_RST
    );
  rx_input_memio_crcll_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(3),
      CE => rx_input_memio_crcll_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_3_FFX_RST,
      O => rx_input_memio_crcll(3)
    );
  rx_input_memio_crcll_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_3_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(0),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_1_FFY_RST,
      O => mac_control_phystat(0)
    );
  mac_control_phystat_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_1_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(1),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_1_FFX_RST,
      O => mac_control_phystat(1)
    );
  mac_control_phystat_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_1_FFX_RST
    );
  rx_input_memio_crcll_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(4),
      CE => rx_input_memio_crcll_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_5_FFY_RST,
      O => rx_input_memio_crcll(4)
    );
  rx_input_memio_crcll_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_5_FFY_RST
    );
  rx_input_memio_crcll_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(5),
      CE => rx_input_memio_crcll_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_5_FFX_RST,
      O => rx_input_memio_crcll(5)
    );
  rx_input_memio_crcll_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_5_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(2),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_3_FFY_RST,
      O => mac_control_phystat(2)
    );
  mac_control_phystat_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_3_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(3),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_3_FFX_RST,
      O => mac_control_phystat(3)
    );
  mac_control_phystat_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_3_FFX_RST
    );
  rx_input_memio_crcll_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(6),
      CE => rx_input_memio_crcll_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_7_FFY_RST,
      O => rx_input_memio_crcll(6)
    );
  rx_input_memio_crcll_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_7_FFY_RST
    );
  rx_input_memio_crcll_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(7),
      CE => rx_input_memio_crcll_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_7_FFX_RST,
      O => rx_input_memio_crcll(7)
    );
  rx_input_memio_crcll_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_7_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(4),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_5_FFY_RST,
      O => mac_control_phystat(4)
    );
  mac_control_phystat_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_5_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(5),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_5_FFX_RST,
      O => mac_control_phystat(5)
    );
  mac_control_phystat_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_5_FFX_RST
    );
  rx_input_memio_crcll_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(8),
      CE => rx_input_memio_crcll_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_9_FFY_RST,
      O => rx_input_memio_crcll(8)
    );
  rx_input_memio_crcll_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_9_FFY_RST
    );
  mac_control_dout_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N75776,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_16_FFY_RST,
      O => mac_control_dout(16)
    );
  mac_control_dout_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_16_FFY_RST
    );
  mac_control_dout_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N76142,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_24_FFY_RST,
      O => mac_control_dout(24)
    );
  mac_control_dout_24_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_24_FFY_RST
    );
  mac_control_dout_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N75186,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_25_FFY_RST,
      O => mac_control_dout(25)
    );
  mac_control_dout_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_25_FFY_RST
    );
  mac_control_dout_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N75898,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_17_FFY_RST,
      O => mac_control_dout(17)
    );
  mac_control_dout_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_17_FFY_RST
    );
  mac_control_dout_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N74835,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_18_FFY_RST,
      O => mac_control_dout(18)
    );
  mac_control_dout_18_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_18_FFY_RST
    );
  mac_control_dout_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N75303,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_26_FFY_RST,
      O => mac_control_dout(26)
    );
  mac_control_dout_26_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_26_FFY_RST
    );
  mac_control_dout_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N74952,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_20_FFY_RST,
      O => mac_control_dout(20)
    );
  mac_control_dout_20_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_20_FFY_RST
    );
  rx_fifocheck_bpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_5_FFY_RST,
      O => rx_fifocheck_bpl(4)
    );
  rx_fifocheck_bpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_5_FFY_RST
    );
  rx_fifocheck_bpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_5_FFX_RST,
      O => rx_fifocheck_bpl(5)
    );
  rx_fifocheck_bpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_5_FFX_RST
    );
  rx_fifocheck_bpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_7_FFY_RST,
      O => rx_fifocheck_bpl(6)
    );
  rx_fifocheck_bpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_7_FFY_RST
    );
  rx_fifocheck_bpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_7_FFX_RST,
      O => rx_fifocheck_bpl(7)
    );
  rx_fifocheck_bpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_7_FFX_RST
    );
  rx_fifocheck_bpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_9_FFY_RST,
      O => rx_fifocheck_bpl(8)
    );
  rx_fifocheck_bpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_9_FFY_RST
    );
  mac_control_dout_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N76020,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_21_FFY_RST,
      O => mac_control_dout(21)
    );
  mac_control_dout_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_21_FFY_RST
    );
  mac_control_dout_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N75537,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_30_FFY_RST,
      O => mac_control_dout(30)
    );
  mac_control_dout_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_30_FFY_RST
    );
  mac_control_dout_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N75069,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_22_FFY_RST,
      O => mac_control_dout(22)
    );
  mac_control_dout_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_22_FFY_RST
    );
  mac_control_dout_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N80026,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_15_FFY_RST,
      O => mac_control_dout(15)
    );
  mac_control_dout_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_15_FFY_RST
    );
  mac_control_dout_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N79056,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_13_FFY_RST,
      O => mac_control_dout(13)
    );
  mac_control_dout_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_13_FFY_RST
    );
  tx_output_crcl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(13),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_13_FFY_RST,
      O => tx_output_crcl(13)
    );
  tx_output_crcl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_13_FFY_RST
    );
  mac_control_phydi_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(19),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_19_FFX_RST,
      O => mac_control_phydi(19)
    );
  mac_control_phydi_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_19_FFX_RST
    );
  mac_control_phydi_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(26),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_27_FFY_RST,
      O => mac_control_phydi(26)
    );
  mac_control_phydi_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_27_FFY_RST
    );
  mac_control_phydi_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(27),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_27_FFX_RST,
      O => mac_control_phydi(27)
    );
  mac_control_phydi_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_27_FFX_RST
    );
  mac_control_phydi_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(28),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_29_FFY_RST,
      O => mac_control_phydi(28)
    );
  mac_control_phydi_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_29_FFY_RST
    );
  mac_control_phydi_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(29),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_29_FFX_RST,
      O => mac_control_phydi(29)
    );
  mac_control_phydi_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_29_FFX_RST
    );
  rx_input_memio_bpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(0),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_1_FFY_RST,
      O => rx_input_memio_bpl(0)
    );
  rx_input_memio_bpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_1_FFY_RST
    );
  rx_input_memio_bpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(1),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_1_FFX_RST,
      O => rx_input_memio_bpl(1)
    );
  rx_input_memio_bpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_1_FFX_RST
    );
  rx_input_memio_bpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(2),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_3_FFY_RST,
      O => rx_input_memio_bpl(2)
    );
  rx_input_memio_bpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_3_FFY_RST
    );
  rx_input_memio_bpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(3),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_3_FFX_RST,
      O => rx_input_memio_bpl(3)
    );
  rx_input_memio_bpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_3_FFX_RST
    );
  rx_input_memio_bpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(4),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_5_FFY_RST,
      O => rx_input_memio_bpl(4)
    );
  rx_input_memio_bpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_5_FFY_RST
    );
  rx_input_memio_bpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(5),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_5_FFX_RST,
      O => rx_input_memio_bpl(5)
    );
  rx_input_memio_bpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_5_FFX_RST
    );
  rx_input_memio_bpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(6),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_7_FFY_RST,
      O => rx_input_memio_bpl(6)
    );
  rx_input_memio_bpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_7_FFY_RST
    );
  rx_input_memio_bpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(7),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_7_FFX_RST,
      O => rx_input_memio_bpl(7)
    );
  rx_input_memio_bpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_7_FFX_RST
    );
  rx_input_memio_bpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(8),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_9_FFY_RST,
      O => rx_input_memio_bpl(8)
    );
  rx_input_memio_bpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_9_FFY_RST
    );
  rx_input_memio_bpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(9),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_9_FFX_RST,
      O => rx_input_memio_bpl(9)
    );
  rx_input_memio_bpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_9_FFX_RST
    );
  mac_control_PHY_status_din_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(10),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_11_FFY_RST,
      O => mac_control_PHY_status_din(10)
    );
  mac_control_PHY_status_din_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_11_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd6_1971 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd6_In,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => mac_control_PHY_status_MII_Interface_cs_FFd6_FFY_SET,
      RST => GND,
      O => mac_control_PHY_status_MII_Interface_cs_FFd6
    );
  mac_control_PHY_status_MII_Interface_cs_FFd6_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => mac_control_PHY_status_MII_Interface_cs_FFd6_FFY_SET
    );
  rx_fifocheck_fbbpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_3_FFY_RST,
      O => rx_fifocheck_fbbpl(2)
    );
  rx_fifocheck_fbbpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_3_FFY_RST
    );
  rx_fifocheck_fbbpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_3_FFX_RST,
      O => rx_fifocheck_fbbpl(3)
    );
  rx_fifocheck_fbbpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_3_FFX_RST
    );
  rx_fifocheck_fbbpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_5_FFY_RST,
      O => rx_fifocheck_fbbpl(4)
    );
  rx_fifocheck_fbbpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_5_FFY_RST
    );
  rx_fifocheck_fbbpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_5_FFX_RST,
      O => rx_fifocheck_fbbpl(5)
    );
  rx_fifocheck_fbbpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_5_FFX_RST
    );
  rx_fifocheck_fbbpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_7_FFY_RST,
      O => rx_fifocheck_fbbpl(6)
    );
  rx_fifocheck_fbbpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_7_FFY_RST
    );
  rx_fifocheck_fbbpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_7_FFX_RST,
      O => rx_fifocheck_fbbpl(7)
    );
  rx_fifocheck_fbbpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_7_FFX_RST
    );
  rx_fifocheck_fbbpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_9_FFY_RST,
      O => rx_fifocheck_fbbpl(8)
    );
  rx_fifocheck_fbbpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_9_FFY_RST
    );
  rx_input_memio_cs_FFd5_1972 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd6,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd6_FFY_RST,
      O => rx_input_memio_cs_FFd5
    );
  rx_input_memio_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd6_FFY_RST
    );
  rx_fifocheck_fbbpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_9_FFX_RST,
      O => rx_fifocheck_fbbpl(9)
    );
  rx_fifocheck_fbbpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_9_FFX_RST
    );
  rx_input_memio_cs_FFd1_1973 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd2,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd2_FFY_RST,
      O => rx_input_memio_cs_FFd1
    );
  rx_input_memio_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd2_FFY_RST
    );
  tx_output_crcl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(23),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_23_FFY_RST,
      O => tx_output_crcl(23)
    );
  tx_output_crcl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_23_FFY_RST
    );
  rx_input_memio_cs_FFd2_1974 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd4,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd2_FFX_RST,
      O => rx_input_memio_cs_FFd2
    );
  rx_input_memio_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd2_FFX_RST
    );
  rx_input_memio_cs_FFd6_1975 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd7,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd6_FFX_RST,
      O => rx_input_memio_cs_FFd6
    );
  rx_input_memio_cs_FFd6_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd6_FFX_RST
    );
  tx_output_crcl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(15),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_15_FFY_RST,
      O => tx_output_crcl(15)
    );
  tx_output_crcl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_15_FFY_RST
    );
  mac_control_dout_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N77167,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_5_FFY_RST,
      O => mac_control_dout(5)
    );
  mac_control_dout_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_5_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(1),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_1_FFX_RST,
      O => mac_control_phydo(1)
    );
  mac_control_phydo_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_1_FFX_RST
    );
  rx_input_memio_crcl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(10),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_10_FFY_RST,
      O => rx_input_memio_crcl(10)
    );
  rx_input_memio_crcl_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_10_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(0),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_1_FFY_RST,
      O => mac_control_phydo(0)
    );
  mac_control_phydo_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_1_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(3),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_3_FFX_RST,
      O => mac_control_phydo(3)
    );
  mac_control_phydo_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_3_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(6),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_7_FFY_RST,
      O => mac_control_phydo(6)
    );
  mac_control_phydo_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_7_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(4),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_5_FFY_RST,
      O => mac_control_phydo(4)
    );
  mac_control_phydo_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_5_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(5),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_5_FFX_RST,
      O => mac_control_phydo(5)
    );
  mac_control_phydo_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_5_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(7),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_7_FFX_RST,
      O => mac_control_phydo(7)
    );
  mac_control_phydo_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_7_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(8),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_9_FFY_RST,
      O => mac_control_phydo(8)
    );
  mac_control_phydo_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_9_FFY_RST
    );
  rx_input_memio_crcl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(8),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_8_FFY_RST,
      O => rx_input_memio_crcl(8)
    );
  rx_input_memio_crcl_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_8_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(9),
      CE => mac_control_PHY_status_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_9_FFX_RST,
      O => mac_control_phydo(9)
    );
  mac_control_phydo_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_9_FFX_RST
    );
  memcontroller_dnl2_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(29),
      CE => memcontroller_dnl2_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_29_FFX_RST,
      O => memcontroller_dnl2(29)
    );
  memcontroller_dnl2_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_29_FFX_RST
    );
  rx_input_memio_datal_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_datal_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_1_FFX_RST,
      O => rx_input_memio_datal(1)
    );
  rx_input_memio_datal_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_1_FFX_RST
    );
  rx_input_memio_datal_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_datal_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_3_FFY_RST,
      O => rx_input_memio_datal(2)
    );
  rx_input_memio_datal_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_3_FFY_RST
    );
  rx_input_memio_datal_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_datal_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_3_FFX_RST,
      O => rx_input_memio_datal(3)
    );
  rx_input_memio_datal_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_3_FFX_RST
    );
  rx_input_memio_datal_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_datal_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_5_FFY_RST,
      O => rx_input_memio_datal(4)
    );
  rx_input_memio_datal_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_5_FFY_RST
    );
  rx_input_memio_datal_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_datal_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_5_FFX_RST,
      O => rx_input_memio_datal(5)
    );
  rx_input_memio_datal_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_5_FFX_RST
    );
  rx_input_memio_datal_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_datal_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_7_FFY_RST,
      O => rx_input_memio_datal(6)
    );
  rx_input_memio_datal_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_7_FFY_RST
    );
  rx_input_memio_datal_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_datal_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_7_FFX_RST,
      O => rx_input_memio_datal(7)
    );
  rx_input_memio_datal_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_7_FFX_RST
    );
  rx_input_memio_addrchk_maceq_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq(1),
      CE => rx_input_memio_addrchk_maceq_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_0_FFY_RST,
      O => rx_input_memio_addrchk_maceq(1)
    );
  rx_input_memio_addrchk_maceq_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_0_FFY_RST
    );
  rx_input_memio_addrchk_maceq_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq_0_rt,
      CE => rx_input_memio_addrchk_maceq_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_0_FFX_RST,
      O => rx_input_memio_addrchk_maceq(0)
    );
  rx_input_memio_addrchk_maceq_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_0_FFX_RST
    );
  rx_input_memio_addrchk_maceq_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq(3),
      CE => rx_input_memio_addrchk_maceq_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_2_FFY_RST,
      O => rx_input_memio_addrchk_maceq(3)
    );
  rx_input_memio_addrchk_maceq_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_2_FFY_RST
    );
  rx_input_memio_addrchk_maceq_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq(5),
      CE => rx_input_memio_addrchk_maceq_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_4_FFY_RST,
      O => rx_input_memio_addrchk_maceq(5)
    );
  rx_input_memio_addrchk_maceq_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_4_FFY_RST
    );
  rx_input_memio_addrchk_datal_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_13_FFX_RST,
      O => rx_input_memio_addrchk_datal(13)
    );
  rx_input_memio_addrchk_datal_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_13_FFX_RST
    );
  rx_input_memio_addrchk_datal_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_23_FFY_RST,
      O => rx_input_memio_addrchk_datal(22)
    );
  rx_input_memio_addrchk_datal_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_23_FFY_RST
    );
  rx_input_memio_addrchk_datal_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_31_FFX_RST,
      O => rx_input_memio_addrchk_datal(31)
    );
  rx_input_memio_addrchk_datal_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_31_FFX_RST
    );
  rx_input_memio_addrchk_datal_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_23_FFX_RST,
      O => rx_input_memio_addrchk_datal(23)
    );
  rx_input_memio_addrchk_datal_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_23_FFX_RST
    );
  rx_input_memio_addrchk_datal_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_15_FFY_RST,
      O => rx_input_memio_addrchk_datal(14)
    );
  rx_input_memio_addrchk_datal_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_15_FFY_RST
    );
  rx_input_memio_addrchk_datal_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_15_FFX_RST,
      O => rx_input_memio_addrchk_datal(15)
    );
  rx_input_memio_addrchk_datal_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_15_FFX_RST
    );
  rx_input_memio_addrchk_datal_40 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_41_FFY_RST,
      O => rx_input_memio_addrchk_datal(40)
    );
  rx_input_memio_addrchk_datal_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_41_FFY_RST
    );
  rx_input_memio_addrchk_datal_32 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_33_FFY_RST,
      O => rx_input_memio_addrchk_datal(32)
    );
  rx_input_memio_addrchk_datal_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_33_FFY_RST
    );
  rx_input_memio_addrchk_datal_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_25_FFY_RST,
      O => rx_input_memio_addrchk_datal(24)
    );
  rx_input_memio_addrchk_datal_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_25_FFY_RST
    );
  rx_input_memio_addrchk_datal_33 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_33_FFX_RST,
      O => rx_input_memio_addrchk_datal(33)
    );
  rx_input_memio_addrchk_datal_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_33_FFX_RST
    );
  rx_input_memio_addrchk_datal_41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_41_FFX_RST,
      O => rx_input_memio_addrchk_datal(41)
    );
  rx_input_memio_addrchk_datal_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_41_FFX_RST
    );
  rx_input_memio_addrchk_datal_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_25_FFX_RST,
      O => rx_input_memio_addrchk_datal(25)
    );
  rx_input_memio_addrchk_datal_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_25_FFX_RST
    );
  rx_input_memio_addrchk_datal_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_17_FFY_RST,
      O => rx_input_memio_addrchk_datal(16)
    );
  rx_input_memio_addrchk_datal_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_17_FFY_RST
    );
  rx_input_memio_addrchk_datal_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_17_FFX_RST,
      O => rx_input_memio_addrchk_datal(17)
    );
  rx_input_memio_addrchk_datal_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_17_FFX_RST
    );
  rx_input_memio_addrchk_datal_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_27_FFY_RST,
      O => rx_input_memio_addrchk_datal(26)
    );
  rx_input_memio_addrchk_datal_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_27_FFY_RST
    );
  rx_input_memio_addrchk_datal_34 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_35_FFY_RST,
      O => rx_input_memio_addrchk_datal(34)
    );
  rx_input_memio_addrchk_datal_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_35_FFY_RST
    );
  rx_input_memio_addrchk_datal_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_27_FFX_RST,
      O => rx_input_memio_addrchk_datal(27)
    );
  rx_input_memio_addrchk_datal_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_27_FFX_RST
    );
  rx_input_memio_crcll_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(9),
      CE => rx_input_memio_crcll_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_9_FFX_RST,
      O => rx_input_memio_crcll(9)
    );
  rx_input_memio_crcll_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_9_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(6),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_7_FFY_RST,
      O => mac_control_phystat(6)
    );
  mac_control_phystat_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_7_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(8),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_9_FFY_RST,
      O => mac_control_phystat(8)
    );
  mac_control_phystat_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_9_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(7),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_7_FFX_RST,
      O => mac_control_phystat(7)
    );
  mac_control_phystat_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_7_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(9),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_9_FFX_RST,
      O => mac_control_phystat(9)
    );
  mac_control_phystat_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_9_FFX_RST
    );
  tx_output_crcl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(17),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_17_FFY_RST,
      O => tx_output_crcl(17)
    );
  tx_output_crcl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_17_FFY_RST
    );
  rx_input_memio_crcl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(12),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_12_FFY_RST,
      O => rx_input_memio_crcl(12)
    );
  rx_input_memio_crcl_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_12_FFY_RST
    );
  rx_fifocheck_fbbpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_11_FFY_RST,
      O => rx_fifocheck_fbbpl(10)
    );
  rx_fifocheck_fbbpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_11_FFY_RST
    );
  rx_fifocheck_fbbpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_11_FFX_RST,
      O => rx_fifocheck_fbbpl(11)
    );
  rx_fifocheck_fbbpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_11_FFX_RST
    );
  rx_fifocheck_fbbpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_13_FFY_RST,
      O => rx_fifocheck_fbbpl(12)
    );
  rx_fifocheck_fbbpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_13_FFY_RST
    );
  rx_fifocheck_fbbpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_13_FFX_RST,
      O => rx_fifocheck_fbbpl(13)
    );
  rx_fifocheck_fbbpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_13_FFX_RST
    );
  rx_fifocheck_fbbpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_15_FFY_RST,
      O => rx_fifocheck_fbbpl(14)
    );
  rx_fifocheck_fbbpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_15_FFY_RST
    );
  mac_control_dout_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N79702,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_7_FFY_RST,
      O => mac_control_dout(7)
    );
  mac_control_dout_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_7_FFY_RST
    );
  mac_control_dout_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N78742,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_9_FFY_RST,
      O => mac_control_dout(9)
    );
  mac_control_dout_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_9_FFY_RST
    );
  tx_output_crcl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(27),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_27_FFY_RST,
      O => tx_output_crcl(27)
    );
  tx_output_crcl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_27_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(23),
      CE => rx_input_memio_addrchk_macaddrl_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_23_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(23)
    );
  rx_input_memio_addrchk_macaddrl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_23_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(15),
      CE => rx_input_memio_addrchk_macaddrl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_15_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(15)
    );
  rx_input_memio_addrchk_macaddrl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_15_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(41),
      CE => rx_input_memio_addrchk_macaddrl_41_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_41_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(41)
    );
  rx_input_memio_addrchk_macaddrl_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_41_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_33 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(33),
      CE => rx_input_memio_addrchk_macaddrl_33_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_33_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(33)
    );
  rx_input_memio_addrchk_macaddrl_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_33_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(25),
      CE => rx_input_memio_addrchk_macaddrl_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_25_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(25)
    );
  rx_input_memio_addrchk_macaddrl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_25_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(17),
      CE => rx_input_memio_addrchk_macaddrl_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_17_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(17)
    );
  rx_input_memio_addrchk_macaddrl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_17_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_43 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(43),
      CE => rx_input_memio_addrchk_macaddrl_43_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_43_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(43)
    );
  rx_input_memio_addrchk_macaddrl_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_43_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_34 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(34),
      CE => rx_input_memio_addrchk_macaddrl_35_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_35_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(34)
    );
  rx_input_memio_addrchk_macaddrl_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_35_FFY_RST
    );
  rx_input_memio_addrchk_datal_35 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_35_FFX_RST,
      O => rx_input_memio_addrchk_datal(35)
    );
  rx_input_memio_addrchk_datal_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_35_FFX_RST
    );
  rx_input_memio_addrchk_datal_42 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_43_FFY_RST,
      O => rx_input_memio_addrchk_datal(42)
    );
  rx_input_memio_addrchk_datal_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_43_FFY_RST
    );
  rx_input_memio_addrchk_datal_43 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_43_FFX_RST,
      O => rx_input_memio_addrchk_datal(43)
    );
  rx_input_memio_addrchk_datal_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_43_FFX_RST
    );
  rx_input_memio_addrchk_datal_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_19_FFY_RST,
      O => rx_input_memio_addrchk_datal(18)
    );
  rx_input_memio_addrchk_datal_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_19_FFY_RST
    );
  rx_input_memio_addrchk_datal_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_19_FFX_RST,
      O => rx_input_memio_addrchk_datal(19)
    );
  rx_input_memio_addrchk_datal_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_19_FFX_RST
    );
  rx_input_memio_addrchk_datal_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_29_FFY_RST,
      O => rx_input_memio_addrchk_datal(28)
    );
  rx_input_memio_addrchk_datal_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_29_FFY_RST
    );
  rx_input_memio_addrchk_datal_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_29_FFX_RST,
      O => rx_input_memio_addrchk_datal(29)
    );
  rx_input_memio_addrchk_datal_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_29_FFX_RST
    );
  rx_input_memio_addrchk_datal_36 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_37_FFY_RST,
      O => rx_input_memio_addrchk_datal(36)
    );
  rx_input_memio_addrchk_datal_37_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_37_FFY_RST
    );
  rx_input_memio_addrchk_datal_37 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_37_FFX_RST,
      O => rx_input_memio_addrchk_datal(37)
    );
  rx_input_memio_addrchk_datal_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_37_FFX_RST
    );
  rx_input_memio_addrchk_datal_44 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_45_FFY_RST,
      O => rx_input_memio_addrchk_datal(44)
    );
  rx_input_memio_addrchk_datal_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_45_FFY_RST
    );
  rx_input_memio_addrchk_datal_45 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_45_FFX_RST,
      O => rx_input_memio_addrchk_datal(45)
    );
  rx_input_memio_addrchk_datal_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_45_FFX_RST
    );
  rx_input_memio_addrchk_datal_38 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_39_FFY_RST,
      O => rx_input_memio_addrchk_datal(38)
    );
  rx_input_memio_addrchk_datal_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_39_FFY_RST
    );
  rx_input_memio_addrchk_datal_39 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_39_FFX_RST,
      O => rx_input_memio_addrchk_datal(39)
    );
  rx_input_memio_addrchk_datal_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_39_FFX_RST
    );
  rx_input_memio_addrchk_datal_46 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_47_FFY_RST,
      O => rx_input_memio_addrchk_datal(46)
    );
  rx_input_memio_addrchk_datal_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_47_FFY_RST
    );
  rx_input_memio_crcll_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(0),
      CE => rx_input_memio_crcll_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_1_FFY_RST,
      O => rx_input_memio_crcll(0)
    );
  rx_input_memio_crcll_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_1_FFY_RST
    );
  rx_input_memio_addrchk_datal_47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_47_FFX_RST,
      O => rx_input_memio_addrchk_datal(47)
    );
  rx_input_memio_addrchk_datal_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_47_FFX_RST
    );
  rx_input_memio_doutl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(1),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_1_FFX_RST,
      O => rx_input_memio_doutl(1)
    );
  rx_input_memio_doutl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_1_FFX_RST
    );
  rx_input_memio_doutl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(0),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_1_FFY_RST,
      O => rx_input_memio_doutl(0)
    );
  rx_input_memio_doutl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_1_FFY_RST
    );
  rx_input_memio_doutl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(2),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_3_FFY_RST,
      O => rx_input_memio_doutl(2)
    );
  rx_input_memio_doutl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_3_FFY_RST
    );
  rx_input_memio_doutl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(3),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_3_FFX_RST,
      O => rx_input_memio_doutl(3)
    );
  rx_input_memio_doutl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_3_FFX_RST
    );
  rx_input_memio_doutl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(4),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_5_FFY_RST,
      O => rx_input_memio_doutl(4)
    );
  rx_input_memio_doutl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_5_FFY_RST
    );
  rx_input_memio_doutl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(5),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_5_FFX_RST,
      O => rx_input_memio_doutl(5)
    );
  rx_input_memio_doutl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_5_FFX_RST
    );
  rx_input_memio_doutl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(6),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_7_FFY_RST,
      O => rx_input_memio_doutl(6)
    );
  rx_input_memio_doutl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_7_FFY_RST
    );
  mac_control_lrxallf_1976 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0238,
      CLK => GTX_CLK_OBUF,
      SET => mac_control_lrxallf_FFY_SET,
      RST => GND,
      O => mac_control_lrxallf
    );
  mac_control_lrxallf_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => mac_control_lrxallf_FFY_SET
    );
  rx_input_memio_doutl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(7),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_7_FFX_RST,
      O => rx_input_memio_doutl(7)
    );
  rx_input_memio_doutl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_7_FFX_RST
    );
  rx_input_memio_doutl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(8),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_9_FFY_RST,
      O => rx_input_memio_doutl(8)
    );
  rx_input_memio_doutl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_9_FFY_RST
    );
  rx_input_memio_doutl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(9),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_9_FFX_RST,
      O => rx_input_memio_doutl(9)
    );
  rx_input_memio_doutl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_9_FFX_RST
    );
  mac_control_dout_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N77375,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_8_FFY_RST,
      O => mac_control_dout(8)
    );
  mac_control_dout_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_8_FFY_RST
    );
  rx_input_memio_wbpl_1977 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd2,
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_wbpl_FFY_RST,
      O => rx_input_memio_wbpl
    );
  rx_input_memio_wbpl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_wbpl_FFY_RST
    );
  rx_input_memio_crcl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(19),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_19_FFY_RST,
      O => rx_input_memio_crcl(19)
    );
  rx_input_memio_crcl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_19_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(13),
      CE => mac_control_PHY_status_MII_Interface_N72822,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_14_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(14)
    );
  mac_control_PHY_status_MII_Interface_dreg_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_14_FFX_RST
    );
  rx_input_memio_dout_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_25_FFY_RST,
      O => rx_input_memio_dout(24)
    );
  rx_input_memio_dout_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_25_FFY_RST
    );
  rx_input_memio_dout_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_25_FFX_RST,
      O => rx_input_memio_dout(25)
    );
  rx_input_memio_dout_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_25_FFX_RST
    );
  rx_input_memio_dout_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_17_FFX_RST,
      O => rx_input_memio_dout(17)
    );
  rx_input_memio_dout_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_17_FFX_RST
    );
  rx_input_memio_dout_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_27_FFY_RST,
      O => rx_input_memio_dout(26)
    );
  rx_input_memio_dout_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_27_FFY_RST
    );
  rx_input_memio_dout_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_27_FFX_RST,
      O => rx_input_memio_dout(27)
    );
  rx_input_memio_dout_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_27_FFX_RST
    );
  rx_input_memio_dout_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_19_FFX_RST,
      O => rx_input_memio_dout(19)
    );
  rx_input_memio_dout_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_19_FFX_RST
    );
  rx_input_memio_dout_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_29_FFX_RST,
      O => rx_input_memio_dout(29)
    );
  rx_input_memio_dout_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_29_FFX_RST
    );
  mac_control_phydi_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_3_FFY_RST,
      O => mac_control_phydi(2)
    );
  mac_control_phydi_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_3_FFY_RST
    );
  mac_control_phydi_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_1_FFX_RST,
      O => mac_control_phydi(1)
    );
  mac_control_phydi_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_1_FFX_RST
    );
  mac_control_phydi_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_5_FFY_RST,
      O => mac_control_phydi(4)
    );
  mac_control_phydi_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_5_FFY_RST
    );
  mac_control_phydi_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_3_FFX_RST,
      O => mac_control_phydi(3)
    );
  mac_control_phydi_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_3_FFX_RST
    );
  mac_control_phydi_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_5_FFX_RST,
      O => mac_control_phydi(5)
    );
  mac_control_phydi_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_5_FFX_RST
    );
  mac_control_phydi_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_7_FFY_RST,
      O => mac_control_phydi(6)
    );
  mac_control_phydi_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_7_FFY_RST
    );
  mac_control_phydi_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_7_FFX_RST,
      O => mac_control_phydi(7)
    );
  mac_control_phydi_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_7_FFX_RST
    );
  mac_control_phydi_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_9_FFY_RST,
      O => mac_control_phydi(8)
    );
  mac_control_phydi_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_9_FFY_RST
    );
  mac_control_phydi_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_9_FFX_RST,
      O => mac_control_phydi(9)
    );
  mac_control_phydi_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_9_FFX_RST
    );
  rx_input_memio_bpen_1978 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd2,
      CE => rx_input_memio_bpen_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpen_FFY_RST,
      O => rx_input_memio_bpen
    );
  rx_input_memio_bpen_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpen_FFY_RST
    );
  rx_input_memio_addrchk_DESTOK : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_n0053,
      CE => rx_input_memio_destok_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_destok_FFY_RST,
      O => rx_input_memio_destok
    );
  rx_input_memio_destok_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_destok_FFY_RST
    );
  rx_output_cs_FFd10_1979 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd10_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd10_FFY_RST,
      O => rx_output_cs_FFd10
    );
  rx_output_cs_FFd10_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd10_FFY_RST
    );
  tx_output_crcl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(18),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_18_FFY_RST,
      O => tx_output_crcl(18)
    );
  tx_output_crcl_18_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_18_FFY_RST
    );
  tx_output_crcl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(26),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_26_FFY_RST,
      O => tx_output_crcl(26)
    );
  tx_output_crcl_26_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_26_FFY_RST
    );
  mac_control_dout_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N79540,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_3_FFY_RST,
      O => mac_control_dout(3)
    );
  mac_control_dout_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_3_FFY_RST
    );
  mac_control_dout_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_N78585,
      CE => mac_control_N70898,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_dout_4_FFY_RST,
      O => mac_control_dout(4)
    );
  mac_control_dout_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_4_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_35 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(35),
      CE => rx_input_memio_addrchk_macaddrl_35_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_35_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(35)
    );
  rx_input_memio_addrchk_macaddrl_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_35_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(27),
      CE => rx_input_memio_addrchk_macaddrl_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_27_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(27)
    );
  rx_input_memio_addrchk_macaddrl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_27_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(19),
      CE => rx_input_memio_addrchk_macaddrl_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_19_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(19)
    );
  rx_input_memio_addrchk_macaddrl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_19_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_45 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(45),
      CE => rx_input_memio_addrchk_macaddrl_45_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_45_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(45)
    );
  rx_input_memio_addrchk_macaddrl_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_45_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_37 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(37),
      CE => rx_input_memio_addrchk_macaddrl_37_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_37_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(37)
    );
  rx_input_memio_addrchk_macaddrl_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_37_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(29),
      CE => rx_input_memio_addrchk_macaddrl_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_29_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(29)
    );
  rx_input_memio_addrchk_macaddrl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_29_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_38 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(38),
      CE => rx_input_memio_addrchk_macaddrl_39_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_39_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(38)
    );
  rx_input_memio_addrchk_macaddrl_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_39_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(47),
      CE => rx_input_memio_addrchk_macaddrl_47_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_47_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(47)
    );
  rx_input_memio_addrchk_macaddrl_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_47_FFX_RST
    );
  slowclock_rxphyerrl_1980 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_rxphyerrl_GROM,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => rxphyerr,
      SRST => slowclock_rxphyerrl_LOGIC_ZERO,
      O => slowclock_rxphyerrl
    );
  rx_input_memio_crcl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(13),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_13_FFY_RST,
      O => rx_input_memio_crcl(13)
    );
  rx_input_memio_crcl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_13_FFY_RST
    );
  tx_input_cs_FFd12_1981 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => tx_input_cs_FFd12_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => tx_input_cs_FFd12_FFY_SET,
      RST => GND,
      O => tx_input_cs_FFd12
    );
  tx_input_cs_FFd12_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF_1,
      O => tx_input_cs_FFd12_FFY_SET
    );
  rx_input_memio_addrchk_macaddrl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(10),
      CE => rx_input_memio_addrchk_macaddrl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_11_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(10)
    );
  rx_input_memio_addrchk_macaddrl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_11_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(11),
      CE => rx_input_memio_addrchk_macaddrl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_11_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(11)
    );
  rx_input_memio_addrchk_macaddrl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_11_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(21),
      CE => rx_input_memio_addrchk_macaddrl_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_21_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(21)
    );
  rx_input_memio_addrchk_macaddrl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_21_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(13),
      CE => rx_input_memio_addrchk_macaddrl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_13_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(13)
    );
  rx_input_memio_addrchk_macaddrl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_13_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(31),
      CE => rx_input_memio_addrchk_macaddrl_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_31_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(31)
    );
  rx_input_memio_addrchk_macaddrl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_31_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(22),
      CE => rx_input_memio_addrchk_macaddrl_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_23_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(22)
    );
  rx_input_memio_addrchk_macaddrl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_23_FFY_RST
    );
  rx_input_memio_crcll_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(15),
      CE => rx_input_memio_crcll_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_15_FFX_RST,
      O => rx_input_memio_crcll(15)
    );
  rx_input_memio_crcll_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_15_FFX_RST
    );
  rx_input_memio_crcll_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(30),
      CE => rx_input_memio_crcll_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_31_FFY_RST,
      O => rx_input_memio_crcll(30)
    );
  rx_input_memio_crcll_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_31_FFY_RST
    );
  rx_input_memio_crcll_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(31),
      CE => rx_input_memio_crcll_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_31_FFX_RST,
      O => rx_input_memio_crcll(31)
    );
  rx_input_memio_crcll_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_31_FFX_RST
    );
  rx_input_memio_crcll_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(22),
      CE => rx_input_memio_crcll_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_23_FFY_RST,
      O => rx_input_memio_crcll(22)
    );
  rx_input_memio_crcll_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_23_FFY_RST
    );
  rx_input_memio_crcll_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(23),
      CE => rx_input_memio_crcll_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_23_FFX_RST,
      O => rx_input_memio_crcll(23)
    );
  rx_input_memio_crcll_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_23_FFX_RST
    );
  rx_input_memio_crcll_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(16),
      CE => rx_input_memio_crcll_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_17_FFY_RST,
      O => rx_input_memio_crcll(16)
    );
  rx_input_memio_crcll_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_17_FFY_RST
    );
  rx_input_memio_crcll_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(24),
      CE => rx_input_memio_crcll_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_25_FFY_RST,
      O => rx_input_memio_crcll(24)
    );
  rx_input_memio_crcll_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_25_FFY_RST
    );
  rx_input_memio_crcll_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(17),
      CE => rx_input_memio_crcll_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_17_FFX_RST,
      O => rx_input_memio_crcll(17)
    );
  rx_input_memio_crcll_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_17_FFX_RST
    );
  rx_input_memio_crcll_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(25),
      CE => rx_input_memio_crcll_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_25_FFX_RST,
      O => rx_input_memio_crcll(25)
    );
  rx_input_memio_crcll_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_25_FFX_RST
    );
  rx_input_memio_crcll_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(26),
      CE => rx_input_memio_crcll_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_27_FFY_RST,
      O => rx_input_memio_crcll(26)
    );
  rx_input_memio_crcll_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_27_FFY_RST
    );
  rx_input_memio_crcll_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(27),
      CE => rx_input_memio_crcll_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_27_FFX_RST,
      O => rx_input_memio_crcll(27)
    );
  rx_input_memio_crcll_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_27_FFX_RST
    );
  rx_input_memio_crcll_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(18),
      CE => rx_input_memio_crcll_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_19_FFY_RST,
      O => rx_input_memio_crcll(18)
    );
  rx_input_memio_crcll_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_19_FFY_RST
    );
  rx_input_memio_crcll_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(19),
      CE => rx_input_memio_crcll_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_19_FFX_RST,
      O => rx_input_memio_crcll(19)
    );
  rx_input_memio_crcll_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_19_FFX_RST
    );
  rx_input_memio_crcll_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(28),
      CE => rx_input_memio_crcll_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_29_FFY_RST,
      O => rx_input_memio_crcll(28)
    );
  rx_input_memio_crcll_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_29_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_39 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(39),
      CE => rx_input_memio_addrchk_macaddrl_39_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_39_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(39)
    );
  rx_input_memio_addrchk_macaddrl_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_39_FFX_RST
    );
  tx_output_crcl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(28),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_28_FFY_RST,
      O => tx_output_crcl(28)
    );
  tx_output_crcl_28_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_28_FFY_RST
    );
  rx_input_memio_crcl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(23),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_23_FFY_RST,
      O => rx_input_memio_crcl(23)
    );
  rx_input_memio_crcl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_23_FFY_RST
    );
  rx_input_memio_crcl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(15),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_15_FFY_RST,
      O => rx_input_memio_crcl(15)
    );
  rx_input_memio_crcl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_15_FFY_RST
    );
  rx_input_memio_crcll_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(29),
      CE => rx_input_memio_crcll_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_29_FFX_RST,
      O => rx_input_memio_crcll(29)
    );
  rx_input_memio_crcll_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_29_FFX_RST
    );
  rx_input_memio_crcl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(24),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_24_FFY_RST,
      O => rx_input_memio_crcl(24)
    );
  rx_input_memio_crcl_24_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_24_FFY_RST
    );
  rx_input_memio_crcl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(16),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_16_FFY_RST,
      O => rx_input_memio_crcl(16)
    );
  rx_input_memio_crcl_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_16_FFY_RST
    );
  rx_input_memio_addrchk_rxallfl_1982 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxallf,
      CE => rx_input_memio_addrchk_rxallfl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_rxallfl_FFY_RST,
      O => rx_input_memio_addrchk_rxallfl
    );
  rx_input_memio_addrchk_rxallfl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_rxallfl_FFY_RST
    );
  tx_fifocheck_bpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_1_FFY_RST,
      O => tx_fifocheck_bpl(0)
    );
  tx_fifocheck_bpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_1_FFY_RST
    );
  tx_fifocheck_bpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_1_FFX_RST,
      O => tx_fifocheck_bpl(1)
    );
  tx_fifocheck_bpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_1_FFX_RST
    );
  tx_fifocheck_bpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_3_FFY_RST,
      O => tx_fifocheck_bpl(2)
    );
  tx_fifocheck_bpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_3_FFY_RST
    );
  tx_fifocheck_bpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_3_FFX_RST,
      O => tx_fifocheck_bpl(3)
    );
  tx_fifocheck_bpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_3_FFX_RST
    );
  tx_fifocheck_bpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_5_FFY_RST,
      O => tx_fifocheck_bpl(4)
    );
  tx_fifocheck_bpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_5_FFY_RST
    );
  tx_fifocheck_bpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_7_FFY_RST,
      O => tx_fifocheck_bpl(6)
    );
  tx_fifocheck_bpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_7_FFY_RST
    );
  tx_fifocheck_bpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_5_FFX_RST,
      O => tx_fifocheck_bpl(5)
    );
  tx_fifocheck_bpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_5_FFX_RST
    );
  tx_fifocheck_bpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_7_FFX_RST,
      O => tx_fifocheck_bpl(7)
    );
  tx_fifocheck_bpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_7_FFX_RST
    );
  tx_fifocheck_bpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_9_FFY_RST,
      O => tx_fifocheck_bpl(8)
    );
  tx_fifocheck_bpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_9_FFY_RST
    );
  tx_fifocheck_bpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_9_FFX_RST,
      O => tx_fifocheck_bpl(9)
    );
  tx_fifocheck_bpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_9_FFX_RST
    );
  tx_output_crcl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(29),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_29_FFY_RST,
      O => tx_output_crcl(29)
    );
  tx_output_crcl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_29_FFY_RST
    );
  rx_input_memio_crcll_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(11),
      CE => rx_input_memio_crcll_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_11_FFX_RST,
      O => rx_input_memio_crcll(11)
    );
  rx_input_memio_crcll_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_11_FFX_RST
    );
  rx_input_memio_crcll_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(10),
      CE => rx_input_memio_crcll_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_11_FFY_RST,
      O => rx_input_memio_crcll(10)
    );
  rx_input_memio_crcll_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_11_FFY_RST
    );
  rx_input_memio_crcll_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(12),
      CE => rx_input_memio_crcll_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_13_FFY_RST,
      O => rx_input_memio_crcll(12)
    );
  rx_input_memio_crcll_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_13_FFY_RST
    );
  rx_input_memio_crcll_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(13),
      CE => rx_input_memio_crcll_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_13_FFX_RST,
      O => rx_input_memio_crcll(13)
    );
  rx_input_memio_crcll_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_13_FFX_RST
    );
  rx_input_memio_crcll_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(20),
      CE => rx_input_memio_crcll_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_21_FFY_RST,
      O => rx_input_memio_crcll(20)
    );
  rx_input_memio_crcll_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_21_FFY_RST
    );
  rx_input_memio_crcll_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(21),
      CE => rx_input_memio_crcll_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_21_FFX_RST,
      O => rx_input_memio_crcll(21)
    );
  rx_input_memio_crcll_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_21_FFX_RST
    );
  rx_input_memio_crcll_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(14),
      CE => rx_input_memio_crcll_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_15_FFY_RST,
      O => rx_input_memio_crcll(14)
    );
  rx_input_memio_crcll_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_15_FFY_RST
    );
  rx_input_memio_doutl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(19),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_19_FFX_RST,
      O => rx_input_memio_doutl(19)
    );
  rx_input_memio_doutl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_19_FFX_RST
    );
  rx_input_memio_doutl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(28),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_29_FFY_RST,
      O => rx_input_memio_doutl(28)
    );
  rx_input_memio_doutl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_29_FFY_RST
    );
  rx_input_memio_doutl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(29),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_29_FFX_RST,
      O => rx_input_memio_doutl(29)
    );
  rx_input_memio_doutl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_29_FFX_RST
    );
  rx_input_fifo_control_d0_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(0),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_1_FFY_RST,
      O => rx_input_fifo_control_d0(0)
    );
  rx_input_fifo_control_d0_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_1_FFY_RST
    );
  rx_input_fifo_control_d0_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(1),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_1_FFX_RST,
      O => rx_input_fifo_control_d0(1)
    );
  rx_input_fifo_control_d0_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_1_FFX_RST
    );
  rx_input_fifo_control_d0_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(3),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_3_FFX_RST,
      O => rx_input_fifo_control_d0(3)
    );
  rx_input_fifo_control_d0_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_3_FFX_RST
    );
  rx_input_fifo_control_d0_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(5),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_5_FFX_RST,
      O => rx_input_fifo_control_d0(5)
    );
  rx_input_fifo_control_d0_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_5_FFX_RST
    );
  rx_input_fifo_control_d1_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(1),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_1_FFX_RST,
      O => rx_input_fifo_control_d1(1)
    );
  rx_input_fifo_control_d1_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_1_FFX_RST
    );
  rx_input_fifo_control_d0_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(6),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_7_FFY_RST,
      O => rx_input_fifo_control_d0(6)
    );
  rx_input_fifo_control_d0_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_7_FFY_RST
    );
  rx_input_fifo_control_d0_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(7),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_7_FFX_RST,
      O => rx_input_fifo_control_d0(7)
    );
  rx_input_fifo_control_d0_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_7_FFX_RST
    );
  rx_input_fifo_control_d1_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(3),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_3_FFX_RST,
      O => rx_input_fifo_control_d1(3)
    );
  rx_input_fifo_control_d1_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_3_FFX_RST
    );
  rx_input_fifo_control_d1_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(4),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_5_FFY_RST,
      O => rx_input_fifo_control_d1(4)
    );
  rx_input_fifo_control_d1_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_5_FFY_RST
    );
  rx_input_fifo_control_d0_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(8),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_8_FFY_RST,
      O => rx_input_fifo_control_d0(8)
    );
  rx_input_fifo_control_d0_8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_8_FFY_RST
    );
  slowclock_RXFSR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_rxfl,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfsr_FFY_RST,
      O => rxfsr
    );
  rxfsr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfsr_FFY_RST
    );
  slowclock_TXFSR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_txfl,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfsr_FFY_RST,
      O => txfsr
    );
  txfsr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfsr_FFY_RST
    );
  rx_input_memio_crcl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(29),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_29_FFY_RST,
      O => rx_input_memio_crcl(29)
    );
  rx_input_memio_crcl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_29_FFY_RST
    );
  rx_input_fifo_control_celll_1983 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_cell,
      CE => rx_input_fifo_control_celll_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_celll_FFY_RST,
      O => rx_input_fifo_control_celll
    );
  rx_input_fifo_control_celll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_celll_FFY_RST
    );
  mac_control_ledrx_rst_1984 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cross,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledrx_rst_FFY_RST,
      O => mac_control_ledrx_rst
    );
  mac_control_ledrx_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_rst_FFY_RST
    );
  mac_control_MACADDR_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(17),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_17_FFX_RST,
      O => macaddr(17)
    );
  macaddr_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_17_FFX_RST
    );
  mac_control_MACADDR_42 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(42),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_43_FFY_RST,
      O => macaddr(42)
    );
  macaddr_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_43_FFY_RST
    );
  mac_control_MACADDR_43 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(43),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_43_FFX_RST,
      O => macaddr(43)
    );
  macaddr_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_43_FFX_RST
    );
  mac_control_MACADDR_34 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(34),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_35_FFY_RST,
      O => macaddr(34)
    );
  macaddr_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_35_FFY_RST
    );
  mac_control_MACADDR_35 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(35),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_35_FFX_RST,
      O => macaddr(35)
    );
  macaddr_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_35_FFX_RST
    );
  mac_control_MACADDR_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(26),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_27_FFY_RST,
      O => macaddr(26)
    );
  macaddr_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_27_FFY_RST
    );
  mac_control_MACADDR_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(27),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_27_FFX_RST,
      O => macaddr(27)
    );
  macaddr_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_27_FFX_RST
    );
  mac_control_MACADDR_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(18),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_19_FFY_RST,
      O => macaddr(18)
    );
  macaddr_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_19_FFY_RST
    );
  mac_control_MACADDR_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(19),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_19_FFX_RST,
      O => macaddr(19)
    );
  macaddr_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_19_FFX_RST
    );
  mac_control_MACADDR_44 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(44),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_45_FFY_RST,
      O => macaddr(44)
    );
  macaddr_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_45_FFY_RST
    );
  mac_control_MACADDR_45 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(45),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_45_FFX_RST,
      O => macaddr(45)
    );
  macaddr_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_45_FFX_RST
    );
  mac_control_MACADDR_36 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(36),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_37_FFY_RST,
      O => macaddr(36)
    );
  macaddr_37_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_37_FFY_RST
    );
  mac_control_MACADDR_37 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(37),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_37_FFX_RST,
      O => macaddr(37)
    );
  macaddr_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_37_FFX_RST
    );
  mac_control_MACADDR_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(28),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_29_FFY_RST,
      O => macaddr(28)
    );
  macaddr_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_29_FFY_RST
    );
  mac_control_MACADDR_46 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(46),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_47_FFY_RST,
      O => macaddr(46)
    );
  macaddr_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_47_FFY_RST
    );
  mac_control_MACADDR_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(29),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_29_FFX_RST,
      O => macaddr(29)
    );
  macaddr_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_29_FFX_RST
    );
  tx_output_bpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(0),
      CE => tx_output_bpl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_1_FFY_RST,
      O => tx_output_bpl(0)
    );
  tx_output_bpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_1_FFY_RST
    );
  tx_output_bpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(1),
      CE => tx_output_bpl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_1_FFX_RST,
      O => tx_output_bpl(1)
    );
  tx_output_bpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_1_FFX_RST
    );
  tx_output_bpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(2),
      CE => tx_output_bpl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_3_FFY_RST,
      O => tx_output_bpl(2)
    );
  tx_output_bpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_3_FFY_RST
    );
  tx_output_bpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(3),
      CE => tx_output_bpl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_3_FFX_RST,
      O => tx_output_bpl(3)
    );
  tx_output_bpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_3_FFX_RST
    );
  tx_output_bpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(4),
      CE => tx_output_bpl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_5_FFY_RST,
      O => tx_output_bpl(4)
    );
  tx_output_bpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_5_FFY_RST
    );
  tx_output_bpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(5),
      CE => tx_output_bpl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_5_FFX_RST,
      O => tx_output_bpl(5)
    );
  tx_output_bpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_5_FFX_RST
    );
  tx_output_bpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(6),
      CE => tx_output_bpl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_7_FFY_RST,
      O => tx_output_bpl(6)
    );
  tx_output_bpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_7_FFY_RST
    );
  tx_output_bpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(7),
      CE => tx_output_bpl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_7_FFX_RST,
      O => tx_output_bpl(7)
    );
  tx_output_bpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_7_FFX_RST
    );
  tx_output_bpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(8),
      CE => tx_output_bpl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_9_FFY_RST,
      O => tx_output_bpl(8)
    );
  tx_output_bpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_9_FFY_RST
    );
  tx_output_bpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(9),
      CE => tx_output_bpl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_9_FFX_RST,
      O => tx_output_bpl(9)
    );
  tx_output_bpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_9_FFX_RST
    );
  mac_control_MACADDR_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(10),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_11_FFY_RST,
      O => macaddr(10)
    );
  macaddr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_11_FFY_RST
    );
  mac_control_MACADDR_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(20),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_21_FFY_RST,
      O => macaddr(20)
    );
  macaddr_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_21_FFY_RST
    );
  rx_input_memio_cs_FFd3_1985 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd3_FFY_RST,
      O => rx_input_memio_cs_FFd3
    );
  rx_input_memio_cs_FFd3_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd3_FFY_RST
    );
  rx_input_memio_cs_FFd4_1986 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd4_FFY_RST,
      O => rx_input_memio_cs_FFd4
    );
  rx_input_memio_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd4_FFY_RST
    );
  mac_control_MACADDR_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(11),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_11_FFX_RST,
      O => macaddr(11)
    );
  macaddr_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_11_FFX_RST
    );
  mac_control_MACADDR_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(21),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_21_FFX_RST,
      O => macaddr(21)
    );
  macaddr_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_21_FFX_RST
    );
  mac_control_MACADDR_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(12),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_13_FFY_RST,
      O => macaddr(12)
    );
  macaddr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_13_FFY_RST
    );
  mac_control_MACADDR_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(13),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_13_FFX_RST,
      O => macaddr(13)
    );
  macaddr_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_13_FFX_RST
    );
  mac_control_MACADDR_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(30),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_31_FFY_RST,
      O => macaddr(30)
    );
  macaddr_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_31_FFY_RST
    );
  mac_control_MACADDR_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(31),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_31_FFX_RST,
      O => macaddr(31)
    );
  macaddr_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_31_FFX_RST
    );
  mac_control_MACADDR_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(22),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_23_FFY_RST,
      O => macaddr(22)
    );
  macaddr_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_23_FFY_RST
    );
  mac_control_MACADDR_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(23),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_23_FFX_RST,
      O => macaddr(23)
    );
  macaddr_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_23_FFX_RST
    );
  mac_control_MACADDR_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(14),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_15_FFY_RST,
      O => macaddr(14)
    );
  macaddr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_15_FFY_RST
    );
  mac_control_MACADDR_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(15),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_15_FFX_RST,
      O => macaddr(15)
    );
  macaddr_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_15_FFX_RST
    );
  mac_control_MACADDR_40 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(40),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_41_FFY_RST,
      O => macaddr(40)
    );
  macaddr_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_41_FFY_RST
    );
  mac_control_MACADDR_41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(41),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_41_FFX_RST,
      O => macaddr(41)
    );
  macaddr_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_41_FFX_RST
    );
  mac_control_MACADDR_32 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(32),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_33_FFY_RST,
      O => macaddr(32)
    );
  macaddr_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_33_FFY_RST
    );
  mac_control_MACADDR_33 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(33),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_33_FFX_RST,
      O => macaddr(33)
    );
  macaddr_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_33_FFX_RST
    );
  mac_control_MACADDR_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(24),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_25_FFY_RST,
      O => macaddr(24)
    );
  macaddr_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_25_FFY_RST
    );
  mac_control_MACADDR_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(16),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_17_FFY_RST,
      O => macaddr(16)
    );
  macaddr_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_17_FFY_RST
    );
  mac_control_MACADDR_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(25),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_25_FFX_RST,
      O => macaddr(25)
    );
  macaddr_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_25_FFX_RST
    );
  mac_control_MACADDR_47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(47),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_47_FFX_RST,
      O => macaddr(47)
    );
  macaddr_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_47_FFX_RST
    );
  mac_control_MACADDR_38 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(38),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_39_FFY_RST,
      O => macaddr(38)
    );
  macaddr_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_39_FFY_RST
    );
  mac_control_MACADDR_39 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(39),
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_39_FFX_RST,
      O => macaddr(39)
    );
  macaddr_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_39_FFX_RST
    );
  mac_control_PHY_status_addrl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(0),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_addrl_1_FFY_RST,
      O => mac_control_PHY_status_addrl(0)
    );
  mac_control_PHY_status_addrl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_addrl_1_FFY_RST
    );
  mac_control_PHY_status_addrl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(1),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_addrl_1_FFX_RST,
      O => mac_control_PHY_status_addrl(1)
    );
  mac_control_PHY_status_addrl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_addrl_1_FFX_RST
    );
  mac_control_PHY_status_addrl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(3),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_addrl_3_FFX_RST,
      O => mac_control_PHY_status_addrl(3)
    );
  mac_control_PHY_status_addrl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_addrl_3_FFX_RST
    );
  tx_output_outsell_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_outsel_1_Q,
      CE => tx_output_outsell_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outsell_1_FFY_RST,
      O => tx_output_outsell(1)
    );
  tx_output_outsell_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outsell_1_FFY_RST
    );
  rx_input_memio_crcl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(17),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_17_FFY_RST,
      O => rx_input_memio_crcl(17)
    );
  rx_input_memio_crcl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_17_FFY_RST
    );
  slowclock_clkcnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_clkcnt_0_BXMUXNOT,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => slowclock_n0002,
      O => slowclock_clkcnt(0)
    );
  mac_control_phydi_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(20),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_21_FFY_RST,
      O => mac_control_phydi(20)
    );
  mac_control_phydi_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_21_FFY_RST
    );
  mac_control_phydi_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(21),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_21_FFX_RST,
      O => mac_control_phydi(21)
    );
  mac_control_phydi_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_21_FFX_RST
    );
  mac_control_phydi_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_13_FFY_RST,
      O => mac_control_phydi(12)
    );
  mac_control_phydi_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_13_FFY_RST
    );
  mac_control_phydi_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_13_FFX_RST,
      O => mac_control_phydi(13)
    );
  mac_control_phydi_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_13_FFX_RST
    );
  mac_control_phydi_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(30),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_31_FFY_RST,
      O => mac_control_phydi(30)
    );
  mac_control_phydi_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_31_FFY_RST
    );
  mac_control_phydi_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(31),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_31_FFX_RST,
      O => mac_control_phydi(31)
    );
  mac_control_phydi_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_31_FFX_RST
    );
  mac_control_phydi_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_15_FFY_RST,
      O => mac_control_phydi(14)
    );
  mac_control_phydi_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_15_FFY_RST
    );
  mac_control_phydi_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_15_FFX_RST,
      O => mac_control_phydi(15)
    );
  mac_control_phydi_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_15_FFX_RST
    );
  mac_control_phydi_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(22),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_23_FFY_RST,
      O => mac_control_phydi(22)
    );
  mac_control_phydi_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_23_FFY_RST
    );
  mac_control_phydi_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(23),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_23_FFX_RST,
      O => mac_control_phydi(23)
    );
  mac_control_phydi_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_23_FFX_RST
    );
  mac_control_phydi_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(16),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_17_FFY_RST,
      O => mac_control_phydi(16)
    );
  mac_control_phydi_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_17_FFY_RST
    );
  mac_control_phydi_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(17),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_17_FFX_RST,
      O => mac_control_phydi(17)
    );
  mac_control_phydi_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_17_FFX_RST
    );
  mac_control_phydi_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(24),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_25_FFY_RST,
      O => mac_control_phydi(24)
    );
  mac_control_phydi_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_25_FFY_RST
    );
  mac_control_phydi_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(25),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_25_FFX_RST,
      O => mac_control_phydi(25)
    );
  mac_control_phydi_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_25_FFX_RST
    );
  mac_control_phydi_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(18),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_19_FFY_RST,
      O => mac_control_phydi(18)
    );
  mac_control_phydi_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_19_FFY_RST
    );
  mac_control_din_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_Mshreg_sinlll_102,
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_1_FFY_RST,
      O => mac_control_din(0)
    );
  mac_control_din_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_1_FFY_RST
    );
  mac_control_din_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_1_FFX_RST,
      O => mac_control_din(1)
    );
  mac_control_din_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_1_FFX_RST
    );
  mac_control_din_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_3_FFY_RST,
      O => mac_control_din(2)
    );
  mac_control_din_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_3_FFY_RST
    );
  mac_control_din_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_3_FFX_RST,
      O => mac_control_din(3)
    );
  mac_control_din_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_3_FFX_RST
    );
  mac_control_din_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_5_FFY_RST,
      O => mac_control_din(4)
    );
  mac_control_din_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_5_FFY_RST
    );
  mac_control_din_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_5_FFX_RST,
      O => mac_control_din(5)
    );
  mac_control_din_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_5_FFX_RST
    );
  mac_control_din_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_7_FFY_RST,
      O => mac_control_din(6)
    );
  mac_control_din_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_7_FFY_RST
    );
  mac_control_din_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_7_FFX_RST,
      O => mac_control_din(7)
    );
  mac_control_din_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_7_FFX_RST
    );
  mac_control_din_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_9_FFY_RST,
      O => mac_control_din(8)
    );
  mac_control_din_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_9_FFY_RST
    );
  mac_control_din_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_din_9_FFX_RST,
      O => mac_control_din(9)
    );
  mac_control_din_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_9_FFX_RST
    );
  memcontroller_oel_1987 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel_BYMUXNOT,
      CE => memcontroller_oel_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_oel_FFY_RST,
      O => memcontroller_oel
    );
  memcontroller_oel_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_oel_FFY_RST
    );
  mac_control_phydi_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_11_FFY_RST,
      O => mac_control_phydi(10)
    );
  mac_control_phydi_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_11_FFY_RST
    );
  mac_control_phydi_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydi_11_FFX_RST,
      O => mac_control_phydi(11)
    );
  mac_control_phydi_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_11_FFX_RST
    );
  slowclock_clkcnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_clkcnt_n0000(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => slowclock_n0002,
      O => slowclock_clkcnt(1)
    );
  tx_output_FBBP_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(1),
      CE => txfbbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_1_FFX_RST,
      O => txfbbp(1)
    );
  txfbbp_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_1_FFX_RST
    );
  tx_output_FBBP_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(2),
      CE => txfbbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_3_FFY_RST,
      O => txfbbp(2)
    );
  txfbbp_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_3_FFY_RST
    );
  tx_output_FBBP_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(3),
      CE => txfbbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_3_FFX_RST,
      O => txfbbp(3)
    );
  txfbbp_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_3_FFX_RST
    );
  tx_output_FBBP_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(4),
      CE => txfbbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_5_FFY_RST,
      O => txfbbp(4)
    );
  txfbbp_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_5_FFY_RST
    );
  tx_output_FBBP_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(5),
      CE => txfbbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_5_FFX_RST,
      O => txfbbp(5)
    );
  txfbbp_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_5_FFX_RST
    );
  tx_output_FBBP_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(6),
      CE => txfbbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_7_FFY_RST,
      O => txfbbp(6)
    );
  txfbbp_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_7_FFY_RST
    );
  tx_output_FBBP_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(7),
      CE => txfbbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_7_FFX_RST,
      O => txfbbp(7)
    );
  txfbbp_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_7_FFX_RST
    );
  tx_output_FBBP_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(8),
      CE => txfbbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_9_FFY_RST,
      O => txfbbp(8)
    );
  txfbbp_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_9_FFY_RST
    );
  tx_output_FBBP_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(9),
      CE => txfbbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_9_FFX_RST,
      O => txfbbp(9)
    );
  txfbbp_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_9_FFX_RST
    );
  rx_input_memio_doutl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(10),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_11_FFY_RST,
      O => rx_input_memio_doutl(10)
    );
  rx_input_memio_doutl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_11_FFY_RST
    );
  rx_input_memio_doutl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(11),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_11_FFX_RST,
      O => rx_input_memio_doutl(11)
    );
  rx_input_memio_doutl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_11_FFX_RST
    );
  mac_control_lrxbcast_1988 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0026,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lrxbcast_FFY_RST,
      O => mac_control_lrxbcast
    );
  mac_control_lrxbcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lrxbcast_FFY_RST
    );
  rx_input_memio_doutl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(20),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_21_FFY_RST,
      O => rx_input_memio_doutl(20)
    );
  rx_input_memio_doutl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_21_FFY_RST
    );
  tx_fifocheck_bpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_11_FFX_RST,
      O => tx_fifocheck_bpl(11)
    );
  tx_fifocheck_bpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_11_FFX_RST
    );
  tx_fifocheck_bpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_13_FFX_RST,
      O => tx_fifocheck_bpl(13)
    );
  tx_fifocheck_bpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_13_FFX_RST
    );
  tx_fifocheck_bpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_13_FFY_RST,
      O => tx_fifocheck_bpl(12)
    );
  tx_fifocheck_bpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_13_FFY_RST
    );
  tx_fifocheck_bpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_15_FFY_RST,
      O => tx_fifocheck_bpl(14)
    );
  tx_fifocheck_bpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_15_FFY_RST
    );
  tx_fifocheck_bpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_15_FFX_RST,
      O => tx_fifocheck_bpl(15)
    );
  tx_fifocheck_bpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_15_FFX_RST
    );
  rx_output_lenr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(14),
      CE => rx_output_lenr_14_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_14_FFY_RST,
      O => rx_output_lenr(14)
    );
  rx_output_lenr_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_14_FFY_RST
    );
  rx_output_lenr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(15),
      CE => rx_output_lenr_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_15_FFY_RST,
      O => rx_output_lenr(15)
    );
  rx_output_lenr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_15_FFY_RST
    );
  tx_output_crcl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034(14),
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_14_FFY_RST,
      O => tx_output_crcl(14)
    );
  tx_output_crcl_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_14_FFY_RST
    );
  rx_input_memio_addrchk_rxmcastl_1989 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxmcast,
      CE => rx_input_memio_addrchk_rxmcastl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_rxmcastl_FFY_RST,
      O => rx_input_memio_addrchk_rxmcastl
    );
  rx_input_memio_addrchk_rxmcastl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_rxmcastl_FFY_RST
    );
  rx_input_memio_doutl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(21),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_21_FFX_RST,
      O => rx_input_memio_doutl(21)
    );
  rx_input_memio_doutl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_21_FFX_RST
    );
  rx_input_memio_doutl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(12),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_13_FFY_RST,
      O => rx_input_memio_doutl(12)
    );
  rx_input_memio_doutl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_13_FFY_RST
    );
  rx_input_memio_doutl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(13),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_13_FFX_RST,
      O => rx_input_memio_doutl(13)
    );
  rx_input_memio_doutl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_13_FFX_RST
    );
  rx_input_memio_doutl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(30),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_31_FFY_RST,
      O => rx_input_memio_doutl(30)
    );
  rx_input_memio_doutl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_31_FFY_RST
    );
  rx_input_memio_doutl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(31),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_31_FFX_RST,
      O => rx_input_memio_doutl(31)
    );
  rx_input_memio_doutl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_31_FFX_RST
    );
  rx_input_memio_doutl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(22),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_23_FFY_RST,
      O => rx_input_memio_doutl(22)
    );
  rx_input_memio_doutl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_23_FFY_RST
    );
  rx_input_memio_doutl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(23),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_23_FFX_RST,
      O => rx_input_memio_doutl(23)
    );
  rx_input_memio_doutl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_23_FFX_RST
    );
  rx_input_memio_doutl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(14),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_15_FFY_RST,
      O => rx_input_memio_doutl(14)
    );
  rx_input_memio_doutl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_15_FFY_RST
    );
  rx_input_memio_doutl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(15),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_15_FFX_RST,
      O => rx_input_memio_doutl(15)
    );
  rx_input_memio_doutl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_15_FFX_RST
    );
  rx_input_memio_doutl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(24),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_25_FFY_RST,
      O => rx_input_memio_doutl(24)
    );
  rx_input_memio_doutl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_25_FFY_RST
    );
  rx_input_memio_doutl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(25),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_25_FFX_RST,
      O => rx_input_memio_doutl(25)
    );
  rx_input_memio_doutl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_25_FFX_RST
    );
  rx_input_memio_doutl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(16),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_17_FFY_RST,
      O => rx_input_memio_doutl(16)
    );
  rx_input_memio_doutl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_17_FFY_RST
    );
  rx_input_memio_doutl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(17),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_17_FFX_RST,
      O => rx_input_memio_doutl(17)
    );
  rx_input_memio_doutl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_17_FFX_RST
    );
  rx_input_memio_doutl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(26),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_27_FFY_RST,
      O => rx_input_memio_doutl(26)
    );
  rx_input_memio_doutl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_27_FFY_RST
    );
  rx_input_memio_doutl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(27),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_27_FFX_RST,
      O => rx_input_memio_doutl(27)
    );
  rx_input_memio_doutl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_27_FFX_RST
    );
  rx_input_memio_doutl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(18),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_19_FFY_RST,
      O => rx_input_memio_doutl(18)
    );
  rx_input_memio_doutl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_19_FFY_RST
    );
  mac_control_PHY_status_din_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(11),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_11_FFX_RST,
      O => mac_control_PHY_status_din(11)
    );
  mac_control_PHY_status_din_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_11_FFX_RST
    );
  mac_control_PHY_status_din_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(12),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_13_FFY_RST,
      O => mac_control_PHY_status_din(12)
    );
  mac_control_PHY_status_din_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_13_FFY_RST
    );
  mac_control_PHY_status_din_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(13),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_13_FFX_RST,
      O => mac_control_PHY_status_din(13)
    );
  mac_control_PHY_status_din_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_13_FFX_RST
    );
  mac_control_PHY_status_din_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(14),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_15_FFY_RST,
      O => mac_control_PHY_status_din(14)
    );
  mac_control_PHY_status_din_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_15_FFY_RST
    );
  mac_control_PHY_status_din_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(15),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_15_FFX_RST,
      O => mac_control_PHY_status_din(15)
    );
  mac_control_PHY_status_din_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_15_FFX_RST
    );
  rx_input_memio_crcl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(18),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_18_FFY_RST,
      O => rx_input_memio_crcl(18)
    );
  rx_input_memio_crcl_18_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_18_FFY_RST
    );
  rx_input_memio_crcl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(26),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_26_FFY_RST,
      O => rx_input_memio_crcl(26)
    );
  rx_input_memio_crcl_26_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_26_FFY_RST
    );
  memcontroller_clknum_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_0_GROM,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_clknum_0_FFY_RST,
      O => memcontroller_clknum(1)
    );
  memcontroller_clknum_0_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_0_FFY_RST
    );
  tx_output_FBBP_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(0),
      CE => txfbbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_1_FFY_RST,
      O => txfbbp(0)
    );
  txfbbp_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_1_FFY_RST
    );
  slowclock_rxfifowerrl_1990 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_rxfifowerrl_GROM,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => rxfifowerr,
      SRST => slowclock_rxfifowerrl_LOGIC_ZERO,
      O => slowclock_rxfifowerrl
    );
  memcontroller_clknum_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_0_BXMUXNOT,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_clknum_0_FFX_RST,
      O => memcontroller_clknum(0)
    );
  memcontroller_clknum_0_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_0_FFX_RST
    );
  rx_input_fifo_control_d2_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(6),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_7_FFY_RST,
      O => rx_input_fifo_control_d2(6)
    );
  rx_input_fifo_control_d2_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_7_FFY_RST
    );
  rx_input_fifo_control_d2_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(7),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_7_FFX_RST,
      O => rx_input_fifo_control_d2(7)
    );
  rx_input_fifo_control_d2_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_7_FFX_RST
    );
  rx_input_fifo_control_d3_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(2),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_3_FFY_RST,
      O => rx_input_fifo_control_d3(2)
    );
  rx_input_fifo_control_d3_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_3_FFY_RST
    );
  rx_input_fifo_control_d3_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(3),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_3_FFX_RST,
      O => rx_input_fifo_control_d3(3)
    );
  rx_input_fifo_control_d3_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_3_FFX_RST
    );
  rx_input_fifo_control_d3_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(4),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_5_FFY_RST,
      O => rx_input_fifo_control_d3(4)
    );
  rx_input_fifo_control_d3_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_5_FFY_RST
    );
  rx_input_fifo_control_d2_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(8),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_8_FFY_RST,
      O => rx_input_fifo_control_d2(8)
    );
  rx_input_fifo_control_d2_8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_8_FFY_RST
    );
  rx_input_fifo_control_d3_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(5),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_5_FFX_RST,
      O => rx_input_fifo_control_d3(5)
    );
  rx_input_fifo_control_d3_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_5_FFX_RST
    );
  rx_input_fifo_control_d2_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1_9_rt,
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_control_d2_9_FFY_SET,
      RST => rx_input_fifo_control_d2_9_FFY_RST,
      O => rx_input_fifo_control_d2(9)
    );
  rx_input_fifo_control_d2_9_FFY_SETOR : X_BUF
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_d2_9_FFY_SET
    );
  rx_input_fifo_control_d2_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_control_d2_9_LOGIC_ZERO,
      I1 => GSR,
      O => rx_input_fifo_control_d2_9_FFY_RST
    );
  rx_input_fifo_control_d3_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(6),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_7_FFY_RST,
      O => rx_input_fifo_control_d3(6)
    );
  rx_input_fifo_control_d3_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_7_FFY_RST
    );
  rx_input_fifo_control_d3_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(7),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_7_FFX_RST,
      O => rx_input_fifo_control_d3(7)
    );
  rx_input_fifo_control_d3_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_7_FFX_RST
    );
  rx_input_fifo_control_d3_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2_9_rt,
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_control_d3_9_FFY_SET,
      RST => rx_input_fifo_control_d3_9_FFY_RST,
      O => rx_input_fifo_control_d3(9)
    );
  rx_input_fifo_control_d3_9_FFY_SETOR : X_BUF
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_d3_9_FFY_SET
    );
  rx_input_fifo_control_d3_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_control_d3_9_LOGIC_ZERO,
      I1 => GSR,
      O => rx_input_fifo_control_d3_9_FFY_RST
    );
  rx_input_fifo_control_d3_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(8),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_8_FFY_RST,
      O => rx_input_fifo_control_d3(8)
    );
  rx_input_fifo_control_d3_8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_8_FFY_RST
    );
  tx_input_MD_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(13),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_13_FFX_RST,
      O => d4(13)
    );
  d4_13_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_13_FFX_RST
    );
  tx_input_MD_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(7),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_23_FFX_RST,
      O => d4(23)
    );
  d4_23_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_23_FFX_RST
    );
  tx_input_MD_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(14),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_15_FFY_RST,
      O => d4(14)
    );
  d4_15_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_15_FFY_RST
    );
  tx_input_MD_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(15),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_15_FFX_RST,
      O => d4(15)
    );
  d4_15_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_15_FFX_RST
    );
  tx_input_MD_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(14),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_31_FFY_RST,
      O => d4(30)
    );
  d4_31_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_31_FFY_RST
    );
  tx_input_MD_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(15),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_31_FFX_RST,
      O => d4(31)
    );
  d4_31_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_31_FFX_RST
    );
  tx_input_MD_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(0),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_17_FFY_RST,
      O => d4(16)
    );
  d4_17_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_17_FFY_RST
    );
  tx_input_MD_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(1),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_17_FFX_RST,
      O => d4(17)
    );
  d4_17_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_17_FFX_RST
    );
  tx_input_MD_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(8),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_25_FFY_RST,
      O => d4(24)
    );
  d4_25_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_25_FFY_RST
    );
  tx_input_MD_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(9),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_25_FFX_RST,
      O => d4(25)
    );
  d4_25_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_25_FFX_RST
    );
  tx_input_MD_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(2),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_19_FFY_RST,
      O => d4(18)
    );
  d4_19_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_19_FFY_RST
    );
  tx_input_MD_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(3),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_19_FFX_RST,
      O => d4(19)
    );
  d4_19_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_19_FFX_RST
    );
  tx_input_MD_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(10),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_27_FFY_RST,
      O => d4(26)
    );
  d4_27_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_27_FFY_RST
    );
  tx_input_MD_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(11),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_27_FFX_RST,
      O => d4(27)
    );
  d4_27_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_27_FFX_RST
    );
  rx_input_fifo_control_cel : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_rd_en_GROM,
      CE => rx_input_fifo_rd_en_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_rd_en_FFY_RST,
      O => rx_input_fifo_rd_en
    );
  rx_input_fifo_rd_en_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_rd_en_FFY_RST
    );
  tx_input_MD_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(12),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_29_FFY_RST,
      O => d4(28)
    );
  d4_29_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_29_FFY_RST
    );
  rx_input_fifo_control_d1_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(5),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_5_FFX_RST,
      O => rx_input_fifo_control_d1(5)
    );
  rx_input_fifo_control_d1_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_5_FFX_RST
    );
  rx_input_fifo_control_d2_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(0),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_1_FFY_RST,
      O => rx_input_fifo_control_d2(0)
    );
  rx_input_fifo_control_d2_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_1_FFY_RST
    );
  rx_input_fifo_control_d2_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(1),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_1_FFX_RST,
      O => rx_input_fifo_control_d2(1)
    );
  rx_input_fifo_control_d2_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_1_FFX_RST
    );
  rx_input_fifo_control_d0_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl_9_rt,
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_control_d0_9_FFY_SET,
      RST => rx_input_fifo_control_d0_9_FFY_RST,
      O => rx_input_fifo_control_d0(9)
    );
  rx_input_fifo_control_d0_9_FFY_SETOR : X_BUF
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_d0_9_FFY_SET
    );
  rx_input_fifo_control_d0_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_control_d0_9_LOGIC_ZERO,
      I1 => GSR,
      O => rx_input_fifo_control_d0_9_FFY_RST
    );
  rx_input_fifo_control_d1_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(6),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_7_FFY_RST,
      O => rx_input_fifo_control_d1(6)
    );
  rx_input_fifo_control_d1_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_7_FFY_RST
    );
  rx_input_fifo_control_d1_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(7),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_7_FFX_RST,
      O => rx_input_fifo_control_d1(7)
    );
  rx_input_fifo_control_d1_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_7_FFX_RST
    );
  rx_input_fifo_control_d2_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(2),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_3_FFY_RST,
      O => rx_input_fifo_control_d2(2)
    );
  rx_input_fifo_control_d2_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_3_FFY_RST
    );
  rx_input_fifo_control_d2_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(3),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_3_FFX_RST,
      O => rx_input_fifo_control_d2(3)
    );
  rx_input_fifo_control_d2_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_3_FFX_RST
    );
  rx_input_fifo_control_d2_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(4),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_5_FFY_RST,
      O => rx_input_fifo_control_d2(4)
    );
  rx_input_fifo_control_d2_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_5_FFY_RST
    );
  rx_input_fifo_control_d1_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(8),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_8_FFY_RST,
      O => rx_input_fifo_control_d1(8)
    );
  rx_input_fifo_control_d1_8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_8_FFY_RST
    );
  rx_input_fifo_control_d2_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(5),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_5_FFX_RST,
      O => rx_input_fifo_control_d2(5)
    );
  rx_input_fifo_control_d2_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_5_FFX_RST
    );
  rx_input_fifo_control_d1_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0_9_rt,
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_control_d1_9_FFY_SET,
      RST => rx_input_fifo_control_d1_9_FFY_RST,
      O => rx_input_fifo_control_d1(9)
    );
  rx_input_fifo_control_d1_9_FFY_SETOR : X_BUF
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_d1_9_FFY_SET
    );
  rx_input_fifo_control_d1_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_control_d1_9_LOGIC_ZERO,
      I1 => GSR,
      O => rx_input_fifo_control_d1_9_FFY_RST
    );
  rx_input_fifo_control_d3_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(0),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_1_FFY_RST,
      O => rx_input_fifo_control_d3(0)
    );
  rx_input_fifo_control_d3_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_1_FFY_RST
    );
  rx_input_fifo_control_d3_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(1),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_1_FFX_RST,
      O => rx_input_fifo_control_d3(1)
    );
  rx_input_fifo_control_d3_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_1_FFX_RST
    );
  rx_input_memio_crcl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(27),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_27_FFY_RST,
      O => rx_input_memio_crcl(27)
    );
  rx_input_memio_crcl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_27_FFY_RST
    );
  mac_control_lrxmcast_1991 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lrxmcast_FFY_RST,
      O => mac_control_lrxmcast
    );
  mac_control_lrxmcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lrxmcast_FFY_RST
    );
  rx_input_GMII_rx_dvll_1992 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_rx_dvl,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_GMII_rx_dvll_FFY_RST,
      O => rx_input_GMII_rx_dvll
    );
  rx_input_GMII_rx_dvll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_GMII_rx_dvll_FFY_RST
    );
  mac_control_lrxucast_1993 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_lrxucast_FFY_RST,
      O => mac_control_lrxucast
    );
  mac_control_lrxucast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lrxucast_FFY_RST
    );
  rx_input_fifo_control_cell_1994 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_rd_en,
      CE => rx_input_fifo_control_cell_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_cell_FFY_RST,
      O => rx_input_fifo_control_cell
    );
  rx_input_fifo_control_cell_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_cell_FFY_RST
    );
  rx_input_memio_crcl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(28),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_28_FFY_RST,
      O => rx_input_memio_crcl(28)
    );
  rx_input_memio_crcl_28_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_28_FFY_RST
    );
  rx_input_memio_crcl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048(14),
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_14_FFY_RST,
      O => rx_input_memio_crcl(14)
    );
  rx_input_memio_crcl_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_14_FFY_RST
    );
  rx_input_memio_addrchk_validmcast_1995 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_mcast(0),
      CE => rx_input_memio_addrchk_validmcast_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_validmcast_FFY_RST,
      O => rx_input_memio_addrchk_validmcast
    );
  rx_input_memio_addrchk_validmcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_validmcast_FFY_RST
    );
  mac_control_ledtx_rst_1996 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cross,
      CE => mac_control_N52198,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_ledtx_rst_FFY_RST,
      O => mac_control_ledtx_rst
    );
  mac_control_ledtx_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_rst_FFY_RST
    );
  tx_input_MA_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_26,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_11_FFY_RST,
      O => addr4ext(10)
    );
  addr4ext_11_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_11_FFY_RST
    );
  tx_input_MA_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_27,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_11_FFX_RST,
      O => addr4ext(11)
    );
  addr4ext_11_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_11_FFX_RST
    );
  tx_input_MA_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_28,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_13_FFY_RST,
      O => addr4ext(12)
    );
  addr4ext_13_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_13_FFY_RST
    );
  tx_input_MA_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_29,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_13_FFX_RST,
      O => addr4ext(13)
    );
  addr4ext_13_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_13_FFX_RST
    );
  tx_input_MA_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_30,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_15_FFY_RST,
      O => addr4ext(14)
    );
  addr4ext_15_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_15_FFY_RST
    );
  tx_input_MA_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_31,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_15_FFX_RST,
      O => addr4ext(15)
    );
  addr4ext_15_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_15_FFX_RST
    );
  tx_input_MD_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(10),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_11_FFY_RST,
      O => d4(10)
    );
  d4_11_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_11_FFY_RST
    );
  tx_input_MD_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(11),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_11_FFX_RST,
      O => d4(11)
    );
  d4_11_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_11_FFX_RST
    );
  mac_control_RXALLF : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lrxallf,
      CE => clkslen,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxallf_FFY_RST,
      O => rxallf
    );
  rxallf_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxallf_FFY_RST
    );
  tx_input_MD_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(4),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_21_FFY_RST,
      O => d4(20)
    );
  d4_21_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_21_FFY_RST
    );
  tx_input_MD_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(5),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_21_FFX_RST,
      O => d4(21)
    );
  d4_21_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_21_FFX_RST
    );
  tx_input_MD_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(6),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_23_FFY_RST,
      O => d4(22)
    );
  d4_23_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_23_FFY_RST
    );
  tx_input_MD_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(12),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_13_FFY_RST,
      O => d4(12)
    );
  d4_13_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_13_FFY_RST
    );
  tx_input_MD_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(13),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_29_FFX_RST,
      O => d4(29)
    );
  d4_29_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_29_FFX_RST
    );
  rx_fifocheck_FIFOFULL : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfifofull_LOGIC_ONE,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_fifocheck_N74128,
      O => rxfifofull
    );
  rx_input_memio_addrchk_rxbcastl_1997 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbcast,
      CE => rx_input_memio_addrchk_rxbcastl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_rxbcastl_FFY_RST,
      O => rx_input_memio_addrchk_rxbcastl
    );
  rx_input_memio_addrchk_rxbcastl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_rxbcastl_FFY_RST
    );
  slowclock_clken : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => slowclock_lclken,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => clkslen_FFY_RST,
      O => clkslen
    );
  clkslen_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => clkslen_FFY_RST
    );
  rx_output_lenr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(10),
      CE => rx_output_lenr_10_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_10_FFY_RST,
      O => rx_output_lenr(10)
    );
  rx_output_lenr_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_10_FFY_RST
    );
  rx_output_lenr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(11),
      CE => rx_output_lenr_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_11_FFY_RST,
      O => rx_output_lenr(11)
    );
  rx_output_lenr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_11_FFY_RST
    );
  rx_output_lenr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(12),
      CE => rx_output_lenr_12_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_12_FFY_RST,
      O => rx_output_lenr(12)
    );
  rx_output_lenr_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_12_FFY_RST
    );
  tx_fifocheck_bpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_11_FFY_RST,
      O => tx_fifocheck_bpl(10)
    );
  tx_fifocheck_bpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_11_FFY_RST
    );
  rx_output_lenr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046(13),
      CE => rx_output_lenr_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_13_FFY_RST,
      O => rx_output_lenr(13)
    );
  rx_output_lenr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_13_FFY_RST
    );
  rx_input_fifo_control_dinl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(0),
      CE => rx_input_fifo_control_dinl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_1_FFY_RST,
      O => rx_input_fifo_control_dinl(0)
    );
  rx_input_fifo_control_dinl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_1_FFY_RST
    );
  rx_input_fifo_control_dinl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(1),
      CE => rx_input_fifo_control_dinl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_1_FFX_RST,
      O => rx_input_fifo_control_dinl(1)
    );
  rx_input_fifo_control_dinl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_1_FFX_RST
    );
  rx_input_fifo_control_dinl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(2),
      CE => rx_input_fifo_control_dinl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_3_FFY_RST,
      O => rx_input_fifo_control_dinl(2)
    );
  rx_input_fifo_control_dinl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_3_FFY_RST
    );
  rx_input_fifo_control_dinl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(3),
      CE => rx_input_fifo_control_dinl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_3_FFX_RST,
      O => rx_input_fifo_control_dinl(3)
    );
  rx_input_fifo_control_dinl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_3_FFX_RST
    );
  rx_input_fifo_control_dinl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(4),
      CE => rx_input_fifo_control_dinl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_5_FFY_RST,
      O => rx_input_fifo_control_dinl(4)
    );
  rx_input_fifo_control_dinl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_5_FFY_RST
    );
  rx_input_fifo_control_dinl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(5),
      CE => rx_input_fifo_control_dinl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_5_FFX_RST,
      O => rx_input_fifo_control_dinl(5)
    );
  rx_input_fifo_control_dinl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_5_FFX_RST
    );
  rx_input_fifo_control_dinl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(6),
      CE => rx_input_fifo_control_dinl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_7_FFY_RST,
      O => rx_input_fifo_control_dinl(6)
    );
  rx_input_fifo_control_dinl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_7_FFY_RST
    );
  rx_input_fifo_control_dinl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(7),
      CE => rx_input_fifo_control_dinl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_7_FFX_RST,
      O => rx_input_fifo_control_dinl(7)
    );
  rx_input_fifo_control_dinl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_7_FFX_RST
    );
  CLKIN_BUF : X_CKBUF
    port map (
      I => CLKIN,
      O => CLKIN_IBUFG
    );
  RX_CLK_BUF : X_CKBUF
    port map (
      I => RX_CLK,
      O => RX_CLK_IBUFG
    );
  CLKIOIN_BUF : X_CKBUF
    port map (
      I => CLKIOIN,
      O => CLKIOIN_IBUFG
    );
  clkio_bufg_BUF : X_CKBUF
    port map (
      I => clkio_to_bufg,
      O => clkio
    );
  clk_bufg_BUF : X_CKBUF
    port map (
      I => clk_to_bufg,
      O => GTX_CLK_OBUF
    );
  clkrx_bufg_BUF : X_CKBUF
    port map (
      I => clkrx_to_bufg,
      O => clkrx
    );
  PWR_VCC_0_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_0_FROM
    );
  PWR_VCC_0_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_0_GROM
    );
  PWR_VCC_0_XUSED : X_BUF
    port map (
      I => PWR_VCC_0_FROM,
      O => GLOBAL_LOGIC1
    );
  PWR_VCC_0_YUSED : X_BUF
    port map (
      I => PWR_VCC_0_GROM,
      O => GLOBAL_LOGIC0_0
    );
  PWR_VCC_1_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_1_FROM
    );
  PWR_VCC_1_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_1_GROM
    );
  PWR_VCC_1_XUSED : X_BUF
    port map (
      I => PWR_VCC_1_FROM,
      O => GLOBAL_LOGIC1_0
    );
  PWR_VCC_1_YUSED : X_BUF
    port map (
      I => PWR_VCC_1_GROM,
      O => GLOBAL_LOGIC0_57
    );
  PWR_VCC_2_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_2_FROM
    );
  PWR_VCC_2_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_2_GROM
    );
  PWR_VCC_2_XUSED : X_BUF
    port map (
      I => PWR_VCC_2_FROM,
      O => GLOBAL_LOGIC1_1
    );
  PWR_VCC_2_YUSED : X_BUF
    port map (
      I => PWR_VCC_2_GROM,
      O => GLOBAL_LOGIC0_56
    );
  PWR_VCC_3_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_3_FROM
    );
  PWR_VCC_3_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_3_GROM
    );
  PWR_VCC_3_XUSED : X_BUF
    port map (
      I => PWR_VCC_3_FROM,
      O => GLOBAL_LOGIC1_2
    );
  PWR_VCC_3_YUSED : X_BUF
    port map (
      I => PWR_VCC_3_GROM,
      O => GLOBAL_LOGIC0_6
    );
  PWR_VCC_4_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_4_FROM
    );
  PWR_VCC_4_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_4_GROM
    );
  PWR_VCC_4_XUSED : X_BUF
    port map (
      I => PWR_VCC_4_FROM,
      O => GLOBAL_LOGIC1_3
    );
  PWR_VCC_4_YUSED : X_BUF
    port map (
      I => PWR_VCC_4_GROM,
      O => GLOBAL_LOGIC0_8
    );
  PWR_VCC_5_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_5_FROM
    );
  PWR_VCC_5_XUSED : X_BUF
    port map (
      I => PWR_VCC_5_FROM,
      O => GLOBAL_LOGIC1_4
    );
  PWR_VCC_6_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_6_FROM
    );
  PWR_VCC_6_XUSED : X_BUF
    port map (
      I => PWR_VCC_6_FROM,
      O => GLOBAL_LOGIC1_5
    );
  PWR_VCC_7_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_7_FROM
    );
  PWR_VCC_7_XUSED : X_BUF
    port map (
      I => PWR_VCC_7_FROM,
      O => GLOBAL_LOGIC1_6
    );
  PWR_VCC_8_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_8_FROM
    );
  PWR_VCC_8_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_8_GROM
    );
  PWR_VCC_8_XUSED : X_BUF
    port map (
      I => PWR_VCC_8_FROM,
      O => GLOBAL_LOGIC1_7
    );
  PWR_VCC_8_YUSED : X_BUF
    port map (
      I => PWR_VCC_8_GROM,
      O => GLOBAL_LOGIC0_47
    );
  PWR_VCC_9_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_9_FROM
    );
  PWR_VCC_9_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_9_GROM
    );
  PWR_VCC_9_XUSED : X_BUF
    port map (
      I => PWR_VCC_9_FROM,
      O => GLOBAL_LOGIC1_8
    );
  PWR_VCC_9_YUSED : X_BUF
    port map (
      I => PWR_VCC_9_GROM,
      O => GLOBAL_LOGIC0_46
    );
  PWR_VCC_10_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_10_FROM
    );
  PWR_VCC_10_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_10_GROM
    );
  PWR_VCC_10_XUSED : X_BUF
    port map (
      I => PWR_VCC_10_FROM,
      O => GLOBAL_LOGIC1_9
    );
  PWR_VCC_10_YUSED : X_BUF
    port map (
      I => PWR_VCC_10_GROM,
      O => GLOBAL_LOGIC0_45
    );
  PWR_VCC_11_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_11_FROM
    );
  PWR_VCC_11_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_11_GROM
    );
  PWR_VCC_11_XUSED : X_BUF
    port map (
      I => PWR_VCC_11_FROM,
      O => GLOBAL_LOGIC1_10
    );
  PWR_VCC_11_YUSED : X_BUF
    port map (
      I => PWR_VCC_11_GROM,
      O => GLOBAL_LOGIC0_44
    );
  PWR_VCC_12_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_12_FROM
    );
  PWR_VCC_12_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_12_GROM
    );
  PWR_VCC_12_XUSED : X_BUF
    port map (
      I => PWR_VCC_12_FROM,
      O => GLOBAL_LOGIC1_11
    );
  PWR_VCC_12_YUSED : X_BUF
    port map (
      I => PWR_VCC_12_GROM,
      O => GLOBAL_LOGIC0_43
    );
  PWR_VCC_13_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_13_FROM
    );
  PWR_VCC_13_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_13_GROM
    );
  PWR_VCC_13_XUSED : X_BUF
    port map (
      I => PWR_VCC_13_FROM,
      O => GLOBAL_LOGIC1_12
    );
  PWR_VCC_13_YUSED : X_BUF
    port map (
      I => PWR_VCC_13_GROM,
      O => GLOBAL_LOGIC0_42
    );
  PWR_VCC_14_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_14_FROM
    );
  PWR_VCC_14_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_14_GROM
    );
  PWR_VCC_14_XUSED : X_BUF
    port map (
      I => PWR_VCC_14_FROM,
      O => GLOBAL_LOGIC1_13
    );
  PWR_VCC_14_YUSED : X_BUF
    port map (
      I => PWR_VCC_14_GROM,
      O => GLOBAL_LOGIC0_41
    );
  PWR_VCC_15_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_15_FROM
    );
  PWR_VCC_15_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_15_GROM
    );
  PWR_VCC_15_XUSED : X_BUF
    port map (
      I => PWR_VCC_15_FROM,
      O => GLOBAL_LOGIC1_14
    );
  PWR_VCC_15_YUSED : X_BUF
    port map (
      I => PWR_VCC_15_GROM,
      O => GLOBAL_LOGIC0_40
    );
  PWR_VCC_16_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_16_FROM
    );
  PWR_VCC_16_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_16_GROM
    );
  PWR_VCC_16_XUSED : X_BUF
    port map (
      I => PWR_VCC_16_FROM,
      O => GLOBAL_LOGIC1_15
    );
  PWR_VCC_16_YUSED : X_BUF
    port map (
      I => PWR_VCC_16_GROM,
      O => GLOBAL_LOGIC0_39
    );
  PWR_VCC_17_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_17_FROM
    );
  PWR_VCC_17_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_17_GROM
    );
  PWR_VCC_17_XUSED : X_BUF
    port map (
      I => PWR_VCC_17_FROM,
      O => GLOBAL_LOGIC1_16
    );
  PWR_VCC_17_YUSED : X_BUF
    port map (
      I => PWR_VCC_17_GROM,
      O => GLOBAL_LOGIC0_36
    );
  PWR_VCC_18_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_18_FROM
    );
  PWR_VCC_18_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_18_GROM
    );
  PWR_VCC_18_XUSED : X_BUF
    port map (
      I => PWR_VCC_18_FROM,
      O => GLOBAL_LOGIC1_17
    );
  PWR_VCC_18_YUSED : X_BUF
    port map (
      I => PWR_VCC_18_GROM,
      O => GLOBAL_LOGIC0_33
    );
  PWR_VCC_19_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_19_FROM
    );
  PWR_VCC_19_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_19_GROM
    );
  PWR_VCC_19_XUSED : X_BUF
    port map (
      I => PWR_VCC_19_FROM,
      O => GLOBAL_LOGIC1_18
    );
  PWR_VCC_19_YUSED : X_BUF
    port map (
      I => PWR_VCC_19_GROM,
      O => GLOBAL_LOGIC0_31
    );
  PWR_VCC_20_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_20_FROM
    );
  PWR_VCC_20_XUSED : X_BUF
    port map (
      I => PWR_VCC_20_FROM,
      O => GLOBAL_LOGIC1_19
    );
  PWR_VCC_21_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_21_FROM
    );
  PWR_VCC_21_XUSED : X_BUF
    port map (
      I => PWR_VCC_21_FROM,
      O => GLOBAL_LOGIC1_20
    );
  PWR_VCC_22_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_22_FROM
    );
  PWR_VCC_22_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_22_GROM
    );
  PWR_VCC_22_XUSED : X_BUF
    port map (
      I => PWR_VCC_22_FROM,
      O => GLOBAL_LOGIC1_21
    );
  PWR_VCC_22_YUSED : X_BUF
    port map (
      I => PWR_VCC_22_GROM,
      O => GLOBAL_LOGIC0_27
    );
  PWR_VCC_23_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_23_FROM
    );
  PWR_VCC_23_XUSED : X_BUF
    port map (
      I => PWR_VCC_23_FROM,
      O => GLOBAL_LOGIC1_22
    );
  PWR_VCC_24_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_24_FROM
    );
  PWR_VCC_24_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_24_GROM
    );
  PWR_VCC_24_XUSED : X_BUF
    port map (
      I => PWR_VCC_24_FROM,
      O => GLOBAL_LOGIC1_23
    );
  PWR_VCC_24_YUSED : X_BUF
    port map (
      I => PWR_VCC_24_GROM,
      O => GLOBAL_LOGIC0_26
    );
  PWR_VCC_25_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_25_FROM
    );
  PWR_VCC_25_XUSED : X_BUF
    port map (
      I => PWR_VCC_25_FROM,
      O => GLOBAL_LOGIC1_24
    );
  PWR_VCC_26_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_26_FROM
    );
  PWR_VCC_26_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_26_GROM
    );
  PWR_VCC_26_XUSED : X_BUF
    port map (
      I => PWR_VCC_26_FROM,
      O => GLOBAL_LOGIC1_25
    );
  PWR_VCC_26_YUSED : X_BUF
    port map (
      I => PWR_VCC_26_GROM,
      O => GLOBAL_LOGIC0_25
    );
  PWR_VCC_27_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_27_FROM
    );
  PWR_VCC_27_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_27_GROM
    );
  PWR_VCC_27_XUSED : X_BUF
    port map (
      I => PWR_VCC_27_FROM,
      O => GLOBAL_LOGIC1_26
    );
  PWR_VCC_27_YUSED : X_BUF
    port map (
      I => PWR_VCC_27_GROM,
      O => GLOBAL_LOGIC0_23
    );
  PWR_VCC_28_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_28_FROM
    );
  PWR_VCC_28_XUSED : X_BUF
    port map (
      I => PWR_VCC_28_FROM,
      O => GLOBAL_LOGIC1_27
    );
  PWR_VCC_29_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_29_FROM
    );
  PWR_VCC_29_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_29_GROM
    );
  PWR_VCC_29_XUSED : X_BUF
    port map (
      I => PWR_VCC_29_FROM,
      O => GLOBAL_LOGIC1_28
    );
  PWR_VCC_29_YUSED : X_BUF
    port map (
      I => PWR_VCC_29_GROM,
      O => GLOBAL_LOGIC0_21
    );
  PWR_VCC_30_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_30_FROM
    );
  PWR_VCC_30_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_30_GROM
    );
  PWR_VCC_30_XUSED : X_BUF
    port map (
      I => PWR_VCC_30_FROM,
      O => GLOBAL_LOGIC1_29
    );
  PWR_VCC_30_YUSED : X_BUF
    port map (
      I => PWR_VCC_30_GROM,
      O => GLOBAL_LOGIC0_20
    );
  PWR_VCC_31_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_31_FROM
    );
  PWR_VCC_31_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_31_GROM
    );
  PWR_VCC_31_XUSED : X_BUF
    port map (
      I => PWR_VCC_31_FROM,
      O => GLOBAL_LOGIC1_30
    );
  PWR_VCC_31_YUSED : X_BUF
    port map (
      I => PWR_VCC_31_GROM,
      O => GLOBAL_LOGIC0_18
    );
  PWR_VCC_32_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_32_FROM
    );
  PWR_VCC_32_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_32_GROM
    );
  PWR_VCC_32_XUSED : X_BUF
    port map (
      I => PWR_VCC_32_FROM,
      O => GLOBAL_LOGIC1_31
    );
  PWR_VCC_32_YUSED : X_BUF
    port map (
      I => PWR_VCC_32_GROM,
      O => GLOBAL_LOGIC0_17
    );
  PWR_VCC_33_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_33_FROM
    );
  PWR_VCC_33_XUSED : X_BUF
    port map (
      I => PWR_VCC_33_FROM,
      O => GLOBAL_LOGIC1_32
    );
  PWR_VCC_34_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_34_FROM
    );
  PWR_VCC_34_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_34_GROM
    );
  PWR_VCC_34_XUSED : X_BUF
    port map (
      I => PWR_VCC_34_FROM,
      O => GLOBAL_LOGIC1_33
    );
  PWR_VCC_34_YUSED : X_BUF
    port map (
      I => PWR_VCC_34_GROM,
      O => GLOBAL_LOGIC0_16
    );
  PWR_VCC_35_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_35_FROM
    );
  PWR_VCC_35_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_35_GROM
    );
  PWR_VCC_35_XUSED : X_BUF
    port map (
      I => PWR_VCC_35_FROM,
      O => GLOBAL_LOGIC1_34
    );
  PWR_VCC_35_YUSED : X_BUF
    port map (
      I => PWR_VCC_35_GROM,
      O => GLOBAL_LOGIC0_15
    );
  PWR_VCC_36_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_36_FROM
    );
  PWR_VCC_36_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_36_GROM
    );
  PWR_VCC_36_XUSED : X_BUF
    port map (
      I => PWR_VCC_36_FROM,
      O => GLOBAL_LOGIC1_35
    );
  PWR_VCC_36_YUSED : X_BUF
    port map (
      I => PWR_VCC_36_GROM,
      O => GLOBAL_LOGIC0_10
    );
  PWR_VCC_37_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_37_FROM
    );
  PWR_VCC_37_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_37_GROM
    );
  PWR_VCC_37_XUSED : X_BUF
    port map (
      I => PWR_VCC_37_FROM,
      O => GLOBAL_LOGIC1_36
    );
  PWR_VCC_37_YUSED : X_BUF
    port map (
      I => PWR_VCC_37_GROM,
      O => GLOBAL_LOGIC0_2
    );
  PWR_VCC_38_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_38_FROM
    );
  PWR_VCC_38_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_38_GROM
    );
  PWR_VCC_38_XUSED : X_BUF
    port map (
      I => PWR_VCC_38_FROM,
      O => GLOBAL_LOGIC1_37
    );
  PWR_VCC_38_YUSED : X_BUF
    port map (
      I => PWR_VCC_38_GROM,
      O => GLOBAL_LOGIC0_1
    );
  PWR_GND_0_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_0_GROM
    );
  PWR_GND_0_YUSED : X_BUF
    port map (
      I => PWR_GND_0_GROM,
      O => GLOBAL_LOGIC0
    );
  PWR_GND_1_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_1_GROM
    );
  PWR_GND_1_YUSED : X_BUF
    port map (
      I => PWR_GND_1_GROM,
      O => GLOBAL_LOGIC0_3
    );
  PWR_GND_2_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_2_GROM
    );
  PWR_GND_2_YUSED : X_BUF
    port map (
      I => PWR_GND_2_GROM,
      O => GLOBAL_LOGIC0_4
    );
  PWR_GND_3_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_3_GROM
    );
  PWR_GND_3_YUSED : X_BUF
    port map (
      I => PWR_GND_3_GROM,
      O => GLOBAL_LOGIC0_5
    );
  PWR_GND_4_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_4_GROM
    );
  PWR_GND_4_YUSED : X_BUF
    port map (
      I => PWR_GND_4_GROM,
      O => GLOBAL_LOGIC0_7
    );
  PWR_GND_5_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_5_GROM
    );
  PWR_GND_5_YUSED : X_BUF
    port map (
      I => PWR_GND_5_GROM,
      O => GLOBAL_LOGIC0_9
    );
  PWR_GND_6_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_6_GROM
    );
  PWR_GND_6_YUSED : X_BUF
    port map (
      I => PWR_GND_6_GROM,
      O => GLOBAL_LOGIC0_11
    );
  PWR_GND_7_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_7_GROM
    );
  PWR_GND_7_YUSED : X_BUF
    port map (
      I => PWR_GND_7_GROM,
      O => GLOBAL_LOGIC0_12
    );
  PWR_GND_8_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_8_GROM
    );
  PWR_GND_8_YUSED : X_BUF
    port map (
      I => PWR_GND_8_GROM,
      O => GLOBAL_LOGIC0_13
    );
  PWR_GND_9_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_9_GROM
    );
  PWR_GND_9_YUSED : X_BUF
    port map (
      I => PWR_GND_9_GROM,
      O => GLOBAL_LOGIC0_14
    );
  PWR_GND_10_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_10_GROM
    );
  PWR_GND_10_YUSED : X_BUF
    port map (
      I => PWR_GND_10_GROM,
      O => GLOBAL_LOGIC0_19
    );
  PWR_GND_11_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_11_GROM
    );
  PWR_GND_11_YUSED : X_BUF
    port map (
      I => PWR_GND_11_GROM,
      O => GLOBAL_LOGIC0_22
    );
  PWR_GND_12_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_12_GROM
    );
  PWR_GND_12_YUSED : X_BUF
    port map (
      I => PWR_GND_12_GROM,
      O => GLOBAL_LOGIC0_24
    );
  PWR_GND_13_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_13_GROM
    );
  PWR_GND_13_YUSED : X_BUF
    port map (
      I => PWR_GND_13_GROM,
      O => GLOBAL_LOGIC0_28
    );
  PWR_GND_14_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_14_GROM
    );
  PWR_GND_14_YUSED : X_BUF
    port map (
      I => PWR_GND_14_GROM,
      O => GLOBAL_LOGIC0_29
    );
  PWR_GND_15_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_15_GROM
    );
  PWR_GND_15_YUSED : X_BUF
    port map (
      I => PWR_GND_15_GROM,
      O => GLOBAL_LOGIC0_30
    );
  PWR_GND_16_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_16_GROM
    );
  PWR_GND_16_YUSED : X_BUF
    port map (
      I => PWR_GND_16_GROM,
      O => GLOBAL_LOGIC0_32
    );
  PWR_GND_17_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_17_GROM
    );
  PWR_GND_17_YUSED : X_BUF
    port map (
      I => PWR_GND_17_GROM,
      O => GLOBAL_LOGIC0_34
    );
  PWR_GND_18_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_18_GROM
    );
  PWR_GND_18_YUSED : X_BUF
    port map (
      I => PWR_GND_18_GROM,
      O => GLOBAL_LOGIC0_35
    );
  PWR_GND_19_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_19_GROM
    );
  PWR_GND_19_YUSED : X_BUF
    port map (
      I => PWR_GND_19_GROM,
      O => GLOBAL_LOGIC0_37
    );
  PWR_GND_20_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_20_GROM
    );
  PWR_GND_20_YUSED : X_BUF
    port map (
      I => PWR_GND_20_GROM,
      O => GLOBAL_LOGIC0_38
    );
  PWR_GND_21_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_21_GROM
    );
  PWR_GND_21_YUSED : X_BUF
    port map (
      I => PWR_GND_21_GROM,
      O => GLOBAL_LOGIC0_48
    );
  PWR_GND_22_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_22_GROM
    );
  PWR_GND_22_YUSED : X_BUF
    port map (
      I => PWR_GND_22_GROM,
      O => GLOBAL_LOGIC0_49
    );
  PWR_GND_23_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_23_GROM
    );
  PWR_GND_23_YUSED : X_BUF
    port map (
      I => PWR_GND_23_GROM,
      O => GLOBAL_LOGIC0_50
    );
  PWR_GND_24_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_24_GROM
    );
  PWR_GND_24_YUSED : X_BUF
    port map (
      I => PWR_GND_24_GROM,
      O => GLOBAL_LOGIC0_51
    );
  PWR_GND_25_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_25_GROM
    );
  PWR_GND_25_YUSED : X_BUF
    port map (
      I => PWR_GND_25_GROM,
      O => GLOBAL_LOGIC0_52
    );
  PWR_GND_26_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_26_GROM
    );
  PWR_GND_26_YUSED : X_BUF
    port map (
      I => PWR_GND_26_GROM,
      O => GLOBAL_LOGIC0_53
    );
  PWR_GND_27_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_27_GROM
    );
  PWR_GND_27_YUSED : X_BUF
    port map (
      I => PWR_GND_27_GROM,
      O => GLOBAL_LOGIC0_54
    );
  PWR_GND_28_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_28_GROM
    );
  PWR_GND_28_YUSED : X_BUF
    port map (
      I => PWR_GND_28_GROM,
      O => GLOBAL_LOGIC0_55
    );
  NlwBlock_network_VCC : X_ONE
    port map (
      O => VCC
    );
  NlwBlock_network_GND : X_ZERO
    port map (
      O => GND
    );
  NlwBlockROC : X_ROC
    generic map (ROC_WIDTH => 100 ns)
    port map (O => GSR);
  NlwBlockTOC : X_TOC
    port map (O => GTS);

end Structure;

