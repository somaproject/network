library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
library UNISIM;
use UNISIM.VComponents.all;

entity rambuffer is
    Port ( CLK : in std_logic;
	 		  RESET : in std_logic; 
           DIN : in std_logic_vector(15 downto 0);
           DOUT : out std_logic_vector(15 downto 0);
           WE : in std_logic;
           ADDR : in std_logic_vector(10 downto 0));
end rambuffer;

architecture Behavioral of rambuffer is
-- RAMBUFFER.VHD -- simple wrapper around BlockSelect+ RAMs to make a 1536x16 ram. 

	signal raddr : std_logic_vector(7 downto 0) := (others => '0');
	signal we0, we1, we2, we3, we4, we5 : std_logic := '0';
	signal dout0, dout1, dout2, dout3, dout4, dout5 : 
			std_logic_vector(15 downto 0) := (others => '0');


	component RAMB4_S16
	  generic (
	       INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
	       INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000");

	  port (DI     : in STD_LOGIC_VECTOR (15 downto 0);
	        EN     : in STD_logic;
	        WE     : in STD_logic;
	        RST    : in STD_logic;
	        CLK    : in STD_logic;
	        ADDR   : in STD_LOGIC_VECTOR (7 downto 0);
	        DO     : out STD_LOGIC_VECTOR (15 downto 0)); 
	end component;

	

begin
	raddr <= ADDR(7 downto 0); 
	we0 <= '1' when WE = '1' and ADDR(9 downto 7) = "000" else '0';
	we1 <= '1' when WE = '1' and ADDR(9 downto 7) = "001" else '0';
	we2 <= '1' when WE = '1' and ADDR(9 downto 7) = "010" else '0';
	we3 <= '1' when WE = '1' and ADDR(9 downto 7) = "011" else '0';
	we4 <= '1' when WE = '1' and ADDR(9 downto 7) = "100" else '0';
	we5 <= '1' when WE = '1' and ADDR(9 downto 7) = "101" else '0';

	DOUT <= dout0 when ADDR(9 downto 7) = "000" else
			  dout1 when ADDR(9 downto 7) = "001" else
			  dout2 when ADDR(9 downto 7) = "010" else
			  dout3 when ADDR(9 downto 7) = "011" else
			  dout4 when ADDR(9 downto 7) = "100" else
			  dout5;

	ram0 : RAMB4_S16 generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
				port map (
				DI => DIN,
				EN => '1',
				WE => we0,
				RST => RESET,
				CLK => CLK,
				ADDR => raddr,
				DO => dout0); 

	ram1 : RAMB4_S16 generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
				port map (
				DI => DIN,
				EN => '1',
				WE => we1,
				RST => RESET,
				CLK => CLK,
				ADDR => raddr,
				DO => dout1); 

	ram2 : RAMB4_S16 generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
				port map (
				DI => DIN,
				EN => '1',
				WE => we2,
				RST => RESET,
				CLK => CLK,
				ADDR => raddr,
				DO => dout2); 

	ram3 : RAMB4_S16 generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
				port map (
				DI => DIN,
				EN => '1',
				WE => we3,
				RST => RESET,
				CLK => CLK,
				ADDR => raddr,
				DO => dout3); 

	ram4 : RAMB4_S16 generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
				port map (
				DI => DIN,
				EN => '1',
				WE => we4,
				RST => RESET,
				CLK => CLK,
				ADDR => raddr,
				DO => dout4); 

	ram5 : RAMB4_S16 generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
				port map (
				DI => DIN,
				EN => '1',
				WE => we5,
				RST => RESET,
				CLK => CLK,
				ADDR => raddr,
				DO => dout5); 

				
				 




end Behavioral;
