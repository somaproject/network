-- Xilinx Vhdl netlist produced by netgen application (version G.25a)
-- Command       : -intstyle ise -s 6 -pcf testsuite.pcf -ngm testsuite.ngm -fn -rpw 100 -tpw 0 -ar Structure -xon false -w -ofmt vhdl -sim testsuite.ncd network_PR.vhd 
-- Input file    : testsuite.ncd
-- Output file   : network_PR.vhd
-- Design name   : testsuite
-- # of Entities : 1
-- Xilinx        : C:/Xilinx
-- Device        : 2s200epq208-6 (PRODUCTION 1.17 2003-09-30)

-- This vhdl netlist is a simulation model and uses simulation 
-- primitives which may not represent the true implementation of the 
-- device, however the netlist is functionally correct and should not 
-- be modified. This file cannot be synthesized and should only be used 
-- with supported simulation tools.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library SIMPRIM;
use SIMPRIM.VCOMPONENTS.ALL;
use SIMPRIM.VPACKAGE.ALL;

entity testsuite is
  port (
    DOUTEN : out STD_LOGIC; 
    MCLK : out STD_LOGIC; 
    LED100 : out STD_LOGIC; 
    TESTOUT : out STD_LOGIC; 
    LED1000 : out STD_LOGIC; 
    PHYRESET : out STD_LOGIC; 
    GTX_CLK : out STD_LOGIC; 
    LEDACT : out STD_LOGIC; 
    SOUT : out STD_LOGIC; 
    MWE : out STD_LOGIC; 
    TX_ER : out STD_LOGIC; 
    TX_EN : out STD_LOGIC; 
    LEDDPX : out STD_LOGIC; 
    MOE : out STD_LOGIC; 
    LEDTX : out STD_LOGIC; 
    LEDRX : out STD_LOGIC; 
    LEDPOWER : out STD_LOGIC; 
    MDC : out STD_LOGIC; 
    MDIO : inout STD_LOGIC; 
    SCS : in STD_LOGIC := 'X'; 
    NEXTFRAME : in STD_LOGIC := 'X'; 
    SCLK : in STD_LOGIC := 'X'; 
    DINEN : in STD_LOGIC := 'X'; 
    IFCLK : in STD_LOGIC := 'X'; 
    CLKIOIN : in STD_LOGIC := 'X'; 
    RX_CLK : in STD_LOGIC := 'X'; 
    NEWFRAME : in STD_LOGIC := 'X'; 
    NEXTF : in STD_LOGIC := 'X'; 
    RESET : in STD_LOGIC := 'X'; 
    CLKIN : in STD_LOGIC := 'X'; 
    CLKFB : in STD_LOGIC := 'X'; 
    RX_ER : in STD_LOGIC := 'X'; 
    RX_DV : in STD_LOGIC := 'X'; 
    SIN : in STD_LOGIC := 'X'; 
    DOUT : out STD_LOGIC_VECTOR ( 15 downto 0 ); 
    TXD : out STD_LOGIC_VECTOR ( 7 downto 0 ); 
    MA : out STD_LOGIC_VECTOR ( 16 downto 0 ); 
    MACDATA : out STD_LOGIC_VECTOR ( 15 downto 0 ); 
    MD : inout STD_LOGIC_VECTOR ( 31 downto 0 ); 
    MACADDR : in STD_LOGIC_VECTOR ( 7 downto 0 ); 
    RXD : in STD_LOGIC_VECTOR ( 7 downto 0 ); 
    DIN : in STD_LOGIC_VECTOR ( 15 downto 0 ) 
  );
end testsuite;

architecture Structure of testsuite is
  signal clk : STD_LOGIC; 
  signal maccontrol_N30273 : STD_LOGIC; 
  signal maccontrol_sclkl : STD_LOGIC; 
  signal memtest2_n0119 : STD_LOGIC; 
  signal memtest2_n0030 : STD_LOGIC; 
  signal ifclk_int : STD_LOGIC; 
  signal MCLK_OBUF : STD_LOGIC; 
  signal RESET_IBUF : STD_LOGIC; 
  signal memcontroller_oel : STD_LOGIC; 
  signal txsim_Mshreg_TX_EN_net129 : STD_LOGIC; 
  signal err : STD_LOGIC; 
  signal Q_n0034 : STD_LOGIC; 
  signal CLKFB_IBUFG : STD_LOGIC; 
  signal CLKIN_IBUFG : STD_LOGIC; 
  signal IFCLK_IBUFG : STD_LOGIC; 
  signal rx_clk_int : STD_LOGIC; 
  signal LEDRX_N1683 : STD_LOGIC; 
  signal RX_CLK_IBUFG : STD_LOGIC; 
  signal maccontrol_n0040 : STD_LOGIC; 
  signal maccontrol_n0041 : STD_LOGIC; 
  signal maccontrol_n0043 : STD_LOGIC; 
  signal testrx_nextfl : STD_LOGIC; 
  signal NEXTF_IBUF : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0011 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_sout : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_sts : STD_LOGIC; 
  signal MDC_OBUF : STD_LOGIC; 
  signal memcontroller_n0116 : STD_LOGIC; 
  signal SCS_IBUF : STD_LOGIC; 
  signal SIN_IBUF : STD_LOGIC; 
  signal maccontrol_n0042 : STD_LOGIC; 
  signal RX_ER_IBUF : STD_LOGIC; 
  signal testrx_rx_dvl : STD_LOGIC; 
  signal RX_DV_IBUF : STD_LOGIC; 
  signal GTX_CLK_OBUF : STD_LOGIC; 
  signal maccontrol_n0045 : STD_LOGIC; 
  signal ifclk_to_bufg : STD_LOGIC; 
  signal rx_clk_to_bufg : STD_LOGIC; 
  signal clk_to_bufg : STD_LOGIC; 
  signal testrx_cs_FFd2 : STD_LOGIC; 
  signal GLOBAL_LOGIC0 : STD_LOGIC; 
  signal memcontroller_clknum_0_2 : STD_LOGIC; 
  signal memcontroller_clknum_1_2 : STD_LOGIC; 
  signal maccontrol_PHY_status_miirw : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE826 : STD_LOGIC; 
  signal maccontrol_n0044 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_225 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_123 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_124 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_227 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_125 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_126 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_229 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_127 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_128 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_231 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_129 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_130 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_233 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_131 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_132 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_133 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_134 : STD_LOGIC; 
  signal maccontrol_n0022 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_cy_184 : STD_LOGIC; 
  signal GLOBAL_LOGIC1 : STD_LOGIC; 
  signal maccontrol_Mshreg_scslll_84 : STD_LOGIC; 
  signal maccontrol_bitcnt_85 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_cy_186 : STD_LOGIC; 
  signal maccontrol_bitcnt_86 : STD_LOGIC; 
  signal maccontrol_bitcnt_87 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_cy_188 : STD_LOGIC; 
  signal maccontrol_bitcnt_88 : STD_LOGIC; 
  signal maccontrol_bitcnt_89 : STD_LOGIC; 
  signal maccontrol_bitcnt_90 : STD_LOGIC; 
  signal maccontrol_N30218 : STD_LOGIC; 
  signal maccontrol_sclkdeltall : STD_LOGIC; 
  signal maccontrol_n00541_1 : STD_LOGIC; 
  signal maccontrol_n0039124_1 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_191 : STD_LOGIC; 
  signal maccontrol_N30228 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1231_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_91 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_193 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_92 : STD_LOGIC; 
  signal maccontrol_N30199 : STD_LOGIC; 
  signal maccontrol_N46337 : STD_LOGIC; 
  signal maccontrol_Ker303141_1 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_93 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_195 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_94 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_95 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_197 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_96 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_97 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_199 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_98 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_99 : STD_LOGIC; 
  signal maccontrol_n0039 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_201 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_100 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_101 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_203 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_102 : STD_LOGIC; 
  signal maccontrol_Ker303141_2 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_103 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_205 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_104 : STD_LOGIC; 
  signal maccontrol_N30285 : STD_LOGIC; 
  signal maccontrol_N46356 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_105 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_207 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_106 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_107 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_209 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_108 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_109 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_211 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_110 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_111 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_213 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_112 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_113 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_215 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_114 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_115 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_217 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_116 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_117 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_219 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_118 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_119 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_221 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_120 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_121 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_122 : STD_LOGIC; 
  signal maccontrol_CHOICE1608 : STD_LOGIC; 
  signal clkslen : STD_LOGIC; 
  signal cnt0_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal cnt0_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal memtest2_Mcompar_n0020_inst_cy_167 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_24_45 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_25_44 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_26_43 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_27_42 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_28_41 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_29_40 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_30_39 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_31_38 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_1 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_3 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_5 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_7 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_9 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_11 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_13 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_15 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0013 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_122 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd5 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_124 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_126 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N41734 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_129 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_0_37 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_1_36 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_2_35 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_3_34 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_131 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_4_33 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_5_32 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_6_31 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_7_30 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_133 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_8_29 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_9_28 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_10_27 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_11_26 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_135 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_12_25 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_13_24 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_14_23 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_15_22 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_137 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_16_21 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_17_20 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_18_19 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_19_18 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_139 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_20_17 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_21_16 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_22_15 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_23_14 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_141 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_24_13 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_25_12 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_26_11 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_27_10 : STD_LOGIC; 
  signal memtest_n0002 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_28_9 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_29_8 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_30_7 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_31_6 : STD_LOGIC; 
  signal testrx_addr_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal testrx_n0008 : STD_LOGIC; 
  signal testrx_addr_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal testrx_addr_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal memcontroller_Ker256691_O : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_87 : STD_LOGIC; 
  signal memtest2_n0011 : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_89 : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_91 : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_93 : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_95 : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_97 : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_99 : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_101 : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_161 : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_163 : STD_LOGIC; 
  signal memtest2_n0025 : STD_LOGIC; 
  signal memtest2_Mcompar_n0017_inst_cy_167 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_0_69 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_1_68 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_2_67 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_3_66 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_4_65 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_5_64 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_6_63 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_7_62 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_25 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_27 : STD_LOGIC; 
  signal memtest2_Mcompar_n0018_inst_cy_167 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_8_61 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_9_60 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_10_59 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_11_58 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_12_57 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_13_56 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_14_55 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_15_54 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_153 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_155 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_157 : STD_LOGIC; 
  signal memtest2_n0027 : STD_LOGIC; 
  signal memtest2_Mcompar_n0019_inst_cy_167 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_16_53 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_17_52 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_18_51 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_19_50 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_20_49 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_21_48 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_22_47 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_23_46 : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_104 : STD_LOGIC; 
  signal txsim_SF22758 : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_106 : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_108 : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_110 : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_112 : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_114 : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_116 : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_118 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_145 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_147 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_149 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut4_16 : STD_LOGIC; 
  signal memtest2_n0028 : STD_LOGIC; 
  signal clken1 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_47 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_49 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_51 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_53 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_55 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_57 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_59 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_61 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_63 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_65 : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_67 : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_71 : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_73 : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_75 : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_77 : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_79 : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_81 : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_83 : STD_LOGIC; 
  signal memtest2_n00511_1 : STD_LOGIC; 
  signal memtest2_n00511_O : STD_LOGIC; 
  signal memtest2_n00511_4 : STD_LOGIC; 
  signal maccontrol_n0012 : STD_LOGIC; 
  signal maccontrol_CHOICE1446 : STD_LOGIC; 
  signal maccontrol_CHOICE1443 : STD_LOGIC; 
  signal maccontrol_CHOICE1439 : STD_LOGIC; 
  signal maccontrol_N30162 : STD_LOGIC; 
  signal maccontrol_N30238 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_0_92_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1426 : STD_LOGIC; 
  signal maccontrol_CHOICE1433 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_14_58_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1055 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_1_58_SW0_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_2_26_2 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_2_26_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1471 : STD_LOGIC; 
  signal maccontrol_CHOICE1474 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_2_58_SW0_O : STD_LOGIC; 
  signal maccontrol_n001223_1 : STD_LOGIC; 
  signal maccontrol_N46555 : STD_LOGIC; 
  signal maccontrol_N46518 : STD_LOGIC; 
  signal maccontrol_CHOICE1269 : STD_LOGIC; 
  signal maccontrol_addr_0_1 : STD_LOGIC; 
  signal maccontrol_addr_1_1 : STD_LOGIC; 
  signal maccontrol_CHOICE1281 : STD_LOGIC; 
  signal maccontrol_CHOICE1266 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_4_32_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_5_26_2 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_5_26_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1507 : STD_LOGIC; 
  signal maccontrol_CHOICE1510 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_5_58_SW0_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_8_58_SW0_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_6_58_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1364 : STD_LOGIC; 
  signal maccontrol_n00691_1 : STD_LOGIC; 
  signal maccontrol_CHOICE1376 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_7_76_SW0_O : STD_LOGIC; 
  signal memtest2_n0116 : STD_LOGIC; 
  signal maccontrol_N46526 : STD_LOGIC; 
  signal maccontrol_CHOICE1288 : STD_LOGIC; 
  signal maccontrol_CHOICE1300 : STD_LOGIC; 
  signal maccontrol_CHOICE1285 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_9_32_O : STD_LOGIC; 
  signal memtest2_n01161_1 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_13_net101 : STD_LOGIC; 
  signal memtest2_n00511_3 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_21_net85 : STD_LOGIC; 
  signal memtest2_n00511_2 : STD_LOGIC; 
  signal maccontrol_N30212 : STD_LOGIC; 
  signal maccontrol_N30192 : STD_LOGIC; 
  signal maccontrol_N30292 : STD_LOGIC; 
  signal maccontrol_n0067 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_13_18_O : STD_LOGIC; 
  signal maccontrol_N46514 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_10_26_2 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_10_26_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1543 : STD_LOGIC; 
  signal maccontrol_CHOICE1546 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_10_58_SW0_O : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd1 : STD_LOGIC; 
  signal maccontrol_PHY_status_n00151_O : STD_LOGIC; 
  signal maccontrol_N46368 : STD_LOGIC; 
  signal maccontrol_N42043 : STD_LOGIC; 
  signal maccontrol_PHY_status_n00151_1 : STD_LOGIC; 
  signal maccontrol_n0069 : STD_LOGIC; 
  signal maccontrol_PHY_status_phyaddrws : STD_LOGIC; 
  signal maccontrol_CHOICE1397 : STD_LOGIC; 
  signal maccontrol_CHOICE1385 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_11_76_SW0_O : STD_LOGIC; 
  signal maccontrol_N46522 : STD_LOGIC; 
  signal maccontrol_CHOICE1307 : STD_LOGIC; 
  signal maccontrol_CHOICE1319 : STD_LOGIC; 
  signal maccontrol_CHOICE1304 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_12_32_O : STD_LOGIC; 
  signal maccontrol_CHOICE1120 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_20_22_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1245 : STD_LOGIC; 
  signal maccontrol_n00671_1 : STD_LOGIC; 
  signal maccontrol_CHOICE1251 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_21_12_O : STD_LOGIC; 
  signal maccontrol_CHOICE1326 : STD_LOGIC; 
  signal maccontrol_CHOICE1338 : STD_LOGIC; 
  signal maccontrol_CHOICE1323 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_13_32_O : STD_LOGIC; 
  signal maccontrol_CHOICE1165 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_30_22_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1129 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_22_22_SW0_O : STD_LOGIC; 
  signal maccontrol_n0068 : STD_LOGIC; 
  signal maccontrol_CHOICE1204 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_23_25_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1184 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_31_25_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1406 : STD_LOGIC; 
  signal maccontrol_CHOICE1418 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_15_76_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1256 : STD_LOGIC; 
  signal maccontrol_CHOICE1262 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_24_12_O : STD_LOGIC; 
  signal maccontrol_CHOICE1223 : STD_LOGIC; 
  signal maccontrol_CHOICE1229 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_16_12_O : STD_LOGIC; 
  signal maccontrol_CHOICE1234 : STD_LOGIC; 
  signal maccontrol_CHOICE1240 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_17_12_O : STD_LOGIC; 
  signal maccontrol_CHOICE1138 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_25_22_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1111 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_18_22_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1147 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_26_22_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1214 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_27_25_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1194 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_19_25_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1156 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_28_22_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1174 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_29_22_SW0_O : STD_LOGIC; 
  signal maccontrol_n0070 : STD_LOGIC; 
  signal maccontrol_n0071 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_6_26_2 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_6_26_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1489 : STD_LOGIC; 
  signal maccontrol_CHOICE1492 : STD_LOGIC; 
  signal maccontrol_n0084 : STD_LOGIC; 
  signal maccontrol_N30305 : STD_LOGIC; 
  signal maccontrol_n0085 : STD_LOGIC; 
  signal maccontrol_n0083 : STD_LOGIC; 
  signal memtest2_Ker2265849_2 : STD_LOGIC; 
  signal memtest2_Ker2265830_O : STD_LOGIC; 
  signal memtest2_N22660 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_9_18_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_14_26_2 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_14_26_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1561 : STD_LOGIC; 
  signal maccontrol_CHOICE1564 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_8_26_2 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_8_26_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1525 : STD_LOGIC; 
  signal maccontrol_CHOICE1528 : STD_LOGIC; 
  signal maccontrol_n00701_1 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_1_26_2 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_1_26_SW0_O : STD_LOGIC; 
  signal maccontrol_CHOICE1453 : STD_LOGIC; 
  signal maccontrol_CHOICE1456 : STD_LOGIC; 
  signal maccontrol_lrxucast : STD_LOGIC; 
  signal maccontrol_CHOICE1429 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_0_11_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O : STD_LOGIC; 
  signal maccontrol_N46462 : STD_LOGIC; 
  signal maccontrol_N30311 : STD_LOGIC; 
  signal maccontrol_sclkdelta : STD_LOGIC; 
  signal maccontrol_N46628 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_4_18_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_3_6_O : STD_LOGIC; 
  signal maccontrol_CHOICE1355 : STD_LOGIC; 
  signal maccontrol_n00397_O : STD_LOGIC; 
  signal maccontrol_CHOICE1582 : STD_LOGIC; 
  signal maccontrol_newcmd : STD_LOGIC; 
  signal maccontrol_N30181 : STD_LOGIC; 
  signal maccontrol_n0034 : STD_LOGIC; 
  signal maccontrol_CHOICE1585 : STD_LOGIC; 
  signal maccontrol_n003923_O : STD_LOGIC; 
  signal maccontrol_CHOICE1589 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_12_18_O : STD_LOGIC; 
  signal maccontrol_N30299 : STD_LOGIC; 
  signal maccontrol_PHY_status_n00171_O : STD_LOGIC; 
  signal maccontrol_PHY_status_n00181_O : STD_LOGIC; 
  signal clken4 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd3 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd4 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0004 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE925 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd6 : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd8 : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd6 : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd3 : STD_LOGIC; 
  signal memcontroller_clknum_1_1 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0010 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0004_2 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0079 : STD_LOGIC; 
  signal memtest2_lfsr_rst : STD_LOGIC; 
  signal clken_n0002 : STD_LOGIC; 
  signal maccontrol_PHY_status_done : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd2 : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd5 : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd4 : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd7 : STD_LOGIC; 
  signal maccontrol_Mshreg_sinlll_83 : STD_LOGIC; 
  signal testrx_cs_FFd3 : STD_LOGIC; 
  signal testrx_n0004 : STD_LOGIC; 
  signal testrx_cs_FFd1 : STD_LOGIC; 
  signal testrx_N41780 : STD_LOGIC; 
  signal maccontrol_sclkll : STD_LOGIC; 
  signal mwe2 : STD_LOGIC; 
  signal memcontroller_oe : STD_LOGIC; 
  signal memtest_lerr : STD_LOGIC; 
  signal maccontrol_PHY_status_n0021 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE784 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE770 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N46672 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N46670 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE793 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N20226 : STD_LOGIC; 
  signal memcontroller_n0005 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd2 : STD_LOGIC; 
  signal maccontrol_PHY_status_n0011 : STD_LOGIC; 
  signal memcontroller_n0007 : STD_LOGIC; 
  signal maccontrol_N46689 : STD_LOGIC; 
  signal maccontrol_CHOICE1368 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_7_40_SW0_O : STD_LOGIC; 
  signal maccontrol_PHY_status_N23512 : STD_LOGIC; 
  signal memtest2_CHOICE1064 : STD_LOGIC; 
  signal memtest2_CHOICE1071 : STD_LOGIC; 
  signal memtest2_CHOICE1067 : STD_LOGIC; 
  signal maccontrol_n0031 : STD_LOGIC; 
  signal maccontrol_n00311_1 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0016 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE920 : STD_LOGIC; 
  signal Q_n0034_2 : STD_LOGIC; 
  signal maccontrol_n0035 : STD_LOGIC; 
  signal maccontrol_n0036 : STD_LOGIC; 
  signal maccontrol_n0037 : STD_LOGIC; 
  signal memcontroller_clknum_0_1 : STD_LOGIC; 
  signal memtest2_CHOICE948 : STD_LOGIC; 
  signal memtest2_CHOICE941 : STD_LOGIC; 
  signal memtest2_n002184_2 : STD_LOGIC; 
  signal memtest2_n002184_SW0_2 : STD_LOGIC; 
  signal testrx_CHOICE930 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE735 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N46530 : STD_LOGIC; 
  signal testrx_CHOICE933 : STD_LOGIC; 
  signal maccontrol_N30206 : STD_LOGIC; 
  signal maccontrol_lrxmcast : STD_LOGIC; 
  signal maccontrol_n0032 : STD_LOGIC; 
  signal maccontrol_lrxbcast : STD_LOGIC; 
  signal maccontrol_lrxallf : STD_LOGIC; 
  signal maccontrol_N46676 : STD_LOGIC; 
  signal maccontrol_N46406 : STD_LOGIC; 
  signal txsim_SF22756 : STD_LOGIC; 
  signal txsim_llltx : STD_LOGIC; 
  signal txsim_N41883 : STD_LOGIC; 
  signal maccontrol_N46681 : STD_LOGIC; 
  signal maccontrol_CHOICE1410 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_15_40_SW0_O : STD_LOGIC; 
  signal memtest_llerr : STD_LOGIC; 
  signal memtest2_n0117 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N20221 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE800 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N41816 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE741 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE749 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE750 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE751 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_sout498_2 : STD_LOGIC; 
  signal maccontrol_n0013 : STD_LOGIC; 
  signal maccontrol_n00131_1 : STD_LOGIC; 
  signal maccontrol_PHY_status_n0019 : STD_LOGIC; 
  signal maccontrol_N46685 : STD_LOGIC; 
  signal maccontrol_CHOICE1347 : STD_LOGIC; 
  signal maccontrol_CHOICE1389 : STD_LOGIC; 
  signal maccontrol_n003963_O : STD_LOGIC; 
  signal maccontrol_CHOICE1603 : STD_LOGIC; 
  signal maccontrol_CHOICE1596 : STD_LOGIC; 
  signal maccontrol_N46402 : STD_LOGIC; 
  signal maccontrol_CHOICE1605 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE831 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE764 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE802 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE812 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE813 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE829 : STD_LOGIC; 
  signal maccontrol_sclkdeltal : STD_LOGIC; 
  signal maccontrol_PHY_status_N23520 : STD_LOGIC; 
  signal maccontrol_PHY_status_n0020 : STD_LOGIC; 
  signal clken_n0005 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE729 : STD_LOGIC; 
  signal maccontrol_n0010 : STD_LOGIC; 
  signal memtest2_N41527 : STD_LOGIC; 
  signal maccontrol_PHY_status_N42089 : STD_LOGIC; 
  signal txsim_CHOICE1098 : STD_LOGIC; 
  signal txsim_CHOICE1105 : STD_LOGIC; 
  signal txsim_N46398 : STD_LOGIC; 
  signal txsim_CHOICE1090 : STD_LOGIC; 
  signal maccontrol_n0011 : STD_LOGIC; 
  signal maccontrol_n0234 : STD_LOGIC; 
  signal maccontrol_PHY_status_start : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_11_40_SW0_O : STD_LOGIC; 
  signal maccontrol_n0033 : STD_LOGIC; 
  signal clken_lclken : STD_LOGIC; 
  signal maccontrol_CHOICE1033 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N46538 : STD_LOGIC; 
  signal maccontrol_CHOICE1041 : STD_LOGIC; 
  signal maccontrol_CHOICE1048 : STD_LOGIC; 
  signal maccontrol_CHOICE1003 : STD_LOGIC; 
  signal maccontrol_CHOICE1018 : STD_LOGIC; 
  signal maccontrol_CHOICE1050 : STD_LOGIC; 
  signal maccontrol_N30316 : STD_LOGIC; 
  signal maccontrol_CHOICE1002 : STD_LOGIC; 
  signal maccontrol_CHOICE1010 : STD_LOGIC; 
  signal maccontrol_PHY_status_rwl : STD_LOGIC; 
  signal maccontrol_CHOICE1017 : STD_LOGIC; 
  signal maccontrol_CHOICE974 : STD_LOGIC; 
  signal maccontrol_CHOICE988 : STD_LOGIC; 
  signal maccontrol_CHOICE981 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_0 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_1 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_2 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_3 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_4 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_5 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_6 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_7 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_8 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_9 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_10 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_11 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_12 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_13 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_14 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_15 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_16 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_17 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_18 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_19 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_20 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_21 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_22 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_23 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_24 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_25 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_26 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_27 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_28 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_29 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_30 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_31 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_32 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_33 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_34 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_35 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_36 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_37 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_38 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_39 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_40 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_41 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_42 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_43 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_44 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_45 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_46 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_0 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_1 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_2 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_3 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_4 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_5 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_6 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_7 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_8 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_9 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_10 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_11 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_12 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_13 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_14 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_15 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_16 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_17 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_18 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_19 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_20 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_21 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_22 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_23 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_24 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_25 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_26 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_27 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_28 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_29 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_30 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_31 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_32 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_33 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_34 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_35 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_36 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_37 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_38 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_39 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_40 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_41 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_42 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_43 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_44 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_45 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_46 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_47 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_48 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_49 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_50 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_51 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_52 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_53 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_54 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_55 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_56 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_57 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_58 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_59 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_60 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_61 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_62 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_63 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_64 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_65 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_66 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_67 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_68 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_69 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_70 : STD_LOGIC; 
  signal GSR : STD_LOGIC; 
  signal GTS : STD_LOGIC; 
  signal SCLK_IFF_RST : STD_LOGIC; 
  signal maccontrol_SCLK_IBUF : STD_LOGIC; 
  signal TESTOUT_OFF_RST : STD_LOGIC; 
  signal TESTOUT_ENABLE : STD_LOGIC; 
  signal TESTOUT_TORGTS : STD_LOGIC; 
  signal TESTOUT_OUTMUX : STD_LOGIC; 
  signal memtest2_ERR : STD_LOGIC; 
  signal TESTOUT_OD : STD_LOGIC; 
  signal TXD_0_OFF_RST : STD_LOGIC; 
  signal TXD_0_ENABLE : STD_LOGIC; 
  signal TXD_0_TORGTS : STD_LOGIC; 
  signal TXD_0_OUTMUX : STD_LOGIC; 
  signal txsim_TXD_0_OBUF : STD_LOGIC; 
  signal TXD_0_OD : STD_LOGIC; 
  signal TXD_1_OFF_RST : STD_LOGIC; 
  signal TXD_1_ENABLE : STD_LOGIC; 
  signal TXD_1_TORGTS : STD_LOGIC; 
  signal TXD_1_OUTMUX : STD_LOGIC; 
  signal txsim_TXD_1_OBUF : STD_LOGIC; 
  signal TXD_1_OD : STD_LOGIC; 
  signal TXD_2_OFF_RST : STD_LOGIC; 
  signal TXD_2_ENABLE : STD_LOGIC; 
  signal TXD_2_TORGTS : STD_LOGIC; 
  signal TXD_2_OUTMUX : STD_LOGIC; 
  signal txsim_TXD_2_OBUF : STD_LOGIC; 
  signal TXD_2_OD : STD_LOGIC; 
  signal TXD_3_OFF_RST : STD_LOGIC; 
  signal TXD_3_ENABLE : STD_LOGIC; 
  signal TXD_3_TORGTS : STD_LOGIC; 
  signal TXD_3_OUTMUX : STD_LOGIC; 
  signal txsim_TXD_3_OBUF : STD_LOGIC; 
  signal TXD_3_OD : STD_LOGIC; 
  signal TXD_4_OFF_RST : STD_LOGIC; 
  signal TXD_4_ENABLE : STD_LOGIC; 
  signal TXD_4_TORGTS : STD_LOGIC; 
  signal TXD_4_OUTMUX : STD_LOGIC; 
  signal txsim_TXD_4_OBUF : STD_LOGIC; 
  signal TXD_4_OD : STD_LOGIC; 
  signal TXD_5_OFF_RST : STD_LOGIC; 
  signal TXD_5_ENABLE : STD_LOGIC; 
  signal TXD_5_TORGTS : STD_LOGIC; 
  signal TXD_5_OUTMUX : STD_LOGIC; 
  signal txsim_TXD_5_OBUF : STD_LOGIC; 
  signal TXD_5_OD : STD_LOGIC; 
  signal TXD_6_OFF_RST : STD_LOGIC; 
  signal TXD_6_ENABLE : STD_LOGIC; 
  signal TXD_6_TORGTS : STD_LOGIC; 
  signal TXD_6_OUTMUX : STD_LOGIC; 
  signal txsim_TXD_6_OBUF : STD_LOGIC; 
  signal TXD_6_OD : STD_LOGIC; 
  signal TXD_7_ENABLE : STD_LOGIC; 
  signal TXD_7_TORGTS : STD_LOGIC; 
  signal TXD_7_OUTMUX : STD_LOGIC; 
  signal txsim_TXD_7_OBUF : STD_LOGIC; 
  signal TXD_7_OD : STD_LOGIC; 
  signal testrx_MACADDR_0_IBUF : STD_LOGIC; 
  signal testrx_MACADDR_1_IBUF : STD_LOGIC; 
  signal testrx_MACADDR_2_IBUF : STD_LOGIC; 
  signal testrx_MACADDR_3_IBUF : STD_LOGIC; 
  signal testrx_MACADDR_4_IBUF : STD_LOGIC; 
  signal testrx_MACADDR_5_IBUF : STD_LOGIC; 
  signal testrx_MACADDR_6_IBUF : STD_LOGIC; 
  signal testrx_MACADDR_7_IBUF : STD_LOGIC; 
  signal MCLK_ENABLE : STD_LOGIC; 
  signal MCLK_TORGTS : STD_LOGIC; 
  signal MCLK_OUTMUX : STD_LOGIC; 
  signal MA_0_ENABLE : STD_LOGIC; 
  signal MA_0_TORGTS : STD_LOGIC; 
  signal MA_0_OUTMUX : STD_LOGIC; 
  signal MA_0_OCEMUXNOT : STD_LOGIC; 
  signal MA_0_OD : STD_LOGIC; 
  signal MA_1_ENABLE : STD_LOGIC; 
  signal MA_1_TORGTS : STD_LOGIC; 
  signal MA_1_OUTMUX : STD_LOGIC; 
  signal MA_1_OCEMUXNOT : STD_LOGIC; 
  signal MA_1_OD : STD_LOGIC; 
  signal MA_2_ENABLE : STD_LOGIC; 
  signal MA_2_TORGTS : STD_LOGIC; 
  signal MA_2_OUTMUX : STD_LOGIC; 
  signal MA_2_OCEMUXNOT : STD_LOGIC; 
  signal MA_2_OD : STD_LOGIC; 
  signal MA_3_ENABLE : STD_LOGIC; 
  signal MA_3_TORGTS : STD_LOGIC; 
  signal MA_3_OUTMUX : STD_LOGIC; 
  signal MA_3_OCEMUXNOT : STD_LOGIC; 
  signal MA_3_OD : STD_LOGIC; 
  signal MA_4_ENABLE : STD_LOGIC; 
  signal MA_4_TORGTS : STD_LOGIC; 
  signal MA_4_OUTMUX : STD_LOGIC; 
  signal MA_4_OCEMUXNOT : STD_LOGIC; 
  signal MA_4_OD : STD_LOGIC; 
  signal TXD_7_OFF_RST : STD_LOGIC; 
  signal MA_5_ENABLE : STD_LOGIC; 
  signal MA_5_TORGTS : STD_LOGIC; 
  signal MA_5_OUTMUX : STD_LOGIC; 
  signal MA_5_OCEMUXNOT : STD_LOGIC; 
  signal MA_5_OD : STD_LOGIC; 
  signal MA_6_ENABLE : STD_LOGIC; 
  signal MA_6_TORGTS : STD_LOGIC; 
  signal MA_6_OUTMUX : STD_LOGIC; 
  signal MA_6_OCEMUXNOT : STD_LOGIC; 
  signal MA_6_OD : STD_LOGIC; 
  signal MA_7_ENABLE : STD_LOGIC; 
  signal MA_7_TORGTS : STD_LOGIC; 
  signal MA_7_OUTMUX : STD_LOGIC; 
  signal MA_7_OCEMUXNOT : STD_LOGIC; 
  signal MA_7_OD : STD_LOGIC; 
  signal MA_8_ENABLE : STD_LOGIC; 
  signal MA_8_TORGTS : STD_LOGIC; 
  signal MA_8_OUTMUX : STD_LOGIC; 
  signal MA_8_OCEMUXNOT : STD_LOGIC; 
  signal MA_8_OD : STD_LOGIC; 
  signal MA_9_ENABLE : STD_LOGIC; 
  signal MA_9_TORGTS : STD_LOGIC; 
  signal MA_9_OUTMUX : STD_LOGIC; 
  signal MA_9_OCEMUXNOT : STD_LOGIC; 
  signal MA_9_OD : STD_LOGIC; 
  signal MD_0_ENABLE : STD_LOGIC; 
  signal MD_0_TORGTS : STD_LOGIC; 
  signal MD_0_OUTMUX : STD_LOGIC; 
  signal MD_0_OD : STD_LOGIC; 
  signal MD_1_ENABLE : STD_LOGIC; 
  signal MD_1_TORGTS : STD_LOGIC; 
  signal MD_1_OUTMUX : STD_LOGIC; 
  signal MD_1_OD : STD_LOGIC; 
  signal TX_EN_ENABLE : STD_LOGIC; 
  signal TX_EN_TORGTS : STD_LOGIC; 
  signal TX_EN_OUTMUX : STD_LOGIC; 
  signal txsim_TX_EN_OBUF : STD_LOGIC; 
  signal TX_EN_OD : STD_LOGIC; 
  signal MD_2_ENABLE : STD_LOGIC; 
  signal MD_2_TORGTS : STD_LOGIC; 
  signal MD_2_OUTMUX : STD_LOGIC; 
  signal MD_2_OD : STD_LOGIC; 
  signal MD_3_ENABLE : STD_LOGIC; 
  signal MD_3_TORGTS : STD_LOGIC; 
  signal MD_3_OUTMUX : STD_LOGIC; 
  signal MD_3_OD : STD_LOGIC; 
  signal MD_4_ENABLE : STD_LOGIC; 
  signal MD_4_TORGTS : STD_LOGIC; 
  signal MD_4_OUTMUX : STD_LOGIC; 
  signal MD_4_OD : STD_LOGIC; 
  signal MD_5_ENABLE : STD_LOGIC; 
  signal MD_5_TORGTS : STD_LOGIC; 
  signal MD_5_OUTMUX : STD_LOGIC; 
  signal MD_5_OD : STD_LOGIC; 
  signal MD_6_ENABLE : STD_LOGIC; 
  signal MD_6_TORGTS : STD_LOGIC; 
  signal MD_6_OUTMUX : STD_LOGIC; 
  signal MD_6_OD : STD_LOGIC; 
  signal MD_7_ENABLE : STD_LOGIC; 
  signal MD_7_TORGTS : STD_LOGIC; 
  signal MD_7_OUTMUX : STD_LOGIC; 
  signal MD_7_OD : STD_LOGIC; 
  signal MD_8_ENABLE : STD_LOGIC; 
  signal MD_8_TORGTS : STD_LOGIC; 
  signal MD_8_OUTMUX : STD_LOGIC; 
  signal MD_8_OD : STD_LOGIC; 
  signal MD_9_ENABLE : STD_LOGIC; 
  signal MD_9_TORGTS : STD_LOGIC; 
  signal MD_9_OUTMUX : STD_LOGIC; 
  signal MD_9_OD : STD_LOGIC; 
  signal LEDACT_ENABLE : STD_LOGIC; 
  signal LEDACT_TORGTS : STD_LOGIC; 
  signal LEDACT_OUTMUX : STD_LOGIC; 
  signal LEDACT_OBUF : STD_LOGIC; 
  signal LEDACT_OCEMUXNOT : STD_LOGIC; 
  signal LEDACT_OD : STD_LOGIC; 
  signal MACADDR_0_IFF_RST : STD_LOGIC; 
  signal LEDDPX_ENABLE : STD_LOGIC; 
  signal LEDDPX_TORGTS : STD_LOGIC; 
  signal LEDDPX_OUTMUX : STD_LOGIC; 
  signal maccontrol_LEDDPX_OBUF : STD_LOGIC; 
  signal LEDDPX_OD : STD_LOGIC; 
  signal LEDRX_ENABLE : STD_LOGIC; 
  signal LEDRX_TORGTS : STD_LOGIC; 
  signal LEDRX_OUTMUX : STD_LOGIC; 
  signal LEDRX_OBUF : STD_LOGIC; 
  signal LEDRX_LOGIC_ONE : STD_LOGIC; 
  signal MA_10_ENABLE : STD_LOGIC; 
  signal MA_10_TORGTS : STD_LOGIC; 
  signal MA_10_OUTMUX : STD_LOGIC; 
  signal MA_10_OCEMUXNOT : STD_LOGIC; 
  signal MA_10_OD : STD_LOGIC; 
  signal MA_11_ENABLE : STD_LOGIC; 
  signal MA_11_TORGTS : STD_LOGIC; 
  signal MA_11_OUTMUX : STD_LOGIC; 
  signal MA_11_OCEMUXNOT : STD_LOGIC; 
  signal MA_11_OD : STD_LOGIC; 
  signal MA_12_ENABLE : STD_LOGIC; 
  signal MA_12_TORGTS : STD_LOGIC; 
  signal MA_12_OUTMUX : STD_LOGIC; 
  signal MA_12_OCEMUXNOT : STD_LOGIC; 
  signal MA_12_OD : STD_LOGIC; 
  signal MA_13_ENABLE : STD_LOGIC; 
  signal MA_13_TORGTS : STD_LOGIC; 
  signal MA_13_OUTMUX : STD_LOGIC; 
  signal MA_13_OCEMUXNOT : STD_LOGIC; 
  signal MA_13_OD : STD_LOGIC; 
  signal MA_14_ENABLE : STD_LOGIC; 
  signal MA_14_TORGTS : STD_LOGIC; 
  signal MA_14_OUTMUX : STD_LOGIC; 
  signal MA_14_OCEMUXNOT : STD_LOGIC; 
  signal MA_14_OD : STD_LOGIC; 
  signal MA_15_ENABLE : STD_LOGIC; 
  signal MA_15_TORGTS : STD_LOGIC; 
  signal MA_15_OUTMUX : STD_LOGIC; 
  signal MA_15_OCEMUXNOT : STD_LOGIC; 
  signal MA_15_OD : STD_LOGIC; 
  signal MA_16_ENABLE : STD_LOGIC; 
  signal MA_16_TORGTS : STD_LOGIC; 
  signal MA_16_OUTMUX : STD_LOGIC; 
  signal MA_16_OCEMUXNOT : STD_LOGIC; 
  signal MA_16_OD : STD_LOGIC; 
  signal SOUT_ENABLE : STD_LOGIC; 
  signal SOUT_TORGTS : STD_LOGIC; 
  signal SOUT_OUTMUX : STD_LOGIC; 
  signal maccontrol_SOUT_OBUF : STD_LOGIC; 
  signal SOUT_OD : STD_LOGIC; 
  signal MACDATA_0_ENABLE : STD_LOGIC; 
  signal MACDATA_0_TORGTS : STD_LOGIC; 
  signal MACDATA_0_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_0_OBUF : STD_LOGIC; 
  signal MACDATA_0_OD : STD_LOGIC; 
  signal MACADDR_1_IFF_RST : STD_LOGIC; 
  signal MACDATA_1_ENABLE : STD_LOGIC; 
  signal MACDATA_1_TORGTS : STD_LOGIC; 
  signal MACDATA_1_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_1_OBUF : STD_LOGIC; 
  signal MACDATA_1_OD : STD_LOGIC; 
  signal MACDATA_2_ENABLE : STD_LOGIC; 
  signal MACDATA_2_TORGTS : STD_LOGIC; 
  signal MACDATA_2_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_2_OBUF : STD_LOGIC; 
  signal MACDATA_2_OD : STD_LOGIC; 
  signal MACDATA_3_ENABLE : STD_LOGIC; 
  signal MACDATA_3_TORGTS : STD_LOGIC; 
  signal MACDATA_3_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_3_OBUF : STD_LOGIC; 
  signal MACDATA_3_OD : STD_LOGIC; 
  signal MACDATA_4_ENABLE : STD_LOGIC; 
  signal MACDATA_4_TORGTS : STD_LOGIC; 
  signal MACDATA_4_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_4_OBUF : STD_LOGIC; 
  signal MACDATA_4_OD : STD_LOGIC; 
  signal MACDATA_5_ENABLE : STD_LOGIC; 
  signal MACDATA_5_TORGTS : STD_LOGIC; 
  signal MACDATA_5_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_5_OBUF : STD_LOGIC; 
  signal MACDATA_5_OD : STD_LOGIC; 
  signal MACDATA_6_ENABLE : STD_LOGIC; 
  signal MACDATA_6_TORGTS : STD_LOGIC; 
  signal MACDATA_6_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_6_OBUF : STD_LOGIC; 
  signal MACDATA_6_OD : STD_LOGIC; 
  signal MACDATA_7_ENABLE : STD_LOGIC; 
  signal MACDATA_7_TORGTS : STD_LOGIC; 
  signal MACDATA_7_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_7_OBUF : STD_LOGIC; 
  signal MACDATA_7_OD : STD_LOGIC; 
  signal MACDATA_8_ENABLE : STD_LOGIC; 
  signal MACDATA_8_TORGTS : STD_LOGIC; 
  signal MACDATA_8_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_8_OBUF : STD_LOGIC; 
  signal MACDATA_8_OD : STD_LOGIC; 
  signal MD_10_ENABLE : STD_LOGIC; 
  signal MD_10_TORGTS : STD_LOGIC; 
  signal MD_10_OUTMUX : STD_LOGIC; 
  signal MD_10_OD : STD_LOGIC; 
  signal MACADDR_2_IFF_RST : STD_LOGIC; 
  signal MACDATA_9_ENABLE : STD_LOGIC; 
  signal MACDATA_9_TORGTS : STD_LOGIC; 
  signal MACDATA_9_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_9_OBUF : STD_LOGIC; 
  signal MACDATA_9_OD : STD_LOGIC; 
  signal MD_11_ENABLE : STD_LOGIC; 
  signal MD_11_TORGTS : STD_LOGIC; 
  signal MD_11_OUTMUX : STD_LOGIC; 
  signal MD_11_OD : STD_LOGIC; 
  signal MD_20_ENABLE : STD_LOGIC; 
  signal MD_20_TORGTS : STD_LOGIC; 
  signal MD_20_OUTMUX : STD_LOGIC; 
  signal MD_20_OD : STD_LOGIC; 
  signal MD_12_ENABLE : STD_LOGIC; 
  signal MD_12_TORGTS : STD_LOGIC; 
  signal MD_12_OUTMUX : STD_LOGIC; 
  signal MD_12_OD : STD_LOGIC; 
  signal MD_21_ENABLE : STD_LOGIC; 
  signal MD_21_TORGTS : STD_LOGIC; 
  signal MD_21_OUTMUX : STD_LOGIC; 
  signal MD_21_OD : STD_LOGIC; 
  signal MD_13_ENABLE : STD_LOGIC; 
  signal MD_13_TORGTS : STD_LOGIC; 
  signal MD_13_OUTMUX : STD_LOGIC; 
  signal MD_13_OD : STD_LOGIC; 
  signal MD_22_ENABLE : STD_LOGIC; 
  signal MD_22_TORGTS : STD_LOGIC; 
  signal MD_22_OUTMUX : STD_LOGIC; 
  signal MD_22_OD : STD_LOGIC; 
  signal MD_14_ENABLE : STD_LOGIC; 
  signal MD_14_TORGTS : STD_LOGIC; 
  signal MD_14_OUTMUX : STD_LOGIC; 
  signal MD_14_OD : STD_LOGIC; 
  signal MD_30_ENABLE : STD_LOGIC; 
  signal MD_30_TORGTS : STD_LOGIC; 
  signal MD_30_OUTMUX : STD_LOGIC; 
  signal MD_30_OD : STD_LOGIC; 
  signal MACADDR_3_IFF_RST : STD_LOGIC; 
  signal MD_23_ENABLE : STD_LOGIC; 
  signal MD_23_TORGTS : STD_LOGIC; 
  signal MD_23_OUTMUX : STD_LOGIC; 
  signal MD_23_OD : STD_LOGIC; 
  signal MD_15_ENABLE : STD_LOGIC; 
  signal MD_15_TORGTS : STD_LOGIC; 
  signal MD_15_OUTMUX : STD_LOGIC; 
  signal MD_15_OD : STD_LOGIC; 
  signal MD_31_ENABLE : STD_LOGIC; 
  signal MD_31_TORGTS : STD_LOGIC; 
  signal MD_31_OUTMUX : STD_LOGIC; 
  signal MD_31_OD : STD_LOGIC; 
  signal MD_24_ENABLE : STD_LOGIC; 
  signal MD_24_TORGTS : STD_LOGIC; 
  signal MD_24_OUTMUX : STD_LOGIC; 
  signal MD_24_OD : STD_LOGIC; 
  signal MD_16_ENABLE : STD_LOGIC; 
  signal MD_16_TORGTS : STD_LOGIC; 
  signal MD_16_OUTMUX : STD_LOGIC; 
  signal MD_16_OD : STD_LOGIC; 
  signal MD_17_ENABLE : STD_LOGIC; 
  signal MD_17_TORGTS : STD_LOGIC; 
  signal MD_17_OUTMUX : STD_LOGIC; 
  signal MD_17_OD : STD_LOGIC; 
  signal MD_25_ENABLE : STD_LOGIC; 
  signal MD_25_TORGTS : STD_LOGIC; 
  signal MD_25_OUTMUX : STD_LOGIC; 
  signal MD_25_OD : STD_LOGIC; 
  signal MD_18_ENABLE : STD_LOGIC; 
  signal MD_18_TORGTS : STD_LOGIC; 
  signal MD_18_OUTMUX : STD_LOGIC; 
  signal MD_18_OD : STD_LOGIC; 
  signal MD_26_ENABLE : STD_LOGIC; 
  signal MD_26_TORGTS : STD_LOGIC; 
  signal MD_26_OUTMUX : STD_LOGIC; 
  signal MD_26_OD : STD_LOGIC; 
  signal MACADDR_4_IFF_RST : STD_LOGIC; 
  signal MD_19_ENABLE : STD_LOGIC; 
  signal MD_19_TORGTS : STD_LOGIC; 
  signal MD_19_OUTMUX : STD_LOGIC; 
  signal MD_19_OD : STD_LOGIC; 
  signal MD_27_ENABLE : STD_LOGIC; 
  signal MD_27_TORGTS : STD_LOGIC; 
  signal MD_27_OUTMUX : STD_LOGIC; 
  signal MD_27_OD : STD_LOGIC; 
  signal PHYRESET_ENABLE : STD_LOGIC; 
  signal PHYRESET_TORGTS : STD_LOGIC; 
  signal PHYRESET_OUTMUX : STD_LOGIC; 
  signal maccontrol_PHYRESET_OBUF : STD_LOGIC; 
  signal PHYRESET_OD : STD_LOGIC; 
  signal MD_28_ENABLE : STD_LOGIC; 
  signal MD_28_TORGTS : STD_LOGIC; 
  signal MD_28_OUTMUX : STD_LOGIC; 
  signal MD_28_OD : STD_LOGIC; 
  signal MD_29_ENABLE : STD_LOGIC; 
  signal MD_29_TORGTS : STD_LOGIC; 
  signal MD_29_OUTMUX : STD_LOGIC; 
  signal MD_29_OD : STD_LOGIC; 
  signal LED100_ENABLE : STD_LOGIC; 
  signal LED100_TORGTS : STD_LOGIC; 
  signal LED100_OUTMUX : STD_LOGIC; 
  signal maccontrol_LED100_OBUF : STD_LOGIC; 
  signal LED100_OD : STD_LOGIC; 
  signal NEXTF_IBUF_0 : STD_LOGIC; 
  signal RESET_IBUF_1 : STD_LOGIC; 
  signal MDIO_ENABLE : STD_LOGIC; 
  signal MDIO_TORGTS : STD_LOGIC; 
  signal MDIO_OUTMUX : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_sin : STD_LOGIC; 
  signal MACADDR_5_IFF_RST : STD_LOGIC; 
  signal MDC_ENABLE : STD_LOGIC; 
  signal MDC_TORGTS : STD_LOGIC; 
  signal MDC_OUTMUX : STD_LOGIC; 
  signal MOE_ENABLE : STD_LOGIC; 
  signal MOE_TORGTS : STD_LOGIC; 
  signal MOE_OUTMUX : STD_LOGIC; 
  signal MOE_LOGIC_ZERO : STD_LOGIC; 
  signal testrx_RXD_0_IBUF : STD_LOGIC; 
  signal testrx_RXD_1_IBUF : STD_LOGIC; 
  signal testrx_RXD_2_IBUF : STD_LOGIC; 
  signal testrx_RXD_3_IBUF : STD_LOGIC; 
  signal testrx_RXD_4_IBUF : STD_LOGIC; 
  signal testrx_RXD_5_IBUF : STD_LOGIC; 
  signal MWE_ENABLE : STD_LOGIC; 
  signal MWE_TORGTS : STD_LOGIC; 
  signal MWE_OUTMUX : STD_LOGIC; 
  signal memcontroller_WEEXT : STD_LOGIC; 
  signal MWE_OCEMUXNOT : STD_LOGIC; 
  signal MWE_OD : STD_LOGIC; 
  signal MACADDR_6_IFF_RST : STD_LOGIC; 
  signal testrx_RXD_6_IBUF : STD_LOGIC; 
  signal SCS_IBUF_2 : STD_LOGIC; 
  signal testrx_RXD_7_IBUF : STD_LOGIC; 
  signal SIN_IBUF_3 : STD_LOGIC; 
  signal LED1000_ENABLE : STD_LOGIC; 
  signal LED1000_TORGTS : STD_LOGIC; 
  signal LED1000_OUTMUX : STD_LOGIC; 
  signal maccontrol_LED1000_OBUF : STD_LOGIC; 
  signal LED1000_OD : STD_LOGIC; 
  signal RX_ER_IBUF_4 : STD_LOGIC; 
  signal RX_DV_IBUF_5 : STD_LOGIC; 
  signal MACDATA_10_ENABLE : STD_LOGIC; 
  signal MACDATA_10_TORGTS : STD_LOGIC; 
  signal MACDATA_10_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_10_OBUF : STD_LOGIC; 
  signal MACDATA_10_OD : STD_LOGIC; 
  signal MACDATA_11_ENABLE : STD_LOGIC; 
  signal MACDATA_11_TORGTS : STD_LOGIC; 
  signal MACDATA_11_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_11_OBUF : STD_LOGIC; 
  signal MACDATA_11_OD : STD_LOGIC; 
  signal MACADDR_7_IFF_RST : STD_LOGIC; 
  signal MACDATA_12_ENABLE : STD_LOGIC; 
  signal MACDATA_12_TORGTS : STD_LOGIC; 
  signal MACDATA_12_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_12_OBUF : STD_LOGIC; 
  signal MACDATA_12_OD : STD_LOGIC; 
  signal MACDATA_13_ENABLE : STD_LOGIC; 
  signal MACDATA_13_TORGTS : STD_LOGIC; 
  signal MACDATA_13_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_13_OBUF : STD_LOGIC; 
  signal MACDATA_13_OD : STD_LOGIC; 
  signal TX_ER_ENABLE : STD_LOGIC; 
  signal TX_ER_TORGTS : STD_LOGIC; 
  signal TX_ER_OUTMUX : STD_LOGIC; 
  signal TX_ER_LOGIC_ZERO : STD_LOGIC; 
  signal MACDATA_14_ENABLE : STD_LOGIC; 
  signal MACDATA_14_TORGTS : STD_LOGIC; 
  signal MACDATA_14_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_14_OBUF : STD_LOGIC; 
  signal MACDATA_14_OD : STD_LOGIC; 
  signal MACDATA_15_ENABLE : STD_LOGIC; 
  signal MACDATA_15_TORGTS : STD_LOGIC; 
  signal MACDATA_15_OUTMUX : STD_LOGIC; 
  signal testrx_MACDATA_15_OBUF : STD_LOGIC; 
  signal MACDATA_15_OD : STD_LOGIC; 
  signal GTX_CLK_ENABLE : STD_LOGIC; 
  signal GTX_CLK_TORGTS : STD_LOGIC; 
  signal GTX_CLK_OUTMUX : STD_LOGIC; 
  signal LEDTX_ENABLE : STD_LOGIC; 
  signal LEDTX_TORGTS : STD_LOGIC; 
  signal LEDTX_OUTMUX : STD_LOGIC; 
  signal maccontrol_LEDTX_OBUF : STD_LOGIC; 
  signal LEDTX_OD : STD_LOGIC; 
  signal LEDPOWER_ENABLE : STD_LOGIC; 
  signal LEDPOWER_TORGTS : STD_LOGIC; 
  signal LEDPOWER_OUTMUX : STD_LOGIC; 
  signal LEDPOWER_OBUF : STD_LOGIC; 
  signal LEDPOWER_OD : STD_LOGIC; 
  signal ifclk_DLL_LOCKED : STD_LOGIC; 
  signal ifclk_DLL_CLKDV : STD_LOGIC; 
  signal ifclk_DLL_CLK2X180 : STD_LOGIC; 
  signal ifclk_DLL_CLK2X : STD_LOGIC; 
  signal ifclk_DLL_CLK270 : STD_LOGIC; 
  signal ifclk_DLL_CLK180 : STD_LOGIC; 
  signal ifclk_DLL_CLK90 : STD_LOGIC; 
  signal clk_DLL_LOCKED : STD_LOGIC; 
  signal clk_DLL_CLKDV : STD_LOGIC; 
  signal clk_DLL_CLK2X180 : STD_LOGIC; 
  signal clk_DLL_CLK2X : STD_LOGIC; 
  signal clk_DLL_CLK270 : STD_LOGIC; 
  signal rxclk_DLL_LOCKED : STD_LOGIC; 
  signal rxclk_DLL_CLKDV : STD_LOGIC; 
  signal rxclk_DLL_CLK2X180 : STD_LOGIC; 
  signal rxclk_DLL_CLK2X : STD_LOGIC; 
  signal rxclk_DLL_CLK270 : STD_LOGIC; 
  signal rxclk_DLL_CLK180 : STD_LOGIC; 
  signal rxclk_DLL_CLK90 : STD_LOGIC; 
  signal testrx_tempram_DOA15 : STD_LOGIC; 
  signal testrx_tempram_DOA14 : STD_LOGIC; 
  signal testrx_tempram_DOA13 : STD_LOGIC; 
  signal testrx_tempram_DOA12 : STD_LOGIC; 
  signal testrx_tempram_DOA11 : STD_LOGIC; 
  signal testrx_tempram_DOA10 : STD_LOGIC; 
  signal testrx_tempram_DOA9 : STD_LOGIC; 
  signal testrx_tempram_DOA8 : STD_LOGIC; 
  signal testrx_tempram_DOA7 : STD_LOGIC; 
  signal testrx_tempram_DOA6 : STD_LOGIC; 
  signal testrx_tempram_DOA5 : STD_LOGIC; 
  signal testrx_tempram_DOA4 : STD_LOGIC; 
  signal testrx_tempram_DOA3 : STD_LOGIC; 
  signal testrx_tempram_DOA2 : STD_LOGIC; 
  signal testrx_tempram_DOA1 : STD_LOGIC; 
  signal testrx_tempram_DOA0 : STD_LOGIC; 
  signal testrx_tempram_DIA15 : STD_LOGIC; 
  signal testrx_tempram_DIA14 : STD_LOGIC; 
  signal testrx_tempram_DIA13 : STD_LOGIC; 
  signal testrx_tempram_DIA12 : STD_LOGIC; 
  signal testrx_tempram_DIA11 : STD_LOGIC; 
  signal testrx_tempram_DIA10 : STD_LOGIC; 
  signal testrx_tempram_DIA9 : STD_LOGIC; 
  signal testrx_tempram_DIA8 : STD_LOGIC; 
  signal testrx_tempram_ADDRB3 : STD_LOGIC; 
  signal testrx_tempram_ADDRB2 : STD_LOGIC; 
  signal testrx_tempram_ADDRB1 : STD_LOGIC; 
  signal testrx_tempram_ADDRB0 : STD_LOGIC; 
  signal testrx_tempram_ADDRA2 : STD_LOGIC; 
  signal testrx_tempram_ADDRA1 : STD_LOGIC; 
  signal testrx_tempram_ADDRA0 : STD_LOGIC; 
  signal testrx_tempram_LOGIC_ZERO : STD_LOGIC; 
  signal testrx_tempram_LOGIC_ONE : STD_LOGIC; 
  signal txsim_rom_DOB15 : STD_LOGIC; 
  signal txsim_rom_DOB14 : STD_LOGIC; 
  signal txsim_rom_DOB13 : STD_LOGIC; 
  signal txsim_rom_DOB12 : STD_LOGIC; 
  signal txsim_rom_DOB11 : STD_LOGIC; 
  signal txsim_rom_DOB10 : STD_LOGIC; 
  signal txsim_rom_DOB9 : STD_LOGIC; 
  signal txsim_rom_DOB8 : STD_LOGIC; 
  signal txsim_rom_DOB7 : STD_LOGIC; 
  signal txsim_rom_DOB6 : STD_LOGIC; 
  signal txsim_rom_DOB5 : STD_LOGIC; 
  signal txsim_rom_DOB4 : STD_LOGIC; 
  signal txsim_rom_DOB3 : STD_LOGIC; 
  signal txsim_rom_DOB2 : STD_LOGIC; 
  signal txsim_rom_DOB1 : STD_LOGIC; 
  signal txsim_rom_DOB0 : STD_LOGIC; 
  signal txsim_rom_DOA15 : STD_LOGIC; 
  signal txsim_rom_DOA14 : STD_LOGIC; 
  signal txsim_rom_DOA13 : STD_LOGIC; 
  signal txsim_rom_DOA12 : STD_LOGIC; 
  signal txsim_rom_DOA11 : STD_LOGIC; 
  signal txsim_rom_DOA10 : STD_LOGIC; 
  signal txsim_rom_DOA9 : STD_LOGIC; 
  signal txsim_rom_DOA8 : STD_LOGIC; 
  signal txsim_rom_DIB15 : STD_LOGIC; 
  signal txsim_rom_DIB14 : STD_LOGIC; 
  signal txsim_rom_DIB13 : STD_LOGIC; 
  signal txsim_rom_DIB12 : STD_LOGIC; 
  signal txsim_rom_DIB11 : STD_LOGIC; 
  signal txsim_rom_DIB10 : STD_LOGIC; 
  signal txsim_rom_DIB9 : STD_LOGIC; 
  signal txsim_rom_DIB8 : STD_LOGIC; 
  signal txsim_rom_DIB7 : STD_LOGIC; 
  signal txsim_rom_DIB6 : STD_LOGIC; 
  signal txsim_rom_DIB5 : STD_LOGIC; 
  signal txsim_rom_DIB4 : STD_LOGIC; 
  signal txsim_rom_DIB3 : STD_LOGIC; 
  signal txsim_rom_DIB2 : STD_LOGIC; 
  signal txsim_rom_DIB1 : STD_LOGIC; 
  signal txsim_rom_DIB0 : STD_LOGIC; 
  signal txsim_rom_DIA15 : STD_LOGIC; 
  signal txsim_rom_DIA14 : STD_LOGIC; 
  signal txsim_rom_DIA13 : STD_LOGIC; 
  signal txsim_rom_DIA12 : STD_LOGIC; 
  signal txsim_rom_DIA11 : STD_LOGIC; 
  signal txsim_rom_DIA10 : STD_LOGIC; 
  signal txsim_rom_DIA9 : STD_LOGIC; 
  signal txsim_rom_DIA8 : STD_LOGIC; 
  signal txsim_rom_ADDRB11 : STD_LOGIC; 
  signal txsim_rom_ADDRB10 : STD_LOGIC; 
  signal txsim_rom_ADDRB9 : STD_LOGIC; 
  signal txsim_rom_ADDRB8 : STD_LOGIC; 
  signal txsim_rom_ADDRB7 : STD_LOGIC; 
  signal txsim_rom_ADDRB6 : STD_LOGIC; 
  signal txsim_rom_ADDRB5 : STD_LOGIC; 
  signal txsim_rom_ADDRB4 : STD_LOGIC; 
  signal txsim_rom_ADDRB3 : STD_LOGIC; 
  signal txsim_rom_ADDRB2 : STD_LOGIC; 
  signal txsim_rom_ADDRB1 : STD_LOGIC; 
  signal txsim_rom_ADDRB0 : STD_LOGIC; 
  signal txsim_rom_ADDRA2 : STD_LOGIC; 
  signal txsim_rom_ADDRA1 : STD_LOGIC; 
  signal txsim_rom_ADDRA0 : STD_LOGIC; 
  signal txsim_rom_LOGIC_ZERO : STD_LOGIC; 
  signal txsim_rom_LOGIC_ONE : STD_LOGIC; 
  signal memcontroller_N46782 : STD_LOGIC; 
  signal memcontroller_N46780 : STD_LOGIC; 
  signal memcontroller_addrn_0_F5MUX : STD_LOGIC; 
  signal memcontroller_N46792 : STD_LOGIC; 
  signal memcontroller_N46790 : STD_LOGIC; 
  signal memcontroller_addrn_2_F5MUX : STD_LOGIC; 
  signal memcontroller_N46797 : STD_LOGIC; 
  signal memcontroller_N46795 : STD_LOGIC; 
  signal memcontroller_addrn_3_F5MUX : STD_LOGIC; 
  signal memcontroller_N46802 : STD_LOGIC; 
  signal memcontroller_N46800 : STD_LOGIC; 
  signal memcontroller_addrn_4_F5MUX : STD_LOGIC; 
  signal memcontroller_N46787 : STD_LOGIC; 
  signal memcontroller_N46785 : STD_LOGIC; 
  signal memcontroller_addrn_1_F5MUX : STD_LOGIC; 
  signal memcontroller_N46807 : STD_LOGIC; 
  signal memcontroller_N46805 : STD_LOGIC; 
  signal memcontroller_addrn_5_F5MUX : STD_LOGIC; 
  signal MA_0_OFF_RST : STD_LOGIC; 
  signal memcontroller_N46812 : STD_LOGIC; 
  signal memcontroller_N46810 : STD_LOGIC; 
  signal memcontroller_addrn_6_F5MUX : STD_LOGIC; 
  signal memcontroller_N46817 : STD_LOGIC; 
  signal memcontroller_N46815 : STD_LOGIC; 
  signal memcontroller_addrn_7_F5MUX : STD_LOGIC; 
  signal memcontroller_N46822 : STD_LOGIC; 
  signal memcontroller_N46820 : STD_LOGIC; 
  signal memcontroller_addrn_8_F5MUX : STD_LOGIC; 
  signal memcontroller_N46827 : STD_LOGIC; 
  signal memcontroller_N46825 : STD_LOGIC; 
  signal memcontroller_addrn_9_F5MUX : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N46762 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N46760 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE826_F5MUX : STD_LOGIC; 
  signal memcontroller_N46832 : STD_LOGIC; 
  signal memcontroller_N46830 : STD_LOGIC; 
  signal memcontroller_addrn_10_F5MUX : STD_LOGIC; 
  signal memcontroller_N46837 : STD_LOGIC; 
  signal memcontroller_N46835 : STD_LOGIC; 
  signal memcontroller_addrn_11_F5MUX : STD_LOGIC; 
  signal memcontroller_N46842 : STD_LOGIC; 
  signal memcontroller_N46840 : STD_LOGIC; 
  signal memcontroller_addrn_12_F5MUX : STD_LOGIC; 
  signal memcontroller_N46847 : STD_LOGIC; 
  signal memcontroller_N46845 : STD_LOGIC; 
  signal memcontroller_addrn_13_F5MUX : STD_LOGIC; 
  signal memcontroller_N46767 : STD_LOGIC; 
  signal memcontroller_N46765 : STD_LOGIC; 
  signal memcontroller_addrn_14_F5MUX : STD_LOGIC; 
  signal memcontroller_N46772 : STD_LOGIC; 
  signal memcontroller_N46770 : STD_LOGIC; 
  signal memcontroller_addrn_15_F5MUX : STD_LOGIC; 
  signal memcontroller_clknum_1_2_rt : STD_LOGIC; 
  signal memcontroller_N46775 : STD_LOGIC; 
  signal memcontroller_addrn_16_F5MUX : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_155 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_123_CYMUXG : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_123_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_156 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_224 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_123_LOGIC_ZERO : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_178 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_157 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_179 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_125_CYMUXG : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_125_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_158 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_226 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_125_CYINIT : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_180 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_159 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_181 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_127_CYMUXG : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_127_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_160 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_228 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_127_CYINIT : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_182 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_161 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_183 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_129_CYMUXG : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_129_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_162 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_230 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_129_CYINIT : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_184 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_163 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_185 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_131_CYMUXG : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_131_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_164 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_232 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_131_CYINIT : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_186 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_133_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_165 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_187 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_lut3_166 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_cy_234 : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_133_CYINIT : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_inst_sum_188 : STD_LOGIC; 
  signal maccontrol_Mshreg_scslll_84_rt : STD_LOGIC; 
  signal maccontrol_bitcnt_85_CYMUXG : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_lut3_117 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_cy_183 : STD_LOGIC; 
  signal maccontrol_bitcnt_85_LOGIC_ZERO : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_sum_139 : STD_LOGIC; 
  signal MA_1_OFF_RST : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_lut3_118 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_sum_140 : STD_LOGIC; 
  signal maccontrol_bitcnt_86_CYMUXG : STD_LOGIC; 
  signal maccontrol_bitcnt_86_LOGIC_ZERO : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_lut3_119 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_cy_185 : STD_LOGIC; 
  signal maccontrol_bitcnt_86_CYINIT : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_sum_141 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_lut3_120 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_sum_142 : STD_LOGIC; 
  signal maccontrol_bitcnt_88_CYMUXG : STD_LOGIC; 
  signal maccontrol_bitcnt_88_LOGIC_ZERO : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_lut3_121 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_cy_187 : STD_LOGIC; 
  signal maccontrol_bitcnt_88_CYINIT : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_sum_143 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_lut3_122 : STD_LOGIC; 
  signal maccontrol_bitcnt_inst_sum_144 : STD_LOGIC; 
  signal maccontrol_bitcnt_90_GROM : STD_LOGIC; 
  signal maccontrol_bitcnt_90_CYINIT : STD_LOGIC; 
  signal maccontrol_N30228_rt : STD_LOGIC; 
  signal maccontrol_phyrstcnt_91_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_91_GROM : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_190 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_91_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_145 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1241_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_146 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_92_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_92_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1251_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_192 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_92_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_147 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1261_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_148 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_94_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_94_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1271_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_194 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_94_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_149 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1281_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_150 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_96_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_96_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1291_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_196 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_96_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_151 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1301_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_152 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_98_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_98_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1311_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_198 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_98_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_153 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1321_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_154 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_100_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_100_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1331_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_200 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_100_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_155 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1341_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_156 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_102_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_102_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1351_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_202 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_102_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_157 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1361_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_158 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_104_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_104_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1371_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_204 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_104_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_159 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1381_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_160 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_106_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_106_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1391_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_206 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_106_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_161 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1401_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_162 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_108_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_108_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1411_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_208 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_108_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_163 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1421_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_164 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_110_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_110_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1431_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_210 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_110_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_165 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1441_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_166 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_112_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_112_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1451_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_212 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_112_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_167 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1461_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_168 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_114_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_114_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1471_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_214 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_114_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_169 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1481_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_170 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_116_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_116_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1491_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_216 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_116_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_171 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1501_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_172 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_118_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_118_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1511_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_218 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_118_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_173 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1521_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_174 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_120_CYMUXG : STD_LOGIC; 
  signal maccontrol_phyrstcnt_120_LOGIC_ONE : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1531_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_cy_220 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_120_CYINIT : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_175 : STD_LOGIC; 
  signal MA_2_OFF_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_lut3_1541_O : STD_LOGIC; 
  signal maccontrol_phyrstcnt_inst_sum_176 : STD_LOGIC; 
  signal maccontrol_phyrstcnt_122_GROM : STD_LOGIC; 
  signal maccontrol_phyrstcnt_122_CYINIT : STD_LOGIC; 
  signal cnt0_Madd_n0000_inst_lut2_24 : STD_LOGIC; 
  signal cnt0_0_CYMUXG : STD_LOGIC; 
  signal cnt0_0_GROM : STD_LOGIC; 
  signal cnt0_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal cnt0_0_LOGIC_ZERO : STD_LOGIC; 
  signal cnt0_2_FROM : STD_LOGIC; 
  signal cnt0_2_CYMUXG : STD_LOGIC; 
  signal cnt0_2_LOGIC_ZERO : STD_LOGIC; 
  signal cnt0_2_GROM : STD_LOGIC; 
  signal cnt0_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal cnt0_2_CYINIT : STD_LOGIC; 
  signal cnt0_4_LOGIC_ZERO : STD_LOGIC; 
  signal cnt0_4_FROM : STD_LOGIC; 
  signal cnt0_5_rt : STD_LOGIC; 
  signal cnt0_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal cnt0_4_CYINIT : STD_LOGIC; 
  signal memtest2_Mcompar_n0020_inst_lut4_25 : STD_LOGIC; 
  signal memtest2_Mcompar_n0020_inst_cy_167_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0020_inst_lut4_26 : STD_LOGIC; 
  signal memtest2_Mcompar_n0020_inst_cy_166 : STD_LOGIC; 
  signal memtest2_Mcompar_n0020_inst_cy_167_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_Mcompar_n0020_inst_cy_167_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_Mcompar_n0020_inst_lut4_27 : STD_LOGIC; 
  signal memtest2_deq_3_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0020_inst_lut4_28 : STD_LOGIC; 
  signal memtest2_Mcompar_n0020_inst_cy_168 : STD_LOGIC; 
  signal memtest2_deq_3_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_deq_3_CYINIT : STD_LOGIC; 
  signal Madd_n0000_inst_lut2_0 : STD_LOGIC; 
  signal cnt_0_CYMUXG : STD_LOGIC; 
  signal cnt_0_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_0 : STD_LOGIC; 
  signal cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_2_FROM : STD_LOGIC; 
  signal cnt_2_CYMUXG : STD_LOGIC; 
  signal cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_2_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_2 : STD_LOGIC; 
  signal cnt_2_CYINIT : STD_LOGIC; 
  signal cnt_4_FROM : STD_LOGIC; 
  signal cnt_4_CYMUXG : STD_LOGIC; 
  signal cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_4_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_4 : STD_LOGIC; 
  signal cnt_4_CYINIT : STD_LOGIC; 
  signal cnt_6_FROM : STD_LOGIC; 
  signal cnt_6_CYMUXG : STD_LOGIC; 
  signal cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_6_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_6 : STD_LOGIC; 
  signal cnt_6_CYINIT : STD_LOGIC; 
  signal cnt_8_FROM : STD_LOGIC; 
  signal cnt_8_CYMUXG : STD_LOGIC; 
  signal cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_8_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_8 : STD_LOGIC; 
  signal cnt_8_CYINIT : STD_LOGIC; 
  signal cnt_10_FROM : STD_LOGIC; 
  signal cnt_10_CYMUXG : STD_LOGIC; 
  signal cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_10_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_10 : STD_LOGIC; 
  signal cnt_10_CYINIT : STD_LOGIC; 
  signal cnt_12_FROM : STD_LOGIC; 
  signal cnt_12_CYMUXG : STD_LOGIC; 
  signal cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_12_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_12 : STD_LOGIC; 
  signal cnt_12_CYINIT : STD_LOGIC; 
  signal cnt_14_FROM : STD_LOGIC; 
  signal cnt_14_CYMUXG : STD_LOGIC; 
  signal cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_14_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_14 : STD_LOGIC; 
  signal cnt_14_CYINIT : STD_LOGIC; 
  signal cnt_16_FROM : STD_LOGIC; 
  signal cnt_16_CYMUXG : STD_LOGIC; 
  signal cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_16_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal cnt_16_CYINIT : STD_LOGIC; 
  signal cnt_18_FROM : STD_LOGIC; 
  signal cnt_18_CYMUXG : STD_LOGIC; 
  signal cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_18_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal cnt_18_CYINIT : STD_LOGIC; 
  signal cnt_20_FROM : STD_LOGIC; 
  signal cnt_20_CYMUXG : STD_LOGIC; 
  signal cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_20_GROM : STD_LOGIC; 
  signal Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal cnt_20_CYINIT : STD_LOGIC; 
  signal cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal cnt_22_FROM : STD_LOGIC; 
  signal cnt_23_rt : STD_LOGIC; 
  signal Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal cnt_22_CYINIT : STD_LOGIC; 
  signal cnt_22_XORG : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd5_rt : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_0_CYMUXG : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_0 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_121 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_121 : STD_LOGIC; 
  signal MA_3_OFF_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_1 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_122 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_1_CYMUXG : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_1_LOGIC_ZERO : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_2 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_123 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_1_CYINIT : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_123 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_3 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_124 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_3_CYMUXG : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_3_LOGIC_ZERO : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_4 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_125 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_3_CYINIT : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_125 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_5 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_126 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_5_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_5_CYINIT : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_0 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_129_CYMUXG : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_1 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_128 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_129_LOGIC_ZERO : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_129_LOGIC_ONE : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_2 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_131_CYMUXG : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_3 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_130 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_131_LOGIC_ZERO : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_131_CYINIT : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_4 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_133_CYMUXG : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_5 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_132 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_133_LOGIC_ZERO : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_133_CYINIT : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_6 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_135_CYMUXG : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_7 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_134 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_135_LOGIC_ZERO : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_135_CYINIT : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_8 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_137_CYMUXG : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_9 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_136 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_137_LOGIC_ZERO : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_137_CYINIT : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_10 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_139_CYMUXG : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_11 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_138 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_139_LOGIC_ZERO : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_139_CYINIT : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_12 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_141_CYMUXG : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_13 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_140 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_141_LOGIC_ZERO : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_141_CYINIT : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_14 : STD_LOGIC; 
  signal memtest_n0002_CYMUXG : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_lut4_15 : STD_LOGIC; 
  signal memtest_Mcompar_n0002_inst_cy_142 : STD_LOGIC; 
  signal memtest_n0002_LOGIC_ZERO : STD_LOGIC; 
  signal memtest_n0002_CYINIT : STD_LOGIC; 
  signal testrx_addr_Madd_n0000_inst_lut2_30 : STD_LOGIC; 
  signal testrx_addr_0_CYMUXG : STD_LOGIC; 
  signal testrx_addr_0_GROM : STD_LOGIC; 
  signal testrx_addr_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal testrx_addr_0_LOGIC_ZERO : STD_LOGIC; 
  signal testrx_addr_2_FROM : STD_LOGIC; 
  signal testrx_addr_2_CYMUXG : STD_LOGIC; 
  signal testrx_addr_2_LOGIC_ZERO : STD_LOGIC; 
  signal testrx_addr_2_GROM : STD_LOGIC; 
  signal testrx_addr_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal testrx_addr_2_CYINIT : STD_LOGIC; 
  signal testrx_addr_4_FROM : STD_LOGIC; 
  signal testrx_addr_4_CYMUXG : STD_LOGIC; 
  signal testrx_addr_4_LOGIC_ZERO : STD_LOGIC; 
  signal testrx_addr_4_GROM : STD_LOGIC; 
  signal testrx_addr_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal testrx_addr_4_CYINIT : STD_LOGIC; 
  signal testrx_addr_6_LOGIC_ZERO : STD_LOGIC; 
  signal testrx_addr_6_FROM : STD_LOGIC; 
  signal testrx_addr_7_rt : STD_LOGIC; 
  signal testrx_addr_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal testrx_addr_6_CYINIT : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_lut2_86 : STD_LOGIC; 
  signal memtest2_cnt_0_CYMUXG : STD_LOGIC; 
  signal memtest2_cnt_0_GROM : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_86 : STD_LOGIC; 
  signal memtest2_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_cnt_2_FROM : STD_LOGIC; 
  signal memtest2_cnt_2_CYMUXG : STD_LOGIC; 
  signal memtest2_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_cnt_2_GROM : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_88 : STD_LOGIC; 
  signal memtest2_cnt_2_CYINIT : STD_LOGIC; 
  signal memtest2_cnt_4_FROM : STD_LOGIC; 
  signal memtest2_cnt_4_CYMUXG : STD_LOGIC; 
  signal memtest2_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_cnt_4_GROM : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_90 : STD_LOGIC; 
  signal memtest2_cnt_4_CYINIT : STD_LOGIC; 
  signal memtest2_cnt_6_FROM : STD_LOGIC; 
  signal memtest2_cnt_6_CYMUXG : STD_LOGIC; 
  signal memtest2_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_cnt_6_GROM : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_92 : STD_LOGIC; 
  signal memtest2_cnt_6_CYINIT : STD_LOGIC; 
  signal MA_4_OFF_RST : STD_LOGIC; 
  signal memtest2_cnt_8_FROM : STD_LOGIC; 
  signal memtest2_cnt_8_CYMUXG : STD_LOGIC; 
  signal memtest2_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_cnt_8_GROM : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_94 : STD_LOGIC; 
  signal memtest2_cnt_8_CYINIT : STD_LOGIC; 
  signal memtest2_cnt_10_FROM : STD_LOGIC; 
  signal memtest2_cnt_10_CYMUXG : STD_LOGIC; 
  signal memtest2_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_cnt_10_GROM : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_96 : STD_LOGIC; 
  signal memtest2_cnt_10_CYINIT : STD_LOGIC; 
  signal memtest2_cnt_12_FROM : STD_LOGIC; 
  signal memtest2_cnt_12_CYMUXG : STD_LOGIC; 
  signal memtest2_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_cnt_12_GROM : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_98 : STD_LOGIC; 
  signal memtest2_cnt_12_CYINIT : STD_LOGIC; 
  signal memtest2_cnt_14_FROM : STD_LOGIC; 
  signal memtest2_cnt_14_CYMUXG : STD_LOGIC; 
  signal memtest2_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_cnt_14_GROM : STD_LOGIC; 
  signal memtest2_cnt_Madd_n0000_inst_cy_100 : STD_LOGIC; 
  signal memtest2_cnt_14_CYINIT : STD_LOGIC; 
  signal memtest2_cnt_16_rt : STD_LOGIC; 
  signal memtest2_cnt_16_CYINIT : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_lut4_22 : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_161_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_lut4_23 : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_160 : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_161_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_161_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_lut4_24 : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_163_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_lut3_6 : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_162 : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_163_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_163_CYINIT : STD_LOGIC; 
  signal memtest2_SIG_0 : STD_LOGIC; 
  signal memtest2_n0025_CYMUXG : STD_LOGIC; 
  signal memtest2_SIG_1 : STD_LOGIC; 
  signal memtest2_Mcompar_n0025_inst_cy_164 : STD_LOGIC; 
  signal memtest2_n0025_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_n0025_CYINIT : STD_LOGIC; 
  signal memtest2_Mcompar_n0017_inst_lut4_25 : STD_LOGIC; 
  signal memtest2_Mcompar_n0017_inst_cy_167_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0017_inst_lut4_26 : STD_LOGIC; 
  signal memtest2_Mcompar_n0017_inst_cy_166 : STD_LOGIC; 
  signal memtest2_Mcompar_n0017_inst_cy_167_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_Mcompar_n0017_inst_cy_167_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_Mcompar_n0017_inst_lut4_27 : STD_LOGIC; 
  signal memtest2_deq_0_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0017_inst_lut4_28 : STD_LOGIC; 
  signal memtest2_Mcompar_n0017_inst_cy_168 : STD_LOGIC; 
  signal memtest2_deq_0_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_deq_0_CYINIT : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_lut2_24 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_1_CYMUXG : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_1_XORG : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_1_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_24 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_1_LOGIC_ZERO : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_2_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_2_XORF : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_2_CYMUXG : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_2_LOGIC_ZERO : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_2_XORG : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_2_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_26 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_2_CYINIT : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_4_LOGIC_ZERO : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_4_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_4_XORF : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_4_XORG : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_statecnt_5_rt : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_28 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0078_4_CYINIT : STD_LOGIC; 
  signal memtest2_Mcompar_n0018_inst_lut4_25 : STD_LOGIC; 
  signal memtest2_Mcompar_n0018_inst_cy_167_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0018_inst_lut4_26 : STD_LOGIC; 
  signal memtest2_Mcompar_n0018_inst_cy_166 : STD_LOGIC; 
  signal memtest2_Mcompar_n0018_inst_cy_167_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_Mcompar_n0018_inst_cy_167_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_Mcompar_n0018_inst_lut4_27 : STD_LOGIC; 
  signal memtest2_deq_1_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0018_inst_lut4_28 : STD_LOGIC; 
  signal memtest2_Mcompar_n0018_inst_cy_168 : STD_LOGIC; 
  signal memtest2_deq_1_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_deq_1_CYINIT : STD_LOGIC; 
  signal memtest2_SIG_2 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_153_CYMUXG : STD_LOGIC; 
  signal memtest2_SIG_3 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_152 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_153_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_153_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_lut4_19 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_155_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_lut4_20 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_154 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_155_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_155_CYINIT : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_lut4_21 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_157_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_lut2_124 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_156 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_157_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_157_CYINIT : STD_LOGIC; 
  signal memtest2_SIG_4 : STD_LOGIC; 
  signal memtest2_n0027_CYMUXG : STD_LOGIC; 
  signal memtest2_SIG_5 : STD_LOGIC; 
  signal memtest2_Mcompar_n0027_inst_cy_158 : STD_LOGIC; 
  signal memtest2_n0027_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_n0027_CYINIT : STD_LOGIC; 
  signal MA_5_OFF_RST : STD_LOGIC; 
  signal memtest2_Mcompar_n0019_inst_lut4_25 : STD_LOGIC; 
  signal memtest2_Mcompar_n0019_inst_cy_167_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0019_inst_lut4_26 : STD_LOGIC; 
  signal memtest2_Mcompar_n0019_inst_cy_166 : STD_LOGIC; 
  signal memtest2_Mcompar_n0019_inst_cy_167_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_Mcompar_n0019_inst_cy_167_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_Mcompar_n0019_inst_lut4_27 : STD_LOGIC; 
  signal memtest2_deq_2_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0019_inst_lut4_28 : STD_LOGIC; 
  signal memtest2_Mcompar_n0019_inst_cy_168 : STD_LOGIC; 
  signal memtest2_deq_2_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_deq_2_CYINIT : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_lut2_103 : STD_LOGIC; 
  signal txsim_counter_0_CYMUXG : STD_LOGIC; 
  signal txsim_counter_0_GROM : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_103 : STD_LOGIC; 
  signal txsim_counter_0_LOGIC_ZERO : STD_LOGIC; 
  signal txsim_counter_2_FROM : STD_LOGIC; 
  signal txsim_counter_2_CYMUXG : STD_LOGIC; 
  signal txsim_counter_2_LOGIC_ZERO : STD_LOGIC; 
  signal txsim_counter_2_GROM : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_105 : STD_LOGIC; 
  signal txsim_counter_2_CYINIT : STD_LOGIC; 
  signal txsim_counter_4_FROM : STD_LOGIC; 
  signal txsim_counter_4_CYMUXG : STD_LOGIC; 
  signal txsim_counter_4_LOGIC_ZERO : STD_LOGIC; 
  signal txsim_counter_4_GROM : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_107 : STD_LOGIC; 
  signal txsim_counter_4_CYINIT : STD_LOGIC; 
  signal txsim_counter_6_FROM : STD_LOGIC; 
  signal txsim_counter_6_CYMUXG : STD_LOGIC; 
  signal txsim_counter_6_LOGIC_ZERO : STD_LOGIC; 
  signal txsim_counter_6_GROM : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_109 : STD_LOGIC; 
  signal txsim_counter_6_CYINIT : STD_LOGIC; 
  signal txsim_counter_8_FROM : STD_LOGIC; 
  signal txsim_counter_8_CYMUXG : STD_LOGIC; 
  signal txsim_counter_8_LOGIC_ZERO : STD_LOGIC; 
  signal txsim_counter_8_GROM : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_111 : STD_LOGIC; 
  signal txsim_counter_8_CYINIT : STD_LOGIC; 
  signal txsim_counter_10_FROM : STD_LOGIC; 
  signal txsim_counter_10_CYMUXG : STD_LOGIC; 
  signal txsim_counter_10_LOGIC_ZERO : STD_LOGIC; 
  signal txsim_counter_10_GROM : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_113 : STD_LOGIC; 
  signal txsim_counter_10_CYINIT : STD_LOGIC; 
  signal txsim_counter_12_FROM : STD_LOGIC; 
  signal txsim_counter_12_CYMUXG : STD_LOGIC; 
  signal txsim_counter_12_LOGIC_ZERO : STD_LOGIC; 
  signal txsim_counter_12_GROM : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_115 : STD_LOGIC; 
  signal txsim_counter_12_CYINIT : STD_LOGIC; 
  signal txsim_counter_14_FROM : STD_LOGIC; 
  signal txsim_counter_14_CYMUXG : STD_LOGIC; 
  signal txsim_counter_14_LOGIC_ZERO : STD_LOGIC; 
  signal txsim_counter_14_GROM : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_117 : STD_LOGIC; 
  signal txsim_counter_14_CYINIT : STD_LOGIC; 
  signal txsim_counter_16_LOGIC_ZERO : STD_LOGIC; 
  signal txsim_counter_16_FROM : STD_LOGIC; 
  signal txsim_counter_17_rt : STD_LOGIC; 
  signal txsim_counter_Madd_n0000_inst_cy_119 : STD_LOGIC; 
  signal txsim_counter_16_CYINIT : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut1_0 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_145_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut1_1 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_144 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_145_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_145_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut2_121 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_147_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut2_122 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_146 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_147_LOGIC_ONE : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_147_CYINIT : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut4_16_FROM : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut4_16_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut4_17 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_148 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut4_16_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut4_16_CYINIT : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut4_18 : STD_LOGIC; 
  signal memtest2_n0028_CYMUXG : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_lut2_123 : STD_LOGIC; 
  signal memtest2_Mcompar_n0028_inst_cy_150 : STD_LOGIC; 
  signal memtest2_n0028_LOGIC_ZERO : STD_LOGIC; 
  signal memtest2_n0028_CYINIT : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_lut2_38 : STD_LOGIC; 
  signal d1_0_CYMUXG : STD_LOGIC; 
  signal d1_0_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal d1_0_LOGIC_ZERO : STD_LOGIC; 
  signal d1_2_FROM : STD_LOGIC; 
  signal d1_2_CYMUXG : STD_LOGIC; 
  signal d1_2_LOGIC_ZERO : STD_LOGIC; 
  signal d1_2_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal d1_2_CYINIT : STD_LOGIC; 
  signal d1_4_FROM : STD_LOGIC; 
  signal d1_4_CYMUXG : STD_LOGIC; 
  signal d1_4_LOGIC_ZERO : STD_LOGIC; 
  signal d1_4_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal d1_4_CYINIT : STD_LOGIC; 
  signal d1_6_FROM : STD_LOGIC; 
  signal d1_6_CYMUXG : STD_LOGIC; 
  signal d1_6_LOGIC_ZERO : STD_LOGIC; 
  signal d1_6_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal d1_6_CYINIT : STD_LOGIC; 
  signal MA_6_OFF_RST : STD_LOGIC; 
  signal d1_8_FROM : STD_LOGIC; 
  signal d1_8_CYMUXG : STD_LOGIC; 
  signal d1_8_LOGIC_ZERO : STD_LOGIC; 
  signal d1_8_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal d1_8_CYINIT : STD_LOGIC; 
  signal d1_10_FROM : STD_LOGIC; 
  signal d1_10_CYMUXG : STD_LOGIC; 
  signal d1_10_LOGIC_ZERO : STD_LOGIC; 
  signal d1_10_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_48 : STD_LOGIC; 
  signal d1_10_CYINIT : STD_LOGIC; 
  signal d1_12_FROM : STD_LOGIC; 
  signal d1_12_CYMUXG : STD_LOGIC; 
  signal d1_12_LOGIC_ZERO : STD_LOGIC; 
  signal d1_12_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_50 : STD_LOGIC; 
  signal d1_12_CYINIT : STD_LOGIC; 
  signal d1_14_FROM : STD_LOGIC; 
  signal d1_14_CYMUXG : STD_LOGIC; 
  signal d1_14_LOGIC_ZERO : STD_LOGIC; 
  signal d1_14_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_52 : STD_LOGIC; 
  signal d1_14_CYINIT : STD_LOGIC; 
  signal d1_16_FROM : STD_LOGIC; 
  signal d1_16_CYMUXG : STD_LOGIC; 
  signal d1_16_LOGIC_ZERO : STD_LOGIC; 
  signal d1_16_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_54 : STD_LOGIC; 
  signal d1_16_CYINIT : STD_LOGIC; 
  signal d1_18_FROM : STD_LOGIC; 
  signal d1_18_CYMUXG : STD_LOGIC; 
  signal d1_18_LOGIC_ZERO : STD_LOGIC; 
  signal d1_18_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_56 : STD_LOGIC; 
  signal d1_18_CYINIT : STD_LOGIC; 
  signal d1_20_FROM : STD_LOGIC; 
  signal d1_20_CYMUXG : STD_LOGIC; 
  signal d1_20_LOGIC_ZERO : STD_LOGIC; 
  signal d1_20_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_58 : STD_LOGIC; 
  signal d1_20_CYINIT : STD_LOGIC; 
  signal d1_22_FROM : STD_LOGIC; 
  signal d1_22_CYMUXG : STD_LOGIC; 
  signal d1_22_LOGIC_ZERO : STD_LOGIC; 
  signal d1_22_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_60 : STD_LOGIC; 
  signal d1_22_CYINIT : STD_LOGIC; 
  signal d1_24_FROM : STD_LOGIC; 
  signal d1_24_CYMUXG : STD_LOGIC; 
  signal d1_24_LOGIC_ZERO : STD_LOGIC; 
  signal d1_24_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_62 : STD_LOGIC; 
  signal d1_24_CYINIT : STD_LOGIC; 
  signal d1_26_FROM : STD_LOGIC; 
  signal d1_26_CYMUXG : STD_LOGIC; 
  signal d1_26_LOGIC_ZERO : STD_LOGIC; 
  signal d1_26_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_64 : STD_LOGIC; 
  signal d1_26_CYINIT : STD_LOGIC; 
  signal d1_28_FROM : STD_LOGIC; 
  signal d1_28_CYMUXG : STD_LOGIC; 
  signal d1_28_LOGIC_ZERO : STD_LOGIC; 
  signal d1_28_GROM : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_66 : STD_LOGIC; 
  signal d1_28_CYINIT : STD_LOGIC; 
  signal d1_30_LOGIC_ZERO : STD_LOGIC; 
  signal d1_30_FROM : STD_LOGIC; 
  signal d1_31_rt : STD_LOGIC; 
  signal memtest_datacnt_Madd_n0000_inst_cy_68 : STD_LOGIC; 
  signal d1_30_CYINIT : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_lut2_70 : STD_LOGIC; 
  signal addr1_0_CYMUXG : STD_LOGIC; 
  signal addr1_0_GROM : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_70 : STD_LOGIC; 
  signal addr1_0_LOGIC_ZERO : STD_LOGIC; 
  signal addr1_2_FROM : STD_LOGIC; 
  signal addr1_2_CYMUXG : STD_LOGIC; 
  signal addr1_2_LOGIC_ZERO : STD_LOGIC; 
  signal addr1_2_GROM : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_72 : STD_LOGIC; 
  signal addr1_2_CYINIT : STD_LOGIC; 
  signal addr1_4_FROM : STD_LOGIC; 
  signal addr1_4_CYMUXG : STD_LOGIC; 
  signal addr1_4_LOGIC_ZERO : STD_LOGIC; 
  signal addr1_4_GROM : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_74 : STD_LOGIC; 
  signal addr1_4_CYINIT : STD_LOGIC; 
  signal addr1_6_FROM : STD_LOGIC; 
  signal addr1_6_CYMUXG : STD_LOGIC; 
  signal addr1_6_LOGIC_ZERO : STD_LOGIC; 
  signal addr1_6_GROM : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_76 : STD_LOGIC; 
  signal addr1_6_CYINIT : STD_LOGIC; 
  signal addr1_8_FROM : STD_LOGIC; 
  signal addr1_8_CYMUXG : STD_LOGIC; 
  signal addr1_8_LOGIC_ZERO : STD_LOGIC; 
  signal addr1_8_GROM : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_78 : STD_LOGIC; 
  signal addr1_8_CYINIT : STD_LOGIC; 
  signal addr1_10_FROM : STD_LOGIC; 
  signal addr1_10_CYMUXG : STD_LOGIC; 
  signal addr1_10_LOGIC_ZERO : STD_LOGIC; 
  signal addr1_10_GROM : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_80 : STD_LOGIC; 
  signal addr1_10_CYINIT : STD_LOGIC; 
  signal addr1_12_FROM : STD_LOGIC; 
  signal addr1_12_CYMUXG : STD_LOGIC; 
  signal addr1_12_LOGIC_ZERO : STD_LOGIC; 
  signal addr1_12_GROM : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_82 : STD_LOGIC; 
  signal addr1_12_CYINIT : STD_LOGIC; 
  signal MA_7_OFF_RST : STD_LOGIC; 
  signal addr1_14_LOGIC_ZERO : STD_LOGIC; 
  signal addr1_14_FROM : STD_LOGIC; 
  signal addr1_15_rt : STD_LOGIC; 
  signal memtest_addrcnt_Madd_n0000_inst_cy_84 : STD_LOGIC; 
  signal addr1_14_CYINIT : STD_LOGIC; 
  signal addr2_13_FROM : STD_LOGIC; 
  signal addr2_13_GROM : STD_LOGIC; 
  signal memtest2_datain_11_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_11_GROM : STD_LOGIC; 
  signal memtest2_datain_30_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_30_FROM : STD_LOGIC; 
  signal memtest2_Mshreg_data4_10_net107 : STD_LOGIC; 
  signal maccontrol_dout_0_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_0_92_O : STD_LOGIC; 
  signal maccontrol_dout_14_FFY_RST : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_14_58_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_1_58_O : STD_LOGIC; 
  signal maccontrol_dout_2_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_2_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_2_58_O : STD_LOGIC; 
  signal maccontrol_dout_3_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_3_76_O : STD_LOGIC; 
  signal maccontrol_dout_4_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_4_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_4_68_O : STD_LOGIC; 
  signal maccontrol_dout_5_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_5_58_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_8_58_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_6_58_O : STD_LOGIC; 
  signal maccontrol_dout_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_7_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_7_76_O : STD_LOGIC; 
  signal d2_0_GROM : STD_LOGIC; 
  signal maccontrol_dout_9_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_9_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_9_68_O : STD_LOGIC; 
  signal d2_3_GROM : STD_LOGIC; 
  signal memtest2_Mshreg_data4_13_56_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_13_56_FROM : STD_LOGIC; 
  signal memtest2_Mshreg_data4_20_net87 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_21_48_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_21_48_FROM : STD_LOGIC; 
  signal memtest2_Mshreg_data4_24_net79 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_13_18_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_13_18_O_GROM : STD_LOGIC; 
  signal maccontrol_dout_10_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_10_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_10_58_O : STD_LOGIC; 
  signal MA_8_OFF_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_phyaddrws_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_phyaddrws_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_phyaddrws_BYMUXNOT : STD_LOGIC; 
  signal maccontrol_dout_11_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_11_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_11_76_O : STD_LOGIC; 
  signal maccontrol_dout_12_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_12_68_O : STD_LOGIC; 
  signal maccontrol_dout_20_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_20_22_O : STD_LOGIC; 
  signal maccontrol_dout_21_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_21_36_O : STD_LOGIC; 
  signal maccontrol_dout_13_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_13_68_O : STD_LOGIC; 
  signal maccontrol_dout_30_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_30_22_O : STD_LOGIC; 
  signal maccontrol_dout_22_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_22_22_O : STD_LOGIC; 
  signal maccontrol_dout_23_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_23_25_O : STD_LOGIC; 
  signal maccontrol_dout_31_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_31_25_O : STD_LOGIC; 
  signal maccontrol_dout_15_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_15_76_O : STD_LOGIC; 
  signal maccontrol_dout_24_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_24_36_O : STD_LOGIC; 
  signal maccontrol_dout_16_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_16_36_O : STD_LOGIC; 
  signal maccontrol_dout_17_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_17_36_O : STD_LOGIC; 
  signal maccontrol_dout_25_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_25_22_O : STD_LOGIC; 
  signal maccontrol_dout_18_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_18_22_O : STD_LOGIC; 
  signal maccontrol_dout_26_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_26_22_O : STD_LOGIC; 
  signal maccontrol_dout_27_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_27_25_O : STD_LOGIC; 
  signal maccontrol_dout_19_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_19_25_O : STD_LOGIC; 
  signal MA_9_OFF_RST : STD_LOGIC; 
  signal maccontrol_dout_28_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_28_22_O : STD_LOGIC; 
  signal maccontrol_dout_29_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_29_22_O : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_6_26_SW0_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_6_26_SW0_O_GROM : STD_LOGIC; 
  signal maccontrol_n0067_FROM : STD_LOGIC; 
  signal maccontrol_n0067_GROM : STD_LOGIC; 
  signal maccontrol_n00691_1_FROM : STD_LOGIC; 
  signal maccontrol_n00691_1_GROM : STD_LOGIC; 
  signal maccontrol_n0083_FROM : STD_LOGIC; 
  signal maccontrol_n0083_GROM : STD_LOGIC; 
  signal MD_0_IFF_RST : STD_LOGIC; 
  signal maccontrol_N30192_FROM : STD_LOGIC; 
  signal maccontrol_N30192_GROM : STD_LOGIC; 
  signal maccontrol_n00671_1_FROM : STD_LOGIC; 
  signal maccontrol_n00671_1_GROM : STD_LOGIC; 
  signal memtest2_Ker2265830_O_FROM : STD_LOGIC; 
  signal memtest2_Ker2265830_O_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_9_18_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_9_18_O_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_14_26_SW0_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_14_26_SW0_O_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_8_26_SW0_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_8_26_SW0_O_GROM : STD_LOGIC; 
  signal maccontrol_n0084_FROM : STD_LOGIC; 
  signal maccontrol_n0084_GROM : STD_LOGIC; 
  signal maccontrol_n00701_1_FROM : STD_LOGIC; 
  signal maccontrol_n00701_1_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_1_26_SW0_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_1_26_SW0_O_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_0_11_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_0_11_O_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O_GROM : STD_LOGIC; 
  signal maccontrol_N30311_FROM : STD_LOGIC; 
  signal maccontrol_N30311_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_4_18_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_4_18_O_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_3_6_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_3_6_O_GROM : STD_LOGIC; 
  signal maccontrol_N30199_FROM : STD_LOGIC; 
  signal maccontrol_N30199_GROM : STD_LOGIC; 
  signal maccontrol_N42043_FROM : STD_LOGIC; 
  signal maccontrol_N42043_GROM : STD_LOGIC; 
  signal MD_1_IFF_RST : STD_LOGIC; 
  signal maccontrol_n00397_O_FROM : STD_LOGIC; 
  signal maccontrol_n00397_O_GROM : STD_LOGIC; 
  signal maccontrol_N30181_FROM : STD_LOGIC; 
  signal maccontrol_N30181_GROM : STD_LOGIC; 
  signal maccontrol_n003923_O_FROM : STD_LOGIC; 
  signal maccontrol_n003923_O_GROM : STD_LOGIC; 
  signal maccontrol_N30292_FROM : STD_LOGIC; 
  signal maccontrol_N30292_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_12_18_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_12_18_O_GROM : STD_LOGIC; 
  signal MD_0_OFF_RST : STD_LOGIC; 
  signal maccontrol_N30299_FROM : STD_LOGIC; 
  signal maccontrol_N30299_GROM : STD_LOGIC; 
  signal maccontrol_phyaddr_31_FROM : STD_LOGIC; 
  signal maccontrol_phyaddr_31_GROM : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_4_net55 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_5_net53 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_11_net105 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_6_net51 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_12_net103 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_7_net49 : STD_LOGIC; 
  signal MD_0_TFF_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_8_net47 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd3_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd3_In : STD_LOGIC; 
  signal memtest2_Mshreg_data4_14_net99 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_22_net83 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_30_net67 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd5_In : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd4_In : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_9_net45 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_15_net97 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_23_net81 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_31_net65 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_16_net95 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_17_net93 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_25_net77 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_18_net91 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_26_net75 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_19_net89 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_27_net73 : STD_LOGIC; 
  signal memcontroller_dnl1_1_CEMUXNOT : STD_LOGIC; 
  signal memtest2_Mshreg_data4_28_41_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_28_net71 : STD_LOGIC; 
  signal memcontroller_dnl1_3_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_5_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_5_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_7_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_7_CEMUXNOT : STD_LOGIC; 
  signal TX_EN_OFF_RST : STD_LOGIC; 
  signal memcontroller_dnl1_9_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_9_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_clknum_1_2_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_1_2_GROM : STD_LOGIC; 
  signal MD_1_OFF_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_29_40_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_29_net69 : STD_LOGIC; 
  signal maccontrol_Mshreg_scslll_net281 : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_statecnt_0_FROM : STD_LOGIC; 
  signal memcontroller_dnl1_11_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_21_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_21_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_13_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_13_CEMUXNOT : STD_LOGIC; 
  signal MD_1_TFF_RST : STD_LOGIC; 
  signal memcontroller_dnl1_31_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_31_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_23_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_23_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_15_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_15_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_25_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_25_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_17_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_17_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_27_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_27_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_19_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_19_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl1_29_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_29_CEMUXNOT : STD_LOGIC; 
  signal memtest2_n0214 : STD_LOGIC; 
  signal clken_clkcnt_2_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd2_In : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd1_In : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd4_In : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd3_In : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd6_In : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd5_In : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd8_In : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd7_In : STD_LOGIC; 
  signal memtest2_Mshreg_data4_0_net127 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_1_net125 : STD_LOGIC; 
  signal maccontrol_Mshreg_sinlll_net279 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_10_net43 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_2_net123 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_11_net41 : STD_LOGIC; 
  signal MD_2_IFF_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_3_net121 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_12_net39 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_20_net23 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_4_net119 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_13_net37 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_21_net21 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_5_net117 : STD_LOGIC; 
  signal testrx_cs_FFd2_FROM : STD_LOGIC; 
  signal testrx_cs_FFd2_In : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_14_net35 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_22_net19 : STD_LOGIC; 
  signal testrx_cs_FFd3_FROM : STD_LOGIC; 
  signal testrx_cs_FFd3_In : STD_LOGIC; 
  signal memtest2_Mshreg_data4_6_net115 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_15_net33 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_23_net17 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_7_net113 : STD_LOGIC; 
  signal txsim_Mshreg_TX_EN_net129_LOGIC_ONE : STD_LOGIC; 
  signal txsim_Mshreg_TX_EN_net129_GSHIFT : STD_LOGIC; 
  signal memtest2_n002184_SW0_2_GROM : STD_LOGIC; 
  signal MA_12_OFF_RST : STD_LOGIC; 
  signal maccontrol_din_13_FFY_RST : STD_LOGIC; 
  signal maccontrol_n0022_FROM : STD_LOGIC; 
  signal maccontrol_n0022_GROM : STD_LOGIC; 
  signal MA_13_OFF_RST : STD_LOGIC; 
  signal memcontroller_oel_BYMUXNOT : STD_LOGIC; 
  signal memcontroller_oel_CEMUXNOT : STD_LOGIC; 
  signal maccontrol_Ker303141_1_FROM : STD_LOGIC; 
  signal maccontrol_Ker303141_1_GROM : STD_LOGIC; 
  signal memtest2_deql_0_FROM : STD_LOGIC; 
  signal memtest2_deq_0_rt : STD_LOGIC; 
  signal memtest2_deql_0_CYINIT : STD_LOGIC; 
  signal txsim_N46398_GROM : STD_LOGIC; 
  signal memtest2_deql_2_FROM : STD_LOGIC; 
  signal memtest2_deq_2_rt : STD_LOGIC; 
  signal memtest2_deql_2_CYINIT : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd6_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd6_In : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_11_40_SW0_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_11_40_SW0_O_GROM : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_16_net31 : STD_LOGIC; 
  signal MD_3_IFF_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_24_net15 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_8_net111 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_17_net29 : STD_LOGIC; 
  signal MD_2_OFF_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_25_net13 : STD_LOGIC; 
  signal memtest2_Mshreg_data4_9_net109 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_26_net11 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_18_net27 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_27_net9 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_19_net25 : STD_LOGIC; 
  signal maccontrol_lsclkdelta : STD_LOGIC; 
  signal memcontroller_oe_FROM : STD_LOGIC; 
  signal memcontroller_wen : STD_LOGIC; 
  signal MD_2_TFF_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_30_net3 : STD_LOGIC; 
  signal memtest2_n0150 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_31_6_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_31_net1 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_28_net7 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_29_net5 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_0_net63 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_1_net61 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_2_net59 : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_3_net57 : STD_LOGIC; 
  signal memtest2_datain_13_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_21_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_15_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_23_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_31_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_25_FFY_RST : STD_LOGIC; 
  signal d2_11_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_26_FFY_RST : STD_LOGIC; 
  signal MD_4_IFF_RST : STD_LOGIC; 
  signal MD_3_OFF_RST : STD_LOGIC; 
  signal err_FFY_RST : STD_LOGIC; 
  signal MD_3_TFF_RST : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_8_26_2_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_8_26_2_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N46670_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N46670_GROM : STD_LOGIC; 
  signal maccontrol_phydo_5_FFY_RST : STD_LOGIC; 
  signal MDC_OBUF_FFY_RST : STD_LOGIC; 
  signal addr4_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydo_9_FFY_RST : STD_LOGIC; 
  signal addr4_3_FFY_RST : STD_LOGIC; 
  signal addr4_7_FFY_RST : STD_LOGIC; 
  signal addr4_9_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_1_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_6_26_2_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_6_26_2_GROM : STD_LOGIC; 
  signal MD_5_IFF_RST : STD_LOGIC; 
  signal memtest2_ldata_7_FFY_RST : STD_LOGIC; 
  signal MD_4_OFF_RST : STD_LOGIC; 
  signal q2_3_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_9_FFY_RST : STD_LOGIC; 
  signal q2_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_N30285_FROM : STD_LOGIC; 
  signal maccontrol_N30285_GROM : STD_LOGIC; 
  signal maccontrol_N30273_FROM : STD_LOGIC; 
  signal maccontrol_N30273_GROM : STD_LOGIC; 
  signal MD_4_TFF_RST : STD_LOGIC; 
  signal q4_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_7_40_SW0_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_7_40_SW0_O_GROM : STD_LOGIC; 
  signal maccontrol_N30212_FROM : STD_LOGIC; 
  signal maccontrol_N30212_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_n00151_1_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_n00151_1_GROM : STD_LOGIC; 
  signal memtest2_CHOICE1064_GROM : STD_LOGIC; 
  signal memtest2_CHOICE1067_FROM : STD_LOGIC; 
  signal memtest2_CHOICE1067_GROM : STD_LOGIC; 
  signal maccontrol_phyaddr_2_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_9_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_9_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydo_11_FFY_RST : STD_LOGIC; 
  signal MD_5_OFF_RST : STD_LOGIC; 
  signal maccontrol_phydo_13_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydo_15_FFY_RST : STD_LOGIC; 
  signal addr4_11_FFY_RST : STD_LOGIC; 
  signal addr4_13_FFY_RST : STD_LOGIC; 
  signal addr4_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_10_26_2_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_10_26_2_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE920_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE920_GROM : STD_LOGIC; 
  signal MD_5_TFF_RST : STD_LOGIC; 
  signal Q_n0034_2_FROM : STD_LOGIC; 
  signal Q_n0034_2_GROM : STD_LOGIC; 
  signal MD_6_IFF_RST : STD_LOGIC; 
  signal memcontroller_dnl2_1_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_1_CEMUXNOT : STD_LOGIC; 
  signal maccontrol_lmacaddr_11_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_3_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_3_CEMUXNOT : STD_LOGIC; 
  signal maccontrol_lmacaddr_13_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_5_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_5_CEMUXNOT : STD_LOGIC; 
  signal maccontrol_lmacaddr_15_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_11_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_7_CEMUXNOT : STD_LOGIC; 
  signal MD_6_OFF_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_41_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_17_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_25_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_0_2_BXMUXNOT : STD_LOGIC; 
  signal memcontroller_clknum_0_2_BYMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_9_CEMUXNOT : STD_LOGIC; 
  signal MD_6_TFF_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_19_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_31_FFY_RST : STD_LOGIC; 
  signal MD_7_IFF_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_29_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_47_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_27_FFY_RST : STD_LOGIC; 
  signal MD_8_IFF_RST : STD_LOGIC; 
  signal MD_7_OFF_RST : STD_LOGIC; 
  signal memtest2_lfsr_rst_FROM : STD_LOGIC; 
  signal memtest2_n0021 : STD_LOGIC; 
  signal MD_7_TFF_RST : STD_LOGIC; 
  signal testrx_CHOICE930_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE735_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE735_GROM : STD_LOGIC; 
  signal testrx_CHOICE933_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1204_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1204_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1543_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1543_GROM : STD_LOGIC; 
  signal maccontrol_n0032_FROM : STD_LOGIC; 
  signal maccontrol_n0032_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1489_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1489_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1546_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1546_GROM : STD_LOGIC; 
  signal maccontrol_N46676_FROM : STD_LOGIC; 
  signal maccontrol_N46676_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1528_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1528_GROM : STD_LOGIC; 
  signal memtest2_CHOICE948_FROM : STD_LOGIC; 
  signal memtest2_CHOICE948_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1385_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1385_GROM : STD_LOGIC; 
  signal MD_8_OFF_RST : STD_LOGIC; 
  signal maccontrol_CHOICE1443_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1443_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1323_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1323_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1326_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1326_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_miiaddr_1_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_miiaddr_1_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_miiaddr_2_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_miiaddr_2_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_miiaddr_4_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_miiaddr_4_GROM : STD_LOGIC; 
  signal MD_8_TFF_RST : STD_LOGIC; 
  signal maccontrol_sclkll_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_25_FFY_RST : STD_LOGIC; 
  signal MD_9_IFF_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_19_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_29_FFY_RST : STD_LOGIC; 
  signal maccontrol_CHOICE1585_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1585_GROM : STD_LOGIC; 
  signal txsim_llltx_FROM : STD_LOGIC; 
  signal txsim_n0002 : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_15_40_SW0_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_15_40_SW0_O_GROM : STD_LOGIC; 
  signal memtest_llerr_BXMUXNOT : STD_LOGIC; 
  signal memtest2_cs_0_BYMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_11_CEMUXNOT : STD_LOGIC; 
  signal MD_9_OFF_RST : STD_LOGIC; 
  signal memcontroller_dnl2_21_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_13_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_31_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_23_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_15_CEMUXNOT : STD_LOGIC; 
  signal MD_9_TFF_RST : STD_LOGIC; 
  signal memcontroller_dnl2_25_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_17_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_27_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_19_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_29_CEMUXNOT : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N20226_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N20226_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N20221_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N20221_GROM : STD_LOGIC; 
  signal LEDACT_OFF_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N41816_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N41816_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE749_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE749_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE751_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE751_GROM : STD_LOGIC; 
  signal maccontrol_phydi_13_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_23_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_25_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_19_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_27_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_29_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_3_FFY_RST : STD_LOGIC; 
  signal testrx_cs_FFd1_FROM : STD_LOGIC; 
  signal testrx_cs_FFd1_In : STD_LOGIC; 
  signal maccontrol_N46681_FROM : STD_LOGIC; 
  signal maccontrol_N46681_GROM : STD_LOGIC; 
  signal LEDDPX_OFF_RST : STD_LOGIC; 
  signal txsim_N41883_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1561_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1561_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1111_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1111_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_din_11_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_13_FFY_RST : STD_LOGIC; 
  signal maccontrol_CHOICE1234_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1234_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1355_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1355_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1174_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1174_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1147_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1147_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1223_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1223_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_10_26_SW0_O_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_10_26_SW0_O_GROM : STD_LOGIC; 
  signal memtest2_Mshreg_data4_13_net101_GSHIFT : STD_LOGIC; 
  signal memtest2_Mshreg_data4_21_net85_GSHIFT : STD_LOGIC; 
  signal maccontrol_CHOICE1256_GROM : STD_LOGIC; 
  signal maccontrol_n0036_FROM : STD_LOGIC; 
  signal maccontrol_n0036_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1156_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1156_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1389_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1389_GROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_14_26_2_FROM : STD_LOGIC; 
  signal maccontrol_Mmux_n0023_Result_14_26_2_GROM : STD_LOGIC; 
  signal maccontrol_N46402_FROM : STD_LOGIC; 
  signal maccontrol_N46402_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1410_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1410_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE802_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE802_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE812_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE812_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE829_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE829_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1319_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1319_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1368_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_N23512_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_N23512_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1240_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1240_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_N23520_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_N23520_GROM : STD_LOGIC; 
  signal MA_10_OFF_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_n0013_GROM : STD_LOGIC; 
  signal clken_clkcnt_0_BXMUXNOT : STD_LOGIC; 
  signal clken_clkcnt_0_FROM : STD_LOGIC; 
  signal maccontrol_n001223_1_FROM : STD_LOGIC; 
  signal maccontrol_n001223_1_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE729_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_CHOICE729_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1338_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1338_GROM : STD_LOGIC; 
  signal MA_11_OFF_RST : STD_LOGIC; 
  signal maccontrol_CHOICE1262_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1262_GROM : STD_LOGIC; 
  signal memtest2_N41527_FROM : STD_LOGIC; 
  signal memtest2_N41527_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_N42089_GROM : STD_LOGIC; 
  signal txsim_CHOICE1098_GROM : STD_LOGIC; 
  signal txsim_CHOICE1090_FROM : STD_LOGIC; 
  signal txsim_CHOICE1090_GROM : STD_LOGIC; 
  signal txsim_CHOICE1105_GROM : STD_LOGIC; 
  signal d2_0_FFY_RST : STD_LOGIC; 
  signal d2_0_FFX_RST : STD_LOGIC; 
  signal d2_3_FFY_RST : STD_LOGIC; 
  signal d2_3_FFX_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_13_56_FFX_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_21_48_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd6_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd8_FFX_SET : STD_LOGIC; 
  signal memtest2_Mshreg_data4_0_69_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_1_68_FFY_RST : STD_LOGIC; 
  signal maccontrol_Mshreg_sinlll_83_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_10_27_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_3_66_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_2_67_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_11_26_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_12_25_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_19_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_29_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd4_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_phyaddrws_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_12_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_20_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_21_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_22_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_13_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_30_FFY_RST : STD_LOGIC; 
  signal MA_14_OFF_RST : STD_LOGIC; 
  signal maccontrol_n00131_1_FROM : STD_LOGIC; 
  signal maccontrol_n00131_1_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1033_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N46538_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_N46538_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1041_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1050_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1050_GROM : STD_LOGIC; 
  signal maccontrol_N30206_FROM : STD_LOGIC; 
  signal maccontrol_N30206_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1048_GROM : STD_LOGIC; 
  signal maccontrol_N30305_FROM : STD_LOGIC; 
  signal maccontrol_N30305_GROM : STD_LOGIC; 
  signal maccontrol_N30228_FROM : STD_LOGIC; 
  signal maccontrol_N30228_GROM : STD_LOGIC; 
  signal MA_15_OFF_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_4_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_6_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_8_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_8_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_10_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_10_FFY_RST : STD_LOGIC; 
  signal memtest_addrcntl_11_FFX_RST : STD_LOGIC; 
  signal memtest_addrcntl_11_FFY_RST : STD_LOGIC; 
  signal memtest_addrcntl_13_FFX_RST : STD_LOGIC; 
  signal memtest_addrcntl_13_FFY_RST : STD_LOGIC; 
  signal maccontrol_CHOICE1002_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1002_GROM : STD_LOGIC; 
  signal memtest_addrcntl_15_FFX_RST : STD_LOGIC; 
  signal memtest_addrcntl_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_CHOICE1608_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1608_GROM : STD_LOGIC; 
  signal clken1_FROM : STD_LOGIC; 
  signal clken1_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_11_FFY_RST : STD_LOGIC; 
  signal maccontrol_n0011_FROM : STD_LOGIC; 
  signal maccontrol_n0011_GROM : STD_LOGIC; 
  signal maccontrol_n003963_O_FROM : STD_LOGIC; 
  signal maccontrol_n003963_O_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_miirw_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_miirw_GROM : STD_LOGIC; 
  signal memcontroller_n0007_FROM : STD_LOGIC; 
  signal memcontroller_n0007_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1017_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1017_GROM : STD_LOGIC; 
  signal MA_16_OFF_RST : STD_LOGIC; 
  signal maccontrol_n00311_1_FROM : STD_LOGIC; 
  signal maccontrol_n00311_1_GROM : STD_LOGIC; 
  signal SOUT_OFF_RST : STD_LOGIC; 
  signal maccontrol_n0043_FROM : STD_LOGIC; 
  signal maccontrol_n0043_GROM : STD_LOGIC; 
  signal maccontrol_n0037_FROM : STD_LOGIC; 
  signal maccontrol_n0037_GROM : STD_LOGIC; 
  signal maccontrol_newcmd_FROM : STD_LOGIC; 
  signal maccontrol_newcmd_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE974_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1055_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE1055_GROM : STD_LOGIC; 
  signal MACDATA_0_OFF_RST : STD_LOGIC; 
  signal maccontrol_CHOICE1596_GROM : STD_LOGIC; 
  signal maccontrol_n0070_FROM : STD_LOGIC; 
  signal maccontrol_n0070_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE981_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE981_GROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd2_FROM : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd2_In : STD_LOGIC; 
  signal maccontrol_CHOICE988_FROM : STD_LOGIC; 
  signal maccontrol_CHOICE988_GROM : STD_LOGIC; 
  signal maccontrol_n0234_GROM : STD_LOGIC; 
  signal maccontrol_CHOICE1603_GROM : STD_LOGIC; 
  signal maccontrol_n0068_GROM : STD_LOGIC; 
  signal memtest2_laddr_3_FFY_RST : STD_LOGIC; 
  signal memtest2_n0117_FROM : STD_LOGIC; 
  signal memtest2_n0117_GROM : STD_LOGIC; 
  signal memtest2_laddr_5_FFY_RST : STD_LOGIC; 
  signal memtest2_laddr_13_FFY_RST : STD_LOGIC; 
  signal memtest2_laddr_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_statecnt_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_statecnt_1_FROM : STD_LOGIC; 
  signal memtest2_CHOICE941_GROM : STD_LOGIC; 
  signal MACDATA_1_OFF_RST : STD_LOGIC; 
  signal LEDRX_N1683_GROM : STD_LOGIC; 
  signal memtest2_n0119_GROM : STD_LOGIC; 
  signal memcontroller_clknum_1_BYMUXNOT : STD_LOGIC; 
  signal maccontrol_N46368_FROM : STD_LOGIC; 
  signal maccontrol_N46368_GROM : STD_LOGIC; 
  signal clken_lclken_LOGIC_ONE : STD_LOGIC; 
  signal MACDATA_2_OFF_RST : STD_LOGIC; 
  signal MACDATA_3_OFF_RST : STD_LOGIC; 
  signal MACDATA_4_OFF_RST : STD_LOGIC; 
  signal MACDATA_5_OFF_RST : STD_LOGIC; 
  signal MACDATA_6_OFF_RST : STD_LOGIC; 
  signal MACDATA_7_OFF_RST : STD_LOGIC; 
  signal MACDATA_8_OFF_RST : STD_LOGIC; 
  signal MD_10_IFF_RST : STD_LOGIC; 
  signal MD_31_TFF_RST : STD_LOGIC; 
  signal MD_24_OFF_RST : STD_LOGIC; 
  signal MD_24_TFF_RST : STD_LOGIC; 
  signal MD_16_IFF_RST : STD_LOGIC; 
  signal MD_16_OFF_RST : STD_LOGIC; 
  signal MD_16_TFF_RST : STD_LOGIC; 
  signal MD_17_IFF_RST : STD_LOGIC; 
  signal MD_25_IFF_RST : STD_LOGIC; 
  signal MD_17_OFF_RST : STD_LOGIC; 
  signal MD_10_OFF_RST : STD_LOGIC; 
  signal MD_10_TFF_RST : STD_LOGIC; 
  signal MACDATA_9_OFF_RST : STD_LOGIC; 
  signal MD_11_IFF_RST : STD_LOGIC; 
  signal MD_11_OFF_RST : STD_LOGIC; 
  signal MD_11_TFF_RST : STD_LOGIC; 
  signal MD_20_IFF_RST : STD_LOGIC; 
  signal MD_12_IFF_RST : STD_LOGIC; 
  signal MD_20_OFF_RST : STD_LOGIC; 
  signal MDIO_IFF_RST : STD_LOGIC; 
  signal RXD_0_IFF_RST : STD_LOGIC; 
  signal RXD_1_IFF_RST : STD_LOGIC; 
  signal RXD_2_IFF_RST : STD_LOGIC; 
  signal RXD_3_IFF_RST : STD_LOGIC; 
  signal RXD_4_IFF_RST : STD_LOGIC; 
  signal RXD_5_IFF_RST : STD_LOGIC; 
  signal MD_28_OFF_RST : STD_LOGIC; 
  signal MD_28_TFF_RST : STD_LOGIC; 
  signal MD_29_IFF_RST : STD_LOGIC; 
  signal MD_29_OFF_RST : STD_LOGIC; 
  signal MD_29_TFF_RST : STD_LOGIC; 
  signal LED100_OFF_RST : STD_LOGIC; 
  signal NEXTF_IFF_RST : STD_LOGIC; 
  signal MD_30_TFF_RST : STD_LOGIC; 
  signal MD_23_OFF_RST : STD_LOGIC; 
  signal MD_23_TFF_RST : STD_LOGIC; 
  signal MD_15_IFF_RST : STD_LOGIC; 
  signal MD_15_OFF_RST : STD_LOGIC; 
  signal MD_15_TFF_RST : STD_LOGIC; 
  signal MD_31_IFF_RST : STD_LOGIC; 
  signal MD_24_IFF_RST : STD_LOGIC; 
  signal MD_31_OFF_RST : STD_LOGIC; 
  signal MWE_OFF_SET : STD_LOGIC; 
  signal RXD_6_IFF_RST : STD_LOGIC; 
  signal RXD_7_IFF_RST : STD_LOGIC; 
  signal LED1000_OFF_RST : STD_LOGIC; 
  signal RX_DV_IFF_RST : STD_LOGIC; 
  signal MACDATA_10_OFF_RST : STD_LOGIC; 
  signal d1_0_FFY_RST : STD_LOGIC; 
  signal d1_2_FFY_RST : STD_LOGIC; 
  signal d1_0_FFX_RST : STD_LOGIC; 
  signal d1_4_FFY_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_123_FFY_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_125_FFY_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_127_FFY_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_123_FFX_RST : STD_LOGIC; 
  signal MACDATA_11_OFF_RST : STD_LOGIC; 
  signal MACDATA_12_OFF_RST : STD_LOGIC; 
  signal MACDATA_13_OFF_RST : STD_LOGIC; 
  signal MACDATA_14_OFF_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_125_FFX_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_127_FFX_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_129_FFY_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_129_FFX_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_131_FFY_RST : STD_LOGIC; 
  signal maccontrol_bitcnt_86_FFX_RST : STD_LOGIC; 
  signal maccontrol_bitcnt_88_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_91_FFY_RST : STD_LOGIC; 
  signal maccontrol_bitcnt_90_FFX_RST : STD_LOGIC; 
  signal maccontrol_bitcnt_88_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_92_FFY_RST : STD_LOGIC; 
  signal MD_26_TFF_RST : STD_LOGIC; 
  signal MD_19_OFF_RST : STD_LOGIC; 
  signal MD_19_TFF_RST : STD_LOGIC; 
  signal MD_27_IFF_RST : STD_LOGIC; 
  signal MD_27_OFF_RST : STD_LOGIC; 
  signal MD_27_TFF_RST : STD_LOGIC; 
  signal PHYRESET_OFF_RST : STD_LOGIC; 
  signal MD_28_IFF_RST : STD_LOGIC; 
  signal MD_13_TFF_RST : STD_LOGIC; 
  signal MD_22_OFF_RST : STD_LOGIC; 
  signal MD_22_TFF_RST : STD_LOGIC; 
  signal MD_14_IFF_RST : STD_LOGIC; 
  signal MD_14_OFF_RST : STD_LOGIC; 
  signal MD_14_TFF_RST : STD_LOGIC; 
  signal MD_30_IFF_RST : STD_LOGIC; 
  signal MD_23_IFF_RST : STD_LOGIC; 
  signal MD_30_OFF_RST : STD_LOGIC; 
  signal cnt_2_FFX_RST : STD_LOGIC; 
  signal cnt_4_FFY_RST : STD_LOGIC; 
  signal cnt_8_FFY_RST : STD_LOGIC; 
  signal cnt_4_FFX_RST : STD_LOGIC; 
  signal cnt_6_FFY_RST : STD_LOGIC; 
  signal MD_20_TFF_RST : STD_LOGIC; 
  signal MD_12_OFF_RST : STD_LOGIC; 
  signal MD_12_TFF_RST : STD_LOGIC; 
  signal MD_21_IFF_RST : STD_LOGIC; 
  signal MD_21_OFF_RST : STD_LOGIC; 
  signal MD_21_TFF_RST : STD_LOGIC; 
  signal MD_13_IFF_RST : STD_LOGIC; 
  signal MD_22_IFF_RST : STD_LOGIC; 
  signal MD_13_OFF_RST : STD_LOGIC; 
  signal cnt_6_FFX_RST : STD_LOGIC; 
  signal cnt_8_FFX_RST : STD_LOGIC; 
  signal cnt_10_FFY_RST : STD_LOGIC; 
  signal cnt_14_FFY_RST : STD_LOGIC; 
  signal cnt_10_FFX_RST : STD_LOGIC; 
  signal cnt_12_FFY_RST : STD_LOGIC; 
  signal MD_17_TFF_RST : STD_LOGIC; 
  signal MD_25_OFF_RST : STD_LOGIC; 
  signal MD_25_TFF_RST : STD_LOGIC; 
  signal MD_18_IFF_RST : STD_LOGIC; 
  signal MD_18_OFF_RST : STD_LOGIC; 
  signal MD_18_TFF_RST : STD_LOGIC; 
  signal MD_26_IFF_RST : STD_LOGIC; 
  signal MD_19_IFF_RST : STD_LOGIC; 
  signal MD_26_OFF_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_110_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_112_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_116_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_112_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_114_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_114_FFX_RST : STD_LOGIC; 
  signal MACDATA_15_OFF_RST : STD_LOGIC; 
  signal LEDTX_OFF_RST : STD_LOGIC; 
  signal LEDPOWER_OFF_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_96_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_98_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_100_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_102_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_100_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_104_FFY_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_131_FFX_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_133_FFY_RST : STD_LOGIC; 
  signal maccontrol_bitcnt_86_FFY_RST : STD_LOGIC; 
  signal maccontrol_ledtx_cnt_133_FFX_RST : STD_LOGIC; 
  signal maccontrol_bitcnt_85_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_27_10_FFY_RST : STD_LOGIC; 
  signal memcontroller_oe_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_19_18_FFY_RST : STD_LOGIC; 
  signal maccontrol_sclkdelta_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_30_7_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_0_37_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_28_9_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_29_8_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_92_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_94_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_94_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_96_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_98_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_102_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_104_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_106_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_106_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_108_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_108_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_110_FFY_RST : STD_LOGIC; 
  signal cnt_0_FFY_RST : STD_LOGIC; 
  signal cnt_0_FFX_RST : STD_LOGIC; 
  signal cnt_2_FFY_RST : STD_LOGIC; 
  signal cnt_12_FFX_RST : STD_LOGIC; 
  signal cnt_14_FFX_RST : STD_LOGIC; 
  signal cnt_16_FFY_RST : STD_LOGIC; 
  signal cnt_16_FFX_RST : STD_LOGIC; 
  signal cnt_18_FFY_RST : STD_LOGIC; 
  signal d1_8_FFX_RST : STD_LOGIC; 
  signal d1_10_FFX_RST : STD_LOGIC; 
  signal d1_12_FFY_RST : STD_LOGIC; 
  signal d1_12_FFX_RST : STD_LOGIC; 
  signal d1_14_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_120_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_122_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_116_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_118_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_118_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyrstcnt_120_FFY_RST : STD_LOGIC; 
  signal d1_18_FFX_RST : STD_LOGIC; 
  signal d1_20_FFX_RST : STD_LOGIC; 
  signal d1_22_FFY_RST : STD_LOGIC; 
  signal d1_26_FFY_RST : STD_LOGIC; 
  signal d1_22_FFX_RST : STD_LOGIC; 
  signal d1_24_FFY_RST : STD_LOGIC; 
  signal d1_2_FFX_RST : STD_LOGIC; 
  signal d1_4_FFX_RST : STD_LOGIC; 
  signal d1_6_FFY_RST : STD_LOGIC; 
  signal d1_10_FFY_RST : STD_LOGIC; 
  signal d1_6_FFX_RST : STD_LOGIC; 
  signal d1_8_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_3_FFY_RST : STD_LOGIC; 
  signal cnt_18_FFX_RST : STD_LOGIC; 
  signal cnt_20_FFY_RST : STD_LOGIC; 
  signal cnt_20_FFX_RST : STD_LOGIC; 
  signal cnt_22_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_mdccnt_0_FFY_RST : STD_LOGIC; 
  signal cnt_22_FFX_RST : STD_LOGIC; 
  signal d1_14_FFX_RST : STD_LOGIC; 
  signal d1_16_FFY_RST : STD_LOGIC; 
  signal d1_20_FFY_RST : STD_LOGIC; 
  signal d1_16_FFX_RST : STD_LOGIC; 
  signal d1_18_FFY_RST : STD_LOGIC; 
  signal d1_30_FFX_RST : STD_LOGIC; 
  signal addr1_0_FFY_RST : STD_LOGIC; 
  signal addr1_4_FFY_RST : STD_LOGIC; 
  signal addr1_0_FFX_RST : STD_LOGIC; 
  signal addr1_2_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_14_FFX_RST : STD_LOGIC; 
  signal maccontrol_dout_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_8_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_8_FFX_RST : STD_LOGIC; 
  signal addr1_8_FFX_RST : STD_LOGIC; 
  signal addr1_10_FFX_RST : STD_LOGIC; 
  signal addr1_12_FFY_RST : STD_LOGIC; 
  signal addr1_12_FFX_RST : STD_LOGIC; 
  signal addr1_14_FFY_RST : STD_LOGIC; 
  signal addr1_14_FFX_RST : STD_LOGIC; 
  signal addr2_13_FFY_RST : STD_LOGIC; 
  signal addr2_13_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_11_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_30_FFX_RST : STD_LOGIC; 
  signal maccontrol_dout_0_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_26_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_27_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_19_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_28_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_29_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_27_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_31_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_23_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_23_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_15_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_15_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_37_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_37_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_45_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_45_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_29_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_25_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_25_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_17_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_39_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_30_39_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd5_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd5_FFX_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_9_28_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_15_54_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_23_46_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_31_38_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_16_53_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_18_51_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_17_52_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_25_44_FFY_RST : STD_LOGIC; 
  signal d1_24_FFX_RST : STD_LOGIC; 
  signal d1_30_FFY_RST : STD_LOGIC; 
  signal d1_26_FFX_RST : STD_LOGIC; 
  signal d1_28_FFY_RST : STD_LOGIC; 
  signal d1_28_FFX_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_1_36_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_2_35_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_3_34_FFY_RST : STD_LOGIC; 
  signal addr2_15_FFY_RST : STD_LOGIC; 
  signal addr2_15_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_13_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_21_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_15_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_23_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_17_FFY_RST : STD_LOGIC; 
  signal addr1_2_FFX_RST : STD_LOGIC; 
  signal addr1_4_FFX_RST : STD_LOGIC; 
  signal addr1_6_FFY_RST : STD_LOGIC; 
  signal addr1_10_FFY_RST : STD_LOGIC; 
  signal addr1_6_FFX_RST : STD_LOGIC; 
  signal addr1_8_FFY_RST : STD_LOGIC; 
  signal memtest2_deql_2_FFY_RST : STD_LOGIC; 
  signal memtest2_deql_2_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd6_FFY_SET : STD_LOGIC; 
  signal maccontrol_din_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_lrxmcast_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_23_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_31_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_24_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_16_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_18_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_17_FFY_RST : STD_LOGIC; 
  signal maccontrol_dout_25_FFY_RST : STD_LOGIC; 
  signal q2_29_FFX_RST : STD_LOGIC; 
  signal q4_11_FFY_RST : STD_LOGIC; 
  signal q4_11_FFX_RST : STD_LOGIC; 
  signal q4_21_FFY_RST : STD_LOGIC; 
  signal q4_21_FFX_RST : STD_LOGIC; 
  signal q4_13_FFY_RST : STD_LOGIC; 
  signal q4_13_FFX_RST : STD_LOGIC; 
  signal q4_31_FFY_RST : STD_LOGIC; 
  signal q4_31_FFX_RST : STD_LOGIC; 
  signal q4_23_FFY_RST : STD_LOGIC; 
  signal q4_23_FFX_RST : STD_LOGIC; 
  signal q4_15_FFY_RST : STD_LOGIC; 
  signal q4_15_FFX_RST : STD_LOGIC; 
  signal q4_25_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_26_43_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_19_50_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_27_42_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_1_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_1_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_3_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_3_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_5_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_7_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_9_FFX_RST : STD_LOGIC; 
  signal memcontroller_clknum_1_2_FFX_RST : STD_LOGIC; 
  signal maccontrol_Mshreg_scslll_84_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_statecnt_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_statecnt_0_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_statecnt_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_statecnt_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_statecnt_5_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_11_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_11_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_21_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_13_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_31_FFX_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_4_33_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_31_FFX_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_5_32_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_11_58_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_6_31_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_12_57_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_7_30_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_8_29_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd3_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_14_55_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_22_47_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_5_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_23_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_15_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_25_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_17_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_27_FFX_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_20_17_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_4_65_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_13_24_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_21_16_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_5_64_FFY_RST : STD_LOGIC; 
  signal testrx_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_14_23_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_22_15_FFY_RST : STD_LOGIC; 
  signal testrx_cs_FFd3_FFY_SET : STD_LOGIC; 
  signal memtest2_Mshreg_data4_6_63_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydo_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydo_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydo_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydo_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydo_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydo_7_FFX_RST : STD_LOGIC; 
  signal addr4_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydo_9_FFX_RST : STD_LOGIC; 
  signal addr4_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_11_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_13_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_21_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_21_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_15_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_23_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_23_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_31_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_31_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_9_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_17_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_9_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_17_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_25_FFX_RST : STD_LOGIC; 
  signal d2_11_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_19_FFY_RST : STD_LOGIC; 
  signal d2_13_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_19_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_27_FFY_RST : STD_LOGIC; 
  signal d2_21_FFY_RST : STD_LOGIC; 
  signal d2_13_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_29_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_29_FFX_RST : STD_LOGIC; 
  signal d2_31_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_15_22_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_23_14_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_7_62_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_16_21_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_24_13_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_8_61_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_17_20_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_25_12_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_18_19_FFY_RST : STD_LOGIC; 
  signal memtest2_Mshreg_data4_9_60_FFY_RST : STD_LOGIC; 
  signal memtest_Mshreg_dataw4_26_11_FFY_RST : STD_LOGIC; 
  signal q4_1_FFX_RST : STD_LOGIC; 
  signal q4_3_FFY_RST : STD_LOGIC; 
  signal q4_3_FFX_RST : STD_LOGIC; 
  signal q4_5_FFY_RST : STD_LOGIC; 
  signal q4_5_FFX_RST : STD_LOGIC; 
  signal q4_7_FFY_RST : STD_LOGIC; 
  signal q4_7_FFX_RST : STD_LOGIC; 
  signal q4_9_FFY_RST : STD_LOGIC; 
  signal q4_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_1_FFY_RST : STD_LOGIC; 
  signal d2_31_FFX_RST : STD_LOGIC; 
  signal d2_22_FFY_RST : STD_LOGIC; 
  signal d2_15_FFY_RST : STD_LOGIC; 
  signal d2_15_FFX_RST : STD_LOGIC; 
  signal d2_25_FFY_RST : STD_LOGIC; 
  signal d2_25_FFX_RST : STD_LOGIC; 
  signal d2_17_FFY_RST : STD_LOGIC; 
  signal d2_17_FFX_RST : STD_LOGIC; 
  signal d2_27_FFY_RST : STD_LOGIC; 
  signal d2_27_FFX_RST : STD_LOGIC; 
  signal d2_19_FFY_RST : STD_LOGIC; 
  signal d2_19_FFX_RST : STD_LOGIC; 
  signal d2_29_FFY_RST : STD_LOGIC; 
  signal d2_29_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydo_1_FFY_RST : STD_LOGIC; 
  signal q4_25_FFX_RST : STD_LOGIC; 
  signal q4_17_FFY_RST : STD_LOGIC; 
  signal q4_17_FFX_RST : STD_LOGIC; 
  signal q4_27_FFY_RST : STD_LOGIC; 
  signal q4_27_FFX_RST : STD_LOGIC; 
  signal q4_19_FFY_RST : STD_LOGIC; 
  signal q4_19_FFX_RST : STD_LOGIC; 
  signal q4_29_FFY_RST : STD_LOGIC; 
  signal q4_29_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_7_FFX_RST : STD_LOGIC; 
  signal q2_3_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_9_FFX_RST : STD_LOGIC; 
  signal q2_5_FFX_RST : STD_LOGIC; 
  signal q2_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_done_FFY_RST : STD_LOGIC; 
  signal q2_7_FFX_RST : STD_LOGIC; 
  signal q2_9_FFY_RST : STD_LOGIC; 
  signal q2_9_FFX_RST : STD_LOGIC; 
  signal addr4_3_FFX_RST : STD_LOGIC; 
  signal addr4_5_FFX_RST : STD_LOGIC; 
  signal addr4_7_FFX_RST : STD_LOGIC; 
  signal addr4_9_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_1_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_3_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_3_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_5_FFX_RST : STD_LOGIC; 
  signal q2_1_FFY_RST : STD_LOGIC; 
  signal q2_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_13_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_21_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_21_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_15_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_30_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_22_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_23_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_17_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_17_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_25_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_27_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_19_FFX_RST : STD_LOGIC; 
  signal testrx_rxdll_7_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_11_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_11_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_11_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_11_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_21_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_21_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_13_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_13_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_21_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_21_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_13_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_13_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_31_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_27_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_29_FFX_RST : STD_LOGIC; 
  signal txsim_llltx_FFY_RST : STD_LOGIC; 
  signal memtest_llerr_FFX_RST : STD_LOGIC; 
  signal testrx_rxdll_1_FFY_RST : STD_LOGIC; 
  signal testrx_rxdll_1_FFX_RST : STD_LOGIC; 
  signal testrx_rxdll_3_FFY_RST : STD_LOGIC; 
  signal testrx_rxdll_5_FFY_RST : STD_LOGIC; 
  signal testrx_rxdll_3_FFX_RST : STD_LOGIC; 
  signal memtest2_cs_0_FFY_SET : STD_LOGIC; 
  signal testrx_rxdll_7_FFY_RST : STD_LOGIC; 
  signal testrx_rxdll_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydo_11_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydo_13_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydo_15_FFX_RST : STD_LOGIC; 
  signal addr4_11_FFX_RST : STD_LOGIC; 
  signal addr4_13_FFX_RST : STD_LOGIC; 
  signal addr4_15_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_23_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_31_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_15_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_11_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_7_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_33_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_33_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_41_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_17_FFX_RST : STD_LOGIC; 
  signal memcontroller_clknum_0_2_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_11_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_21_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_21_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_13_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_23_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_31_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_25_FFX_RST : STD_LOGIC; 
  signal memcontroller_clknum_0_2_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_21_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_21_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_13_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_13_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_9_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_35_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_35_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_43_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_43_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_19_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_27_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_17_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_39_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_47_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_27_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_19_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_19_FFX_RST : STD_LOGIC; 
  signal memtest2_ldata_29_FFY_RST : STD_LOGIC; 
  signal memtest2_ldata_29_FFX_RST : STD_LOGIC; 
  signal q2_11_FFY_RST : STD_LOGIC; 
  signal q2_11_FFX_RST : STD_LOGIC; 
  signal q2_21_FFY_RST : STD_LOGIC; 
  signal q2_21_FFX_RST : STD_LOGIC; 
  signal q2_13_FFY_RST : STD_LOGIC; 
  signal q2_31_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_11_FFY_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_11_FFX_RST : STD_LOGIC; 
  signal maccontrol_phyaddr_13_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_29_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_11_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_11_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_13_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_21_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_21_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_22_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_15_FFX_RST : STD_LOGIC; 
  signal q2_13_FFX_RST : STD_LOGIC; 
  signal q2_31_FFX_RST : STD_LOGIC; 
  signal q2_23_FFY_RST : STD_LOGIC; 
  signal q2_23_FFX_RST : STD_LOGIC; 
  signal q2_15_FFY_RST : STD_LOGIC; 
  signal q2_15_FFX_RST : STD_LOGIC; 
  signal q2_25_FFY_RST : STD_LOGIC; 
  signal q2_25_FFX_RST : STD_LOGIC; 
  signal q2_17_FFY_RST : STD_LOGIC; 
  signal q2_17_FFX_RST : STD_LOGIC; 
  signal memtest2_lfsr_rst_FFY_RST : STD_LOGIC; 
  signal q2_27_FFX_RST : STD_LOGIC; 
  signal q2_27_FFY_RST : STD_LOGIC; 
  signal q2_19_FFY_RST : STD_LOGIC; 
  signal q2_29_FFY_RST : STD_LOGIC; 
  signal q2_19_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_31_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_23_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_23_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_15_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_15_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_31_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_31_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_23_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_23_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_15_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_15_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_25_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_25_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_17_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_25_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_17_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_9_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_sclkdeltall_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_addrl_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_31_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_31_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_17_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_17_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_25_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_19_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_27_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_29_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_1_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_25_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_17_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_17_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_27_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_27_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_19_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_19_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_27_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_27_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_19_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_19_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_29_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_29_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_29_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_9_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_9_FFX_RST : STD_LOGIC; 
  signal testrx_cs_FFd1_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_12_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_1_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_1_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_2_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_3_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_5_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_5_FFX_RST : STD_LOGIC; 
  signal memtest2_datain_7_FFY_RST : STD_LOGIC; 
  signal memtest2_datain_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_17_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_25_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_25_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_19_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_19_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_27_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_27_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_29_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_29_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_14_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_12_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_11_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_14_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_13_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_15_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_addrl_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_addrl_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_addrl_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_addrl_4_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_9_FFY_RST : STD_LOGIC; 
  signal maccontrol_lmacaddr_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_addr_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_addr_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_addr_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_addr_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_addr_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_addr_5_FFX_RST : STD_LOGIC; 
  signal memtest_lerr_FFY_RST : STD_LOGIC; 
  signal maccontrol_addr_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_addr_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_lrxbcast_FFY_RST : STD_LOGIC; 
  signal maccontrol_addr_0_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_addr_1_1_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_11_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_13_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_13_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_dout_15_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_11_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_11_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_1_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_3_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_3_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_5_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_5_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_7_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_7_FFX_RST : STD_LOGIC; 
  signal memtest_dataw1_9_FFY_RST : STD_LOGIC; 
  signal memtest_dataw1_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_phydi_2_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_3_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_11_FFY_RST : STD_LOGIC; 
  signal maccontrol_phydi_5_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_din_9_FFY_RST : STD_LOGIC; 
  signal maccontrol_din_9_FFX_RST : STD_LOGIC; 
  signal clkslen_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_7_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_9_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_din_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_sclkdeltal_FFY_RST : STD_LOGIC; 
  signal memcontroller_oel_FFY_RST : STD_LOGIC; 
  signal maccontrol_lrxallf_FFY_SET : STD_LOGIC; 
  signal memtest2_deql_0_FFY_RST : STD_LOGIC; 
  signal memtest2_deql_0_FFX_RST : STD_LOGIC; 
  signal txsim_ltxd_1_FFY_RST : STD_LOGIC; 
  signal txsim_ltxd_1_FFX_RST : STD_LOGIC; 
  signal txsim_ltxd_3_FFY_RST : STD_LOGIC; 
  signal txsim_ltxd_3_FFX_RST : STD_LOGIC; 
  signal txsim_ltxd_5_FFY_RST : STD_LOGIC; 
  signal txsim_ltxd_5_FFX_RST : STD_LOGIC; 
  signal txsim_ltxd_7_FFY_RST : STD_LOGIC; 
  signal txsim_ltxd_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_2_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_2_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_4_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_dreg_6_FFY_RST : STD_LOGIC; 
  signal addr2_1_FFY_RST : STD_LOGIC; 
  signal addr2_1_FFX_RST : STD_LOGIC; 
  signal addr2_3_FFY_RST : STD_LOGIC; 
  signal addr2_3_FFX_RST : STD_LOGIC; 
  signal addr2_5_FFY_RST : STD_LOGIC; 
  signal addr2_5_FFX_RST : STD_LOGIC; 
  signal addr2_7_FFY_RST : STD_LOGIC; 
  signal addr2_7_FFX_RST : STD_LOGIC; 
  signal mwe2_FFY_RST : STD_LOGIC; 
  signal addr2_9_FFY_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_rwl_FFY_RST : STD_LOGIC; 
  signal addr2_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_29_FFX_RST : STD_LOGIC; 
  signal memtest_addrcntl_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_PHY_status_MII_Interface_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal maccontrol_lrxucast_FFY_RST : STD_LOGIC; 
  signal memtest2_laddr_1_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_13_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_21_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_21_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_13_FFX_RST : STD_LOGIC; 
  signal memtest_addrcntl_1_FFY_RST : STD_LOGIC; 
  signal memtest_addrcntl_1_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_23_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_23_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_31_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_31_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_15_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_15_FFX_RST : STD_LOGIC; 
  signal memtest_addrcntl_3_FFY_RST : STD_LOGIC; 
  signal memtest_addrcntl_3_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_25_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_17_FFY_RST : STD_LOGIC; 
  signal memtest2_laddr_1_FFX_RST : STD_LOGIC; 
  signal memtest2_laddr_3_FFX_RST : STD_LOGIC; 
  signal memtest2_laddr_11_FFY_RST : STD_LOGIC; 
  signal memtest2_laddr_11_FFX_RST : STD_LOGIC; 
  signal memtest2_laddr_5_FFX_RST : STD_LOGIC; 
  signal memtest2_laddr_13_FFX_RST : STD_LOGIC; 
  signal memtest2_laddr_7_FFY_RST : STD_LOGIC; 
  signal memtest2_laddr_7_FFX_RST : STD_LOGIC; 
  signal memtest2_laddr_15_FFX_RST : STD_LOGIC; 
  signal memtest2_laddr_9_FFY_RST : STD_LOGIC; 
  signal memtest2_laddr_9_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_25_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_17_FFX_RST : STD_LOGIC; 
  signal memtest_addrcntl_5_FFY_RST : STD_LOGIC; 
  signal memtest_addrcntl_5_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_27_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_27_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_19_FFY_RST : STD_LOGIC; 
  signal maccontrol_phystat_19_FFX_RST : STD_LOGIC; 
  signal memtest_addrcntl_7_FFY_RST : STD_LOGIC; 
  signal memtest_addrcntl_7_FFX_RST : STD_LOGIC; 
  signal maccontrol_phystat_29_FFY_RST : STD_LOGIC; 
  signal memtest_addrcntl_9_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_1_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_1_FFX_RST : STD_LOGIC; 
  signal d2_1_FFY_RST : STD_LOGIC; 
  signal d2_2_FFY_RST : STD_LOGIC; 
  signal d2_5_FFY_RST : STD_LOGIC; 
  signal d2_5_FFX_RST : STD_LOGIC; 
  signal d2_7_FFY_RST : STD_LOGIC; 
  signal d2_7_FFX_RST : STD_LOGIC; 
  signal d2_9_FFY_RST : STD_LOGIC; 
  signal d2_9_FFX_RST : STD_LOGIC; 
  signal addr2_11_FFY_RST : STD_LOGIC; 
  signal addr2_11_FFX_RST : STD_LOGIC; 
  signal ifclk_bufg_CE : STD_LOGIC; 
  signal rx_clk_bufg_CE : STD_LOGIC; 
  signal clk_bufg_CE : STD_LOGIC; 
  signal PWR_VCC_0_FROM : STD_LOGIC; 
  signal PWR_VCC_0_GROM : STD_LOGIC; 
  signal PWR_VCC_1_FROM : STD_LOGIC; 
  signal PWR_VCC_2_FROM : STD_LOGIC; 
  signal PWR_VCC_3_FROM : STD_LOGIC; 
  signal PWR_VCC_4_FROM : STD_LOGIC; 
  signal PWR_VCC_5_FROM : STD_LOGIC; 
  signal PWR_VCC_5_GROM : STD_LOGIC; 
  signal PWR_VCC_6_FROM : STD_LOGIC; 
  signal PWR_VCC_7_FROM : STD_LOGIC; 
  signal PWR_VCC_7_GROM : STD_LOGIC; 
  signal PWR_VCC_8_FROM : STD_LOGIC; 
  signal PWR_VCC_9_FROM : STD_LOGIC; 
  signal PWR_VCC_10_FROM : STD_LOGIC; 
  signal PWR_VCC_11_FROM : STD_LOGIC; 
  signal PWR_VCC_12_FROM : STD_LOGIC; 
  signal PWR_VCC_13_FROM : STD_LOGIC; 
  signal PWR_VCC_14_FROM : STD_LOGIC; 
  signal PWR_VCC_15_FROM : STD_LOGIC; 
  signal PWR_VCC_16_FROM : STD_LOGIC; 
  signal PWR_VCC_17_FROM : STD_LOGIC; 
  signal PWR_VCC_18_FROM : STD_LOGIC; 
  signal PWR_VCC_18_GROM : STD_LOGIC; 
  signal PWR_VCC_19_FROM : STD_LOGIC; 
  signal PWR_VCC_19_GROM : STD_LOGIC; 
  signal PWR_VCC_20_FROM : STD_LOGIC; 
  signal PWR_VCC_21_FROM : STD_LOGIC; 
  signal PWR_VCC_22_FROM : STD_LOGIC; 
  signal PWR_VCC_23_FROM : STD_LOGIC; 
  signal PWR_VCC_24_FROM : STD_LOGIC; 
  signal PWR_VCC_25_FROM : STD_LOGIC; 
  signal PWR_VCC_26_FROM : STD_LOGIC; 
  signal PWR_VCC_27_FROM : STD_LOGIC; 
  signal PWR_VCC_28_FROM : STD_LOGIC; 
  signal PWR_VCC_28_GROM : STD_LOGIC; 
  signal PWR_VCC_29_FROM : STD_LOGIC; 
  signal PWR_VCC_29_GROM : STD_LOGIC; 
  signal PWR_VCC_30_FROM : STD_LOGIC; 
  signal PWR_VCC_31_FROM : STD_LOGIC; 
  signal PWR_VCC_32_FROM : STD_LOGIC; 
  signal PWR_VCC_32_GROM : STD_LOGIC; 
  signal PWR_VCC_33_FROM : STD_LOGIC; 
  signal PWR_VCC_33_GROM : STD_LOGIC; 
  signal PWR_VCC_34_FROM : STD_LOGIC; 
  signal PWR_VCC_34_GROM : STD_LOGIC; 
  signal PWR_VCC_35_FROM : STD_LOGIC; 
  signal PWR_VCC_35_GROM : STD_LOGIC; 
  signal PWR_VCC_36_FROM : STD_LOGIC; 
  signal PWR_VCC_37_FROM : STD_LOGIC; 
  signal PWR_VCC_37_GROM : STD_LOGIC; 
  signal PWR_VCC_38_FROM : STD_LOGIC; 
  signal PWR_VCC_38_GROM : STD_LOGIC; 
  signal PWR_VCC_39_FROM : STD_LOGIC; 
  signal PWR_VCC_39_GROM : STD_LOGIC; 
  signal PWR_VCC_40_FROM : STD_LOGIC; 
  signal PWR_VCC_40_GROM : STD_LOGIC; 
  signal PWR_VCC_41_FROM : STD_LOGIC; 
  signal PWR_VCC_41_GROM : STD_LOGIC; 
  signal PWR_VCC_42_FROM : STD_LOGIC; 
  signal PWR_VCC_42_GROM : STD_LOGIC; 
  signal PWR_VCC_43_FROM : STD_LOGIC; 
  signal PWR_VCC_44_FROM : STD_LOGIC; 
  signal PWR_VCC_45_FROM : STD_LOGIC; 
  signal PWR_VCC_46_FROM : STD_LOGIC; 
  signal PWR_VCC_46_GROM : STD_LOGIC; 
  signal PWR_VCC_47_FROM : STD_LOGIC; 
  signal PWR_GND_0_GROM : STD_LOGIC; 
  signal PWR_GND_1_GROM : STD_LOGIC; 
  signal PWR_GND_2_GROM : STD_LOGIC; 
  signal PWR_GND_3_GROM : STD_LOGIC; 
  signal PWR_GND_4_GROM : STD_LOGIC; 
  signal PWR_GND_5_GROM : STD_LOGIC; 
  signal PWR_GND_6_GROM : STD_LOGIC; 
  signal PWR_GND_7_GROM : STD_LOGIC; 
  signal PWR_GND_8_GROM : STD_LOGIC; 
  signal PWR_GND_9_GROM : STD_LOGIC; 
  signal PWR_GND_10_GROM : STD_LOGIC; 
  signal PWR_GND_11_GROM : STD_LOGIC; 
  signal PWR_GND_12_GROM : STD_LOGIC; 
  signal PWR_GND_13_GROM : STD_LOGIC; 
  signal PWR_GND_14_GROM : STD_LOGIC; 
  signal PWR_GND_15_GROM : STD_LOGIC; 
  signal PWR_GND_16_GROM : STD_LOGIC; 
  signal PWR_GND_17_GROM : STD_LOGIC; 
  signal PWR_GND_18_GROM : STD_LOGIC; 
  signal PWR_GND_19_GROM : STD_LOGIC; 
  signal PWR_GND_20_GROM : STD_LOGIC; 
  signal PWR_GND_21_GROM : STD_LOGIC; 
  signal PWR_GND_22_GROM : STD_LOGIC; 
  signal PWR_GND_23_GROM : STD_LOGIC; 
  signal PWR_GND_24_GROM : STD_LOGIC; 
  signal PWR_GND_25_GROM : STD_LOGIC; 
  signal PWR_GND_26_GROM : STD_LOGIC; 
  signal PWR_GND_27_GROM : STD_LOGIC; 
  signal PWR_GND_28_GROM : STD_LOGIC; 
  signal PWR_GND_29_GROM : STD_LOGIC; 
  signal PWR_GND_30_GROM : STD_LOGIC; 
  signal PWR_GND_31_GROM : STD_LOGIC; 
  signal PWR_GND_32_GROM : STD_LOGIC; 
  signal PWR_GND_33_GROM : STD_LOGIC; 
  signal PWR_GND_34_GROM : STD_LOGIC; 
  signal PWR_GND_35_GROM : STD_LOGIC; 
  signal PWR_GND_36_GROM : STD_LOGIC; 
  signal PWR_GND_37_GROM : STD_LOGIC; 
  signal PWR_GND_38_GROM : STD_LOGIC; 
  signal PWR_GND_39_GROM : STD_LOGIC; 
  signal PWR_GND_40_GROM : STD_LOGIC; 
  signal PWR_GND_41_GROM : STD_LOGIC; 
  signal PWR_GND_42_GROM : STD_LOGIC; 
  signal PWR_GND_43_GROM : STD_LOGIC; 
  signal PWR_GND_44_GROM : STD_LOGIC; 
  signal PWR_GND_45_GROM : STD_LOGIC; 
  signal PWR_GND_46_GROM : STD_LOGIC; 
  signal PWR_GND_47_GROM : STD_LOGIC; 
  signal PWR_GND_48_GROM : STD_LOGIC; 
  signal PWR_GND_49_GROM : STD_LOGIC; 
  signal PWR_GND_50_GROM : STD_LOGIC; 
  signal PWR_GND_51_GROM : STD_LOGIC; 
  signal PWR_GND_52_GROM : STD_LOGIC; 
  signal PWR_GND_53_GROM : STD_LOGIC; 
  signal GND : STD_LOGIC; 
  signal VCC : STD_LOGIC; 
  signal txsim_ltxd : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal testrx_macaddrl : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal memcontroller_addrn : STD_LOGIC_VECTOR ( 16 downto 0 ); 
  signal memcontroller_qn : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_dnl2 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal maccontrol_phystat : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal maccontrol_dout : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal testrx_lmacdata : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal maccontrol_PHY_status_MII_Interface_dreg : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal testrx_rxdl : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal Q_n0000 : STD_LOGIC_VECTOR ( 23 downto 1 ); 
  signal testrx_addr : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal testrx_rxdll : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal txsim_counter : STD_LOGIC_VECTOR ( 17 downto 0 ); 
  signal txsim_ramout : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal addr4 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal addr2 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal addr1 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal maccontrol_PHY_status_MII_Interface_statecnt : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal maccontrol_PHY_status_din : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal cnt0 : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal memtest2_datain : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memtest2_deq : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal cnt : STD_LOGIC_VECTOR ( 23 downto 0 ); 
  signal maccontrol_PHY_status_MII_Interface_mdccnt : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal q4 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memtest2_cnt : STD_LOGIC_VECTOR ( 16 downto 0 ); 
  signal maccontrol_PHY_status_MII_Interface_n0078 : STD_LOGIC_VECTOR ( 5 downto 1 ); 
  signal d1 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memtest2_laddr : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal memcontroller_clknum : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal memtest2_cs : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal q2 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memtest2_ldata : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal maccontrol_addr : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal maccontrol_phyaddr : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal d2 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal maccontrol_phydo : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal maccontrol_lmacaddr : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal maccontrol_phydi : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memtest_dataw1 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_dnl1 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_clknum_n0001 : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal memtest2_datalfsr : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal clken_clkcnt : STD_LOGIC_VECTOR ( 2 downto 0 ); 
  signal memtest2_addrlfsr : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal maccontrol_PHY_status_dout : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal memtest_addrcntl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal maccontrol_din : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal maccontrol_PHY_status_addrl : STD_LOGIC_VECTOR ( 4 downto 0 ); 
  signal maccontrol_PHY_status_miiaddr : STD_LOGIC_VECTOR ( 4 downto 0 ); 
  signal memtest2_deql : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal memcontroller_ADDREXT : STD_LOGIC_VECTOR ( 16 downto 0 ); 
  signal memcontroller_ts : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_dnout : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_q : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal cnt0_n0000 : STD_LOGIC_VECTOR ( 5 downto 1 ); 
  signal testrx_addr_n0000 : STD_LOGIC_VECTOR ( 7 downto 1 ); 
  signal memtest2_cnt_n0000 : STD_LOGIC_VECTOR ( 16 downto 1 ); 
  signal txsim_counter_n0000 : STD_LOGIC_VECTOR ( 17 downto 1 ); 
  signal memtest_datacnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal memtest_addrcnt_n0000 : STD_LOGIC_VECTOR ( 15 downto 1 ); 
  signal memcontroller_dn : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal maccontrol_PHY_status_MII_Interface_n0014 : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal clken_clkcnt_n0000 : STD_LOGIC_VECTOR ( 2 downto 1 ); 
begin
  SCLK_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => SCLK_IFF_RST
    );
  maccontrol_sclkl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_SCLK_IBUF,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => SCLK_IFF_RST,
      O => maccontrol_sclkl
    );
  maccontrol_SCLK_IBUF_7 : X_BUF
    port map (
      I => SCLK,
      O => maccontrol_SCLK_IBUF
    );
  TESTOUT_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TESTOUT_OFF_RST
    );
  memtest2_ERR_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TESTOUT_OD,
      CE => memtest2_n0119,
      CLK => clk,
      SET => GND,
      RST => TESTOUT_OFF_RST,
      O => memtest2_ERR
    );
  memtest2_TESTOUT_OBUF : X_TRI
    port map (
      I => TESTOUT_OUTMUX,
      CTL => TESTOUT_ENABLE,
      O => TESTOUT
    );
  TESTOUT_ENABLEINV : X_INV
    port map (
      I => TESTOUT_TORGTS,
      O => TESTOUT_ENABLE
    );
  TESTOUT_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TESTOUT_TORGTS
    );
  TESTOUT_OUTMUX_9 : X_BUF
    port map (
      I => memtest2_ERR,
      O => TESTOUT_OUTMUX
    );
  TESTOUT_OMUX : X_BUF
    port map (
      I => memtest2_n0030,
      O => TESTOUT_OD
    );
  TXD_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_0_OFF_RST
    );
  txsim_TXD_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_0_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => TXD_0_OFF_RST,
      O => txsim_TXD_0_OBUF
    );
  txsim_TXD_0_OBUF_10 : X_TRI
    port map (
      I => TXD_0_OUTMUX,
      CTL => TXD_0_ENABLE,
      O => TXD(0)
    );
  TXD_0_ENABLEINV : X_INV
    port map (
      I => TXD_0_TORGTS,
      O => TXD_0_ENABLE
    );
  TXD_0_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_0_TORGTS
    );
  TXD_0_OUTMUX_11 : X_BUF
    port map (
      I => txsim_TXD_0_OBUF,
      O => TXD_0_OUTMUX
    );
  TXD_0_OMUX : X_BUF
    port map (
      I => txsim_ltxd(0),
      O => TXD_0_OD
    );
  TXD_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_1_OFF_RST
    );
  txsim_TXD_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_1_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => TXD_1_OFF_RST,
      O => txsim_TXD_1_OBUF
    );
  txsim_TXD_1_OBUF_12 : X_TRI
    port map (
      I => TXD_1_OUTMUX,
      CTL => TXD_1_ENABLE,
      O => TXD(1)
    );
  TXD_1_ENABLEINV : X_INV
    port map (
      I => TXD_1_TORGTS,
      O => TXD_1_ENABLE
    );
  TXD_1_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_1_TORGTS
    );
  TXD_1_OUTMUX_13 : X_BUF
    port map (
      I => txsim_TXD_1_OBUF,
      O => TXD_1_OUTMUX
    );
  TXD_1_OMUX : X_BUF
    port map (
      I => txsim_ltxd(1),
      O => TXD_1_OD
    );
  TXD_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_2_OFF_RST
    );
  txsim_TXD_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_2_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => TXD_2_OFF_RST,
      O => txsim_TXD_2_OBUF
    );
  txsim_TXD_2_OBUF_14 : X_TRI
    port map (
      I => TXD_2_OUTMUX,
      CTL => TXD_2_ENABLE,
      O => TXD(2)
    );
  TXD_2_ENABLEINV : X_INV
    port map (
      I => TXD_2_TORGTS,
      O => TXD_2_ENABLE
    );
  TXD_2_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_2_TORGTS
    );
  TXD_2_OUTMUX_15 : X_BUF
    port map (
      I => txsim_TXD_2_OBUF,
      O => TXD_2_OUTMUX
    );
  TXD_2_OMUX : X_BUF
    port map (
      I => txsim_ltxd(2),
      O => TXD_2_OD
    );
  TXD_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_3_OFF_RST
    );
  txsim_TXD_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_3_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => TXD_3_OFF_RST,
      O => txsim_TXD_3_OBUF
    );
  txsim_TXD_3_OBUF_16 : X_TRI
    port map (
      I => TXD_3_OUTMUX,
      CTL => TXD_3_ENABLE,
      O => TXD(3)
    );
  TXD_3_ENABLEINV : X_INV
    port map (
      I => TXD_3_TORGTS,
      O => TXD_3_ENABLE
    );
  TXD_3_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_3_TORGTS
    );
  TXD_3_OUTMUX_17 : X_BUF
    port map (
      I => txsim_TXD_3_OBUF,
      O => TXD_3_OUTMUX
    );
  TXD_3_OMUX : X_BUF
    port map (
      I => txsim_ltxd(3),
      O => TXD_3_OD
    );
  TXD_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_4_OFF_RST
    );
  txsim_TXD_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_4_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => TXD_4_OFF_RST,
      O => txsim_TXD_4_OBUF
    );
  txsim_TXD_4_OBUF_18 : X_TRI
    port map (
      I => TXD_4_OUTMUX,
      CTL => TXD_4_ENABLE,
      O => TXD(4)
    );
  TXD_4_ENABLEINV : X_INV
    port map (
      I => TXD_4_TORGTS,
      O => TXD_4_ENABLE
    );
  TXD_4_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_4_TORGTS
    );
  TXD_4_OUTMUX_19 : X_BUF
    port map (
      I => txsim_TXD_4_OBUF,
      O => TXD_4_OUTMUX
    );
  TXD_4_OMUX : X_BUF
    port map (
      I => txsim_ltxd(4),
      O => TXD_4_OD
    );
  TXD_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_5_OFF_RST
    );
  txsim_TXD_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_5_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => TXD_5_OFF_RST,
      O => txsim_TXD_5_OBUF
    );
  txsim_TXD_5_OBUF_20 : X_TRI
    port map (
      I => TXD_5_OUTMUX,
      CTL => TXD_5_ENABLE,
      O => TXD(5)
    );
  TXD_5_ENABLEINV : X_INV
    port map (
      I => TXD_5_TORGTS,
      O => TXD_5_ENABLE
    );
  TXD_5_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_5_TORGTS
    );
  TXD_5_OUTMUX_21 : X_BUF
    port map (
      I => txsim_TXD_5_OBUF,
      O => TXD_5_OUTMUX
    );
  TXD_5_OMUX : X_BUF
    port map (
      I => txsim_ltxd(5),
      O => TXD_5_OD
    );
  TXD_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_6_OFF_RST
    );
  txsim_TXD_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_6_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => TXD_6_OFF_RST,
      O => txsim_TXD_6_OBUF
    );
  txsim_TXD_6_OBUF_22 : X_TRI
    port map (
      I => TXD_6_OUTMUX,
      CTL => TXD_6_ENABLE,
      O => TXD(6)
    );
  TXD_6_ENABLEINV : X_INV
    port map (
      I => TXD_6_TORGTS,
      O => TXD_6_ENABLE
    );
  TXD_6_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_6_TORGTS
    );
  TXD_6_OUTMUX_23 : X_BUF
    port map (
      I => txsim_TXD_6_OBUF,
      O => TXD_6_OUTMUX
    );
  TXD_6_OMUX : X_BUF
    port map (
      I => txsim_ltxd(6),
      O => TXD_6_OD
    );
  txsim_TXD_7_OBUF_24 : X_TRI
    port map (
      I => TXD_7_OUTMUX,
      CTL => TXD_7_ENABLE,
      O => TXD(7)
    );
  TXD_7_ENABLEINV : X_INV
    port map (
      I => TXD_7_TORGTS,
      O => TXD_7_ENABLE
    );
  TXD_7_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_7_TORGTS
    );
  TXD_7_OUTMUX_25 : X_BUF
    port map (
      I => txsim_TXD_7_OBUF,
      O => TXD_7_OUTMUX
    );
  TXD_7_OMUX : X_BUF
    port map (
      I => txsim_ltxd(7),
      O => TXD_7_OD
    );
  testrx_MACADDR_0_IBUF_26 : X_BUF
    port map (
      I => MACADDR(0),
      O => testrx_MACADDR_0_IBUF
    );
  testrx_MACADDR_1_IBUF_27 : X_BUF
    port map (
      I => MACADDR(1),
      O => testrx_MACADDR_1_IBUF
    );
  testrx_MACADDR_2_IBUF_28 : X_BUF
    port map (
      I => MACADDR(2),
      O => testrx_MACADDR_2_IBUF
    );
  testrx_MACADDR_3_IBUF_29 : X_BUF
    port map (
      I => MACADDR(3),
      O => testrx_MACADDR_3_IBUF
    );
  testrx_MACADDR_4_IBUF_30 : X_BUF
    port map (
      I => MACADDR(4),
      O => testrx_MACADDR_4_IBUF
    );
  testrx_MACADDR_5_IBUF_31 : X_BUF
    port map (
      I => MACADDR(5),
      O => testrx_MACADDR_5_IBUF
    );
  testrx_MACADDR_6_IBUF_32 : X_BUF
    port map (
      I => MACADDR(6),
      O => testrx_MACADDR_6_IBUF
    );
  testrx_MACADDR_7_IBUF_33 : X_BUF
    port map (
      I => MACADDR(7),
      O => testrx_MACADDR_7_IBUF
    );
  MCLK_OBUF_34 : X_TRI
    port map (
      I => MCLK_OUTMUX,
      CTL => MCLK_ENABLE,
      O => MCLK
    );
  MCLK_ENABLEINV : X_INV
    port map (
      I => MCLK_TORGTS,
      O => MCLK_ENABLE
    );
  MCLK_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MCLK_TORGTS
    );
  MCLK_OUTMUX_35 : X_BUF
    port map (
      I => MCLK_OBUF,
      O => MCLK_OUTMUX
    );
  memcontroller_MA_0_OBUF : X_TRI
    port map (
      I => MA_0_OUTMUX,
      CTL => MA_0_ENABLE,
      O => MA(0)
    );
  MA_0_ENABLEINV : X_INV
    port map (
      I => MA_0_TORGTS,
      O => MA_0_ENABLE
    );
  MA_0_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_0_TORGTS
    );
  MA_0_OUTMUX_36 : X_BUF
    port map (
      I => memcontroller_ADDREXT(0),
      O => MA_0_OUTMUX
    );
  MA_0_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_0_OCEMUXNOT
    );
  MA_0_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(0),
      O => MA_0_OD
    );
  memcontroller_MA_1_OBUF : X_TRI
    port map (
      I => MA_1_OUTMUX,
      CTL => MA_1_ENABLE,
      O => MA(1)
    );
  MA_1_ENABLEINV : X_INV
    port map (
      I => MA_1_TORGTS,
      O => MA_1_ENABLE
    );
  MA_1_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_1_TORGTS
    );
  MA_1_OUTMUX_37 : X_BUF
    port map (
      I => memcontroller_ADDREXT(1),
      O => MA_1_OUTMUX
    );
  MA_1_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_1_OCEMUXNOT
    );
  MA_1_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(1),
      O => MA_1_OD
    );
  memcontroller_MA_2_OBUF : X_TRI
    port map (
      I => MA_2_OUTMUX,
      CTL => MA_2_ENABLE,
      O => MA(2)
    );
  MA_2_ENABLEINV : X_INV
    port map (
      I => MA_2_TORGTS,
      O => MA_2_ENABLE
    );
  MA_2_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_2_TORGTS
    );
  MA_2_OUTMUX_38 : X_BUF
    port map (
      I => memcontroller_ADDREXT(2),
      O => MA_2_OUTMUX
    );
  MA_2_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_2_OCEMUXNOT
    );
  MA_2_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(2),
      O => MA_2_OD
    );
  memcontroller_MA_3_OBUF : X_TRI
    port map (
      I => MA_3_OUTMUX,
      CTL => MA_3_ENABLE,
      O => MA(3)
    );
  MA_3_ENABLEINV : X_INV
    port map (
      I => MA_3_TORGTS,
      O => MA_3_ENABLE
    );
  MA_3_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_3_TORGTS
    );
  MA_3_OUTMUX_39 : X_BUF
    port map (
      I => memcontroller_ADDREXT(3),
      O => MA_3_OUTMUX
    );
  MA_3_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_3_OCEMUXNOT
    );
  MA_3_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(3),
      O => MA_3_OD
    );
  memcontroller_MA_4_OBUF : X_TRI
    port map (
      I => MA_4_OUTMUX,
      CTL => MA_4_ENABLE,
      O => MA(4)
    );
  MA_4_ENABLEINV : X_INV
    port map (
      I => MA_4_TORGTS,
      O => MA_4_ENABLE
    );
  MA_4_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_4_TORGTS
    );
  MA_4_OUTMUX_40 : X_BUF
    port map (
      I => memcontroller_ADDREXT(4),
      O => MA_4_OUTMUX
    );
  MA_4_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_4_OCEMUXNOT
    );
  MA_4_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(4),
      O => MA_4_OD
    );
  txsim_TXD_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_7_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => TXD_7_OFF_RST,
      O => txsim_TXD_7_OBUF
    );
  TXD_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_7_OFF_RST
    );
  memcontroller_MA_5_OBUF : X_TRI
    port map (
      I => MA_5_OUTMUX,
      CTL => MA_5_ENABLE,
      O => MA(5)
    );
  MA_5_ENABLEINV : X_INV
    port map (
      I => MA_5_TORGTS,
      O => MA_5_ENABLE
    );
  MA_5_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_5_TORGTS
    );
  MA_5_OUTMUX_41 : X_BUF
    port map (
      I => memcontroller_ADDREXT(5),
      O => MA_5_OUTMUX
    );
  MA_5_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_5_OCEMUXNOT
    );
  MA_5_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(5),
      O => MA_5_OD
    );
  memcontroller_MA_6_OBUF : X_TRI
    port map (
      I => MA_6_OUTMUX,
      CTL => MA_6_ENABLE,
      O => MA(6)
    );
  MA_6_ENABLEINV : X_INV
    port map (
      I => MA_6_TORGTS,
      O => MA_6_ENABLE
    );
  MA_6_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_6_TORGTS
    );
  MA_6_OUTMUX_42 : X_BUF
    port map (
      I => memcontroller_ADDREXT(6),
      O => MA_6_OUTMUX
    );
  MA_6_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_6_OCEMUXNOT
    );
  MA_6_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(6),
      O => MA_6_OD
    );
  memcontroller_MA_7_OBUF : X_TRI
    port map (
      I => MA_7_OUTMUX,
      CTL => MA_7_ENABLE,
      O => MA(7)
    );
  MA_7_ENABLEINV : X_INV
    port map (
      I => MA_7_TORGTS,
      O => MA_7_ENABLE
    );
  MA_7_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_7_TORGTS
    );
  MA_7_OUTMUX_43 : X_BUF
    port map (
      I => memcontroller_ADDREXT(7),
      O => MA_7_OUTMUX
    );
  MA_7_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_7_OCEMUXNOT
    );
  MA_7_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(7),
      O => MA_7_OD
    );
  memcontroller_MA_8_OBUF : X_TRI
    port map (
      I => MA_8_OUTMUX,
      CTL => MA_8_ENABLE,
      O => MA(8)
    );
  MA_8_ENABLEINV : X_INV
    port map (
      I => MA_8_TORGTS,
      O => MA_8_ENABLE
    );
  MA_8_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_8_TORGTS
    );
  MA_8_OUTMUX_44 : X_BUF
    port map (
      I => memcontroller_ADDREXT(8),
      O => MA_8_OUTMUX
    );
  MA_8_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_8_OCEMUXNOT
    );
  MA_8_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(8),
      O => MA_8_OD
    );
  memcontroller_MA_9_OBUF : X_TRI
    port map (
      I => MA_9_OUTMUX,
      CTL => MA_9_ENABLE,
      O => MA(9)
    );
  MA_9_ENABLEINV : X_INV
    port map (
      I => MA_9_TORGTS,
      O => MA_9_ENABLE
    );
  MA_9_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_9_TORGTS
    );
  MA_9_OUTMUX_45 : X_BUF
    port map (
      I => memcontroller_ADDREXT(9),
      O => MA_9_OUTMUX
    );
  MA_9_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_9_OCEMUXNOT
    );
  MA_9_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(9),
      O => MA_9_OD
    );
  memcontroller_qdout0_OBUFT : X_TRI
    port map (
      I => MD_0_OUTMUX,
      CTL => MD_0_ENABLE,
      O => MD(0)
    );
  MD_0_ENABLEINV : X_INV
    port map (
      I => MD_0_TORGTS,
      O => MD_0_ENABLE
    );
  MD_0_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_0_TORGTS
    );
  MD_0_OUTMUX_46 : X_BUF
    port map (
      I => memcontroller_dnout(0),
      O => MD_0_OUTMUX
    );
  MD_0_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(0),
      O => MD_0_OD
    );
  memcontroller_qdout0_IBUF : X_BUF
    port map (
      I => MD(0),
      O => memcontroller_q(0)
    );
  memcontroller_qdout1_OBUFT : X_TRI
    port map (
      I => MD_1_OUTMUX,
      CTL => MD_1_ENABLE,
      O => MD(1)
    );
  MD_1_ENABLEINV : X_INV
    port map (
      I => MD_1_TORGTS,
      O => MD_1_ENABLE
    );
  MD_1_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(1),
      O => MD_1_TORGTS
    );
  MD_1_OUTMUX_47 : X_BUF
    port map (
      I => memcontroller_dnout(1),
      O => MD_1_OUTMUX
    );
  MD_1_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(1),
      O => MD_1_OD
    );
  memcontroller_qdout1_IBUF : X_BUF
    port map (
      I => MD(1),
      O => memcontroller_q(1)
    );
  txsim_TX_EN_OBUF_48 : X_TRI
    port map (
      I => TX_EN_OUTMUX,
      CTL => TX_EN_ENABLE,
      O => TX_EN
    );
  TX_EN_ENABLEINV : X_INV
    port map (
      I => TX_EN_TORGTS,
      O => TX_EN_ENABLE
    );
  TX_EN_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TX_EN_TORGTS
    );
  TX_EN_OUTMUX_49 : X_BUF
    port map (
      I => txsim_TX_EN_OBUF,
      O => TX_EN_OUTMUX
    );
  TX_EN_OMUX : X_BUF
    port map (
      I => txsim_Mshreg_TX_EN_net129,
      O => TX_EN_OD
    );
  memcontroller_qdout2_OBUFT : X_TRI
    port map (
      I => MD_2_OUTMUX,
      CTL => MD_2_ENABLE,
      O => MD(2)
    );
  MD_2_ENABLEINV : X_INV
    port map (
      I => MD_2_TORGTS,
      O => MD_2_ENABLE
    );
  MD_2_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(2),
      O => MD_2_TORGTS
    );
  MD_2_OUTMUX_50 : X_BUF
    port map (
      I => memcontroller_dnout(2),
      O => MD_2_OUTMUX
    );
  MD_2_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(2),
      O => MD_2_OD
    );
  memcontroller_qdout2_IBUF : X_BUF
    port map (
      I => MD(2),
      O => memcontroller_q(2)
    );
  memcontroller_qdout3_OBUFT : X_TRI
    port map (
      I => MD_3_OUTMUX,
      CTL => MD_3_ENABLE,
      O => MD(3)
    );
  MD_3_ENABLEINV : X_INV
    port map (
      I => MD_3_TORGTS,
      O => MD_3_ENABLE
    );
  MD_3_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(3),
      O => MD_3_TORGTS
    );
  MD_3_OUTMUX_51 : X_BUF
    port map (
      I => memcontroller_dnout(3),
      O => MD_3_OUTMUX
    );
  MD_3_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(3),
      O => MD_3_OD
    );
  memcontroller_qdout3_IBUF : X_BUF
    port map (
      I => MD(3),
      O => memcontroller_q(3)
    );
  memcontroller_qdout4_OBUFT : X_TRI
    port map (
      I => MD_4_OUTMUX,
      CTL => MD_4_ENABLE,
      O => MD(4)
    );
  MD_4_ENABLEINV : X_INV
    port map (
      I => MD_4_TORGTS,
      O => MD_4_ENABLE
    );
  MD_4_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(4),
      O => MD_4_TORGTS
    );
  MD_4_OUTMUX_52 : X_BUF
    port map (
      I => memcontroller_dnout(4),
      O => MD_4_OUTMUX
    );
  MD_4_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(4),
      O => MD_4_OD
    );
  memcontroller_qdout4_IBUF : X_BUF
    port map (
      I => MD(4),
      O => memcontroller_q(4)
    );
  memcontroller_qdout5_OBUFT : X_TRI
    port map (
      I => MD_5_OUTMUX,
      CTL => MD_5_ENABLE,
      O => MD(5)
    );
  MD_5_ENABLEINV : X_INV
    port map (
      I => MD_5_TORGTS,
      O => MD_5_ENABLE
    );
  MD_5_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(5),
      O => MD_5_TORGTS
    );
  MD_5_OUTMUX_53 : X_BUF
    port map (
      I => memcontroller_dnout(5),
      O => MD_5_OUTMUX
    );
  MD_5_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(5),
      O => MD_5_OD
    );
  memcontroller_qdout5_IBUF : X_BUF
    port map (
      I => MD(5),
      O => memcontroller_q(5)
    );
  memcontroller_qdout6_OBUFT : X_TRI
    port map (
      I => MD_6_OUTMUX,
      CTL => MD_6_ENABLE,
      O => MD(6)
    );
  MD_6_ENABLEINV : X_INV
    port map (
      I => MD_6_TORGTS,
      O => MD_6_ENABLE
    );
  MD_6_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(6),
      O => MD_6_TORGTS
    );
  MD_6_OUTMUX_54 : X_BUF
    port map (
      I => memcontroller_dnout(6),
      O => MD_6_OUTMUX
    );
  MD_6_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(6),
      O => MD_6_OD
    );
  memcontroller_qdout6_IBUF : X_BUF
    port map (
      I => MD(6),
      O => memcontroller_q(6)
    );
  memcontroller_qdout7_OBUFT : X_TRI
    port map (
      I => MD_7_OUTMUX,
      CTL => MD_7_ENABLE,
      O => MD(7)
    );
  MD_7_ENABLEINV : X_INV
    port map (
      I => MD_7_TORGTS,
      O => MD_7_ENABLE
    );
  MD_7_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(7),
      O => MD_7_TORGTS
    );
  MD_7_OUTMUX_55 : X_BUF
    port map (
      I => memcontroller_dnout(7),
      O => MD_7_OUTMUX
    );
  MD_7_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(7),
      O => MD_7_OD
    );
  memcontroller_qdout7_IBUF : X_BUF
    port map (
      I => MD(7),
      O => memcontroller_q(7)
    );
  memcontroller_qdout8_OBUFT : X_TRI
    port map (
      I => MD_8_OUTMUX,
      CTL => MD_8_ENABLE,
      O => MD(8)
    );
  MD_8_ENABLEINV : X_INV
    port map (
      I => MD_8_TORGTS,
      O => MD_8_ENABLE
    );
  MD_8_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(8),
      O => MD_8_TORGTS
    );
  MD_8_OUTMUX_56 : X_BUF
    port map (
      I => memcontroller_dnout(8),
      O => MD_8_OUTMUX
    );
  MD_8_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(8),
      O => MD_8_OD
    );
  memcontroller_qdout8_IBUF : X_BUF
    port map (
      I => MD(8),
      O => memcontroller_q(8)
    );
  memcontroller_qdout9_OBUFT : X_TRI
    port map (
      I => MD_9_OUTMUX,
      CTL => MD_9_ENABLE,
      O => MD(9)
    );
  MD_9_ENABLEINV : X_INV
    port map (
      I => MD_9_TORGTS,
      O => MD_9_ENABLE
    );
  MD_9_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(9),
      O => MD_9_TORGTS
    );
  MD_9_OUTMUX_57 : X_BUF
    port map (
      I => memcontroller_dnout(9),
      O => MD_9_OUTMUX
    );
  MD_9_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(9),
      O => MD_9_OD
    );
  memcontroller_qdout9_IBUF : X_BUF
    port map (
      I => MD(9),
      O => memcontroller_q(9)
    );
  LEDACT_OBUF_58 : X_TRI
    port map (
      I => LEDACT_OUTMUX,
      CTL => LEDACT_ENABLE,
      O => LEDACT
    );
  LEDACT_ENABLEINV : X_INV
    port map (
      I => LEDACT_TORGTS,
      O => LEDACT_ENABLE
    );
  LEDACT_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDACT_TORGTS
    );
  LEDACT_OUTMUX_59 : X_BUF
    port map (
      I => LEDACT_OBUF,
      O => LEDACT_OUTMUX
    );
  LEDACT_OCEMUX : X_INV
    port map (
      I => err,
      O => LEDACT_OCEMUXNOT
    );
  LEDACT_OMUX : X_BUF
    port map (
      I => Q_n0034,
      O => LEDACT_OD
    );
  testrx_macaddrl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_MACADDR_0_IBUF,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACADDR_0_IFF_RST,
      O => testrx_macaddrl(0)
    );
  MACADDR_0_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACADDR_0_IFF_RST
    );
  maccontrol_LEDDPX_OBUF_60 : X_TRI
    port map (
      I => LEDDPX_OUTMUX,
      CTL => LEDDPX_ENABLE,
      O => LEDDPX
    );
  LEDDPX_ENABLEINV : X_INV
    port map (
      I => LEDDPX_TORGTS,
      O => LEDDPX_ENABLE
    );
  LEDDPX_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDDPX_TORGTS
    );
  LEDDPX_OUTMUX_61 : X_BUF
    port map (
      I => maccontrol_LEDDPX_OBUF,
      O => LEDDPX_OUTMUX
    );
  LEDDPX_OMUX : X_BUF
    port map (
      I => maccontrol_phystat(1),
      O => LEDDPX_OD
    );
  LEDRX_LOGIC_ONE_62 : X_ONE
    port map (
      O => LEDRX_LOGIC_ONE
    );
  LEDRX_OBUF_63 : X_TRI
    port map (
      I => LEDRX_OUTMUX,
      CTL => LEDRX_ENABLE,
      O => LEDRX
    );
  LEDRX_ENABLEINV : X_INV
    port map (
      I => LEDRX_TORGTS,
      O => LEDRX_ENABLE
    );
  LEDRX_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDRX_TORGTS
    );
  LEDRX_OUTMUX_64 : X_BUF
    port map (
      I => LEDRX_OBUF,
      O => LEDRX_OUTMUX
    );
  memcontroller_MA_10_OBUF : X_TRI
    port map (
      I => MA_10_OUTMUX,
      CTL => MA_10_ENABLE,
      O => MA(10)
    );
  MA_10_ENABLEINV : X_INV
    port map (
      I => MA_10_TORGTS,
      O => MA_10_ENABLE
    );
  MA_10_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_10_TORGTS
    );
  MA_10_OUTMUX_65 : X_BUF
    port map (
      I => memcontroller_ADDREXT(10),
      O => MA_10_OUTMUX
    );
  MA_10_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_10_OCEMUXNOT
    );
  MA_10_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(10),
      O => MA_10_OD
    );
  memcontroller_MA_11_OBUF : X_TRI
    port map (
      I => MA_11_OUTMUX,
      CTL => MA_11_ENABLE,
      O => MA(11)
    );
  MA_11_ENABLEINV : X_INV
    port map (
      I => MA_11_TORGTS,
      O => MA_11_ENABLE
    );
  MA_11_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_11_TORGTS
    );
  MA_11_OUTMUX_66 : X_BUF
    port map (
      I => memcontroller_ADDREXT(11),
      O => MA_11_OUTMUX
    );
  MA_11_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_11_OCEMUXNOT
    );
  MA_11_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(11),
      O => MA_11_OD
    );
  memcontroller_MA_12_OBUF : X_TRI
    port map (
      I => MA_12_OUTMUX,
      CTL => MA_12_ENABLE,
      O => MA(12)
    );
  MA_12_ENABLEINV : X_INV
    port map (
      I => MA_12_TORGTS,
      O => MA_12_ENABLE
    );
  MA_12_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_12_TORGTS
    );
  MA_12_OUTMUX_67 : X_BUF
    port map (
      I => memcontroller_ADDREXT(12),
      O => MA_12_OUTMUX
    );
  MA_12_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_12_OCEMUXNOT
    );
  MA_12_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(12),
      O => MA_12_OD
    );
  memcontroller_MA_13_OBUF : X_TRI
    port map (
      I => MA_13_OUTMUX,
      CTL => MA_13_ENABLE,
      O => MA(13)
    );
  MA_13_ENABLEINV : X_INV
    port map (
      I => MA_13_TORGTS,
      O => MA_13_ENABLE
    );
  MA_13_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_13_TORGTS
    );
  MA_13_OUTMUX_68 : X_BUF
    port map (
      I => memcontroller_ADDREXT(13),
      O => MA_13_OUTMUX
    );
  MA_13_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_13_OCEMUXNOT
    );
  MA_13_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(13),
      O => MA_13_OD
    );
  memcontroller_MA_14_OBUF : X_TRI
    port map (
      I => MA_14_OUTMUX,
      CTL => MA_14_ENABLE,
      O => MA(14)
    );
  MA_14_ENABLEINV : X_INV
    port map (
      I => MA_14_TORGTS,
      O => MA_14_ENABLE
    );
  MA_14_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_14_TORGTS
    );
  MA_14_OUTMUX_69 : X_BUF
    port map (
      I => memcontroller_ADDREXT(14),
      O => MA_14_OUTMUX
    );
  MA_14_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_14_OCEMUXNOT
    );
  MA_14_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(14),
      O => MA_14_OD
    );
  memcontroller_MA_15_OBUF : X_TRI
    port map (
      I => MA_15_OUTMUX,
      CTL => MA_15_ENABLE,
      O => MA(15)
    );
  MA_15_ENABLEINV : X_INV
    port map (
      I => MA_15_TORGTS,
      O => MA_15_ENABLE
    );
  MA_15_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_15_TORGTS
    );
  MA_15_OUTMUX_70 : X_BUF
    port map (
      I => memcontroller_ADDREXT(15),
      O => MA_15_OUTMUX
    );
  MA_15_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_15_OCEMUXNOT
    );
  MA_15_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(15),
      O => MA_15_OD
    );
  memcontroller_MA_16_OBUF : X_TRI
    port map (
      I => MA_16_OUTMUX,
      CTL => MA_16_ENABLE,
      O => MA(16)
    );
  MA_16_ENABLEINV : X_INV
    port map (
      I => MA_16_TORGTS,
      O => MA_16_ENABLE
    );
  MA_16_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_16_TORGTS
    );
  MA_16_OUTMUX_71 : X_BUF
    port map (
      I => memcontroller_ADDREXT(16),
      O => MA_16_OUTMUX
    );
  MA_16_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MA_16_OCEMUXNOT
    );
  MA_16_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(16),
      O => MA_16_OD
    );
  maccontrol_SOUT_OBUF_72 : X_TRI
    port map (
      I => SOUT_OUTMUX,
      CTL => SOUT_ENABLE,
      O => SOUT
    );
  SOUT_ENABLEINV : X_INV
    port map (
      I => SOUT_TORGTS,
      O => SOUT_ENABLE
    );
  SOUT_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => SOUT_TORGTS
    );
  SOUT_OUTMUX_73 : X_BUF
    port map (
      I => maccontrol_SOUT_OBUF,
      O => SOUT_OUTMUX
    );
  SOUT_OMUX : X_BUF
    port map (
      I => maccontrol_dout(31),
      O => SOUT_OD
    );
  testrx_MACDATA_0_OBUF_74 : X_TRI
    port map (
      I => MACDATA_0_OUTMUX,
      CTL => MACDATA_0_ENABLE,
      O => MACDATA(0)
    );
  MACDATA_0_ENABLEINV : X_INV
    port map (
      I => MACDATA_0_TORGTS,
      O => MACDATA_0_ENABLE
    );
  MACDATA_0_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_0_TORGTS
    );
  MACDATA_0_OUTMUX_75 : X_BUF
    port map (
      I => testrx_MACDATA_0_OBUF,
      O => MACDATA_0_OUTMUX
    );
  MACDATA_0_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(0),
      O => MACDATA_0_OD
    );
  testrx_macaddrl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_MACADDR_1_IBUF,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACADDR_1_IFF_RST,
      O => testrx_macaddrl(1)
    );
  MACADDR_1_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACADDR_1_IFF_RST
    );
  testrx_MACDATA_1_OBUF_76 : X_TRI
    port map (
      I => MACDATA_1_OUTMUX,
      CTL => MACDATA_1_ENABLE,
      O => MACDATA(1)
    );
  MACDATA_1_ENABLEINV : X_INV
    port map (
      I => MACDATA_1_TORGTS,
      O => MACDATA_1_ENABLE
    );
  MACDATA_1_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_1_TORGTS
    );
  MACDATA_1_OUTMUX_77 : X_BUF
    port map (
      I => testrx_MACDATA_1_OBUF,
      O => MACDATA_1_OUTMUX
    );
  MACDATA_1_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(1),
      O => MACDATA_1_OD
    );
  testrx_MACDATA_2_OBUF_78 : X_TRI
    port map (
      I => MACDATA_2_OUTMUX,
      CTL => MACDATA_2_ENABLE,
      O => MACDATA(2)
    );
  MACDATA_2_ENABLEINV : X_INV
    port map (
      I => MACDATA_2_TORGTS,
      O => MACDATA_2_ENABLE
    );
  MACDATA_2_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_2_TORGTS
    );
  MACDATA_2_OUTMUX_79 : X_BUF
    port map (
      I => testrx_MACDATA_2_OBUF,
      O => MACDATA_2_OUTMUX
    );
  MACDATA_2_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(2),
      O => MACDATA_2_OD
    );
  testrx_MACDATA_3_OBUF_80 : X_TRI
    port map (
      I => MACDATA_3_OUTMUX,
      CTL => MACDATA_3_ENABLE,
      O => MACDATA(3)
    );
  MACDATA_3_ENABLEINV : X_INV
    port map (
      I => MACDATA_3_TORGTS,
      O => MACDATA_3_ENABLE
    );
  MACDATA_3_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_3_TORGTS
    );
  MACDATA_3_OUTMUX_81 : X_BUF
    port map (
      I => testrx_MACDATA_3_OBUF,
      O => MACDATA_3_OUTMUX
    );
  MACDATA_3_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(3),
      O => MACDATA_3_OD
    );
  testrx_MACDATA_4_OBUF_82 : X_TRI
    port map (
      I => MACDATA_4_OUTMUX,
      CTL => MACDATA_4_ENABLE,
      O => MACDATA(4)
    );
  MACDATA_4_ENABLEINV : X_INV
    port map (
      I => MACDATA_4_TORGTS,
      O => MACDATA_4_ENABLE
    );
  MACDATA_4_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_4_TORGTS
    );
  MACDATA_4_OUTMUX_83 : X_BUF
    port map (
      I => testrx_MACDATA_4_OBUF,
      O => MACDATA_4_OUTMUX
    );
  MACDATA_4_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(4),
      O => MACDATA_4_OD
    );
  testrx_MACDATA_5_OBUF_84 : X_TRI
    port map (
      I => MACDATA_5_OUTMUX,
      CTL => MACDATA_5_ENABLE,
      O => MACDATA(5)
    );
  MACDATA_5_ENABLEINV : X_INV
    port map (
      I => MACDATA_5_TORGTS,
      O => MACDATA_5_ENABLE
    );
  MACDATA_5_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_5_TORGTS
    );
  MACDATA_5_OUTMUX_85 : X_BUF
    port map (
      I => testrx_MACDATA_5_OBUF,
      O => MACDATA_5_OUTMUX
    );
  MACDATA_5_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(5),
      O => MACDATA_5_OD
    );
  testrx_MACDATA_6_OBUF_86 : X_TRI
    port map (
      I => MACDATA_6_OUTMUX,
      CTL => MACDATA_6_ENABLE,
      O => MACDATA(6)
    );
  MACDATA_6_ENABLEINV : X_INV
    port map (
      I => MACDATA_6_TORGTS,
      O => MACDATA_6_ENABLE
    );
  MACDATA_6_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_6_TORGTS
    );
  MACDATA_6_OUTMUX_87 : X_BUF
    port map (
      I => testrx_MACDATA_6_OBUF,
      O => MACDATA_6_OUTMUX
    );
  MACDATA_6_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(6),
      O => MACDATA_6_OD
    );
  testrx_MACDATA_7_OBUF_88 : X_TRI
    port map (
      I => MACDATA_7_OUTMUX,
      CTL => MACDATA_7_ENABLE,
      O => MACDATA(7)
    );
  MACDATA_7_ENABLEINV : X_INV
    port map (
      I => MACDATA_7_TORGTS,
      O => MACDATA_7_ENABLE
    );
  MACDATA_7_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_7_TORGTS
    );
  MACDATA_7_OUTMUX_89 : X_BUF
    port map (
      I => testrx_MACDATA_7_OBUF,
      O => MACDATA_7_OUTMUX
    );
  MACDATA_7_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(7),
      O => MACDATA_7_OD
    );
  testrx_MACDATA_8_OBUF_90 : X_TRI
    port map (
      I => MACDATA_8_OUTMUX,
      CTL => MACDATA_8_ENABLE,
      O => MACDATA(8)
    );
  MACDATA_8_ENABLEINV : X_INV
    port map (
      I => MACDATA_8_TORGTS,
      O => MACDATA_8_ENABLE
    );
  MACDATA_8_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_8_TORGTS
    );
  MACDATA_8_OUTMUX_91 : X_BUF
    port map (
      I => testrx_MACDATA_8_OBUF,
      O => MACDATA_8_OUTMUX
    );
  MACDATA_8_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(8),
      O => MACDATA_8_OD
    );
  memcontroller_qdout10_OBUFT : X_TRI
    port map (
      I => MD_10_OUTMUX,
      CTL => MD_10_ENABLE,
      O => MD(10)
    );
  MD_10_ENABLEINV : X_INV
    port map (
      I => MD_10_TORGTS,
      O => MD_10_ENABLE
    );
  MD_10_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(10),
      O => MD_10_TORGTS
    );
  MD_10_OUTMUX_92 : X_BUF
    port map (
      I => memcontroller_dnout(10),
      O => MD_10_OUTMUX
    );
  MD_10_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(10),
      O => MD_10_OD
    );
  memcontroller_qdout10_IBUF : X_BUF
    port map (
      I => MD(10),
      O => memcontroller_q(10)
    );
  testrx_macaddrl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_MACADDR_2_IBUF,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACADDR_2_IFF_RST,
      O => testrx_macaddrl(2)
    );
  MACADDR_2_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACADDR_2_IFF_RST
    );
  testrx_MACDATA_9_OBUF_93 : X_TRI
    port map (
      I => MACDATA_9_OUTMUX,
      CTL => MACDATA_9_ENABLE,
      O => MACDATA(9)
    );
  MACDATA_9_ENABLEINV : X_INV
    port map (
      I => MACDATA_9_TORGTS,
      O => MACDATA_9_ENABLE
    );
  MACDATA_9_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_9_TORGTS
    );
  MACDATA_9_OUTMUX_94 : X_BUF
    port map (
      I => testrx_MACDATA_9_OBUF,
      O => MACDATA_9_OUTMUX
    );
  MACDATA_9_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(9),
      O => MACDATA_9_OD
    );
  memcontroller_qdout11_OBUFT : X_TRI
    port map (
      I => MD_11_OUTMUX,
      CTL => MD_11_ENABLE,
      O => MD(11)
    );
  MD_11_ENABLEINV : X_INV
    port map (
      I => MD_11_TORGTS,
      O => MD_11_ENABLE
    );
  MD_11_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(11),
      O => MD_11_TORGTS
    );
  MD_11_OUTMUX_95 : X_BUF
    port map (
      I => memcontroller_dnout(11),
      O => MD_11_OUTMUX
    );
  MD_11_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(11),
      O => MD_11_OD
    );
  memcontroller_qdout11_IBUF : X_BUF
    port map (
      I => MD(11),
      O => memcontroller_q(11)
    );
  memcontroller_qdout20_OBUFT : X_TRI
    port map (
      I => MD_20_OUTMUX,
      CTL => MD_20_ENABLE,
      O => MD(20)
    );
  MD_20_ENABLEINV : X_INV
    port map (
      I => MD_20_TORGTS,
      O => MD_20_ENABLE
    );
  MD_20_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(20),
      O => MD_20_TORGTS
    );
  MD_20_OUTMUX_96 : X_BUF
    port map (
      I => memcontroller_dnout(20),
      O => MD_20_OUTMUX
    );
  MD_20_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(20),
      O => MD_20_OD
    );
  memcontroller_qdout20_IBUF : X_BUF
    port map (
      I => MD(20),
      O => memcontroller_q(20)
    );
  memcontroller_qdout12_OBUFT : X_TRI
    port map (
      I => MD_12_OUTMUX,
      CTL => MD_12_ENABLE,
      O => MD(12)
    );
  MD_12_ENABLEINV : X_INV
    port map (
      I => MD_12_TORGTS,
      O => MD_12_ENABLE
    );
  MD_12_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(12),
      O => MD_12_TORGTS
    );
  MD_12_OUTMUX_97 : X_BUF
    port map (
      I => memcontroller_dnout(12),
      O => MD_12_OUTMUX
    );
  MD_12_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(12),
      O => MD_12_OD
    );
  memcontroller_qdout12_IBUF : X_BUF
    port map (
      I => MD(12),
      O => memcontroller_q(12)
    );
  memcontroller_qdout21_OBUFT : X_TRI
    port map (
      I => MD_21_OUTMUX,
      CTL => MD_21_ENABLE,
      O => MD(21)
    );
  MD_21_ENABLEINV : X_INV
    port map (
      I => MD_21_TORGTS,
      O => MD_21_ENABLE
    );
  MD_21_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(21),
      O => MD_21_TORGTS
    );
  MD_21_OUTMUX_98 : X_BUF
    port map (
      I => memcontroller_dnout(21),
      O => MD_21_OUTMUX
    );
  MD_21_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(21),
      O => MD_21_OD
    );
  memcontroller_qdout21_IBUF : X_BUF
    port map (
      I => MD(21),
      O => memcontroller_q(21)
    );
  memcontroller_qdout13_OBUFT : X_TRI
    port map (
      I => MD_13_OUTMUX,
      CTL => MD_13_ENABLE,
      O => MD(13)
    );
  MD_13_ENABLEINV : X_INV
    port map (
      I => MD_13_TORGTS,
      O => MD_13_ENABLE
    );
  MD_13_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(13),
      O => MD_13_TORGTS
    );
  MD_13_OUTMUX_99 : X_BUF
    port map (
      I => memcontroller_dnout(13),
      O => MD_13_OUTMUX
    );
  MD_13_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(13),
      O => MD_13_OD
    );
  memcontroller_qdout13_IBUF : X_BUF
    port map (
      I => MD(13),
      O => memcontroller_q(13)
    );
  memcontroller_qdout22_OBUFT : X_TRI
    port map (
      I => MD_22_OUTMUX,
      CTL => MD_22_ENABLE,
      O => MD(22)
    );
  MD_22_ENABLEINV : X_INV
    port map (
      I => MD_22_TORGTS,
      O => MD_22_ENABLE
    );
  MD_22_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(22),
      O => MD_22_TORGTS
    );
  MD_22_OUTMUX_100 : X_BUF
    port map (
      I => memcontroller_dnout(22),
      O => MD_22_OUTMUX
    );
  MD_22_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(22),
      O => MD_22_OD
    );
  memcontroller_qdout22_IBUF : X_BUF
    port map (
      I => MD(22),
      O => memcontroller_q(22)
    );
  memcontroller_qdout14_OBUFT : X_TRI
    port map (
      I => MD_14_OUTMUX,
      CTL => MD_14_ENABLE,
      O => MD(14)
    );
  MD_14_ENABLEINV : X_INV
    port map (
      I => MD_14_TORGTS,
      O => MD_14_ENABLE
    );
  MD_14_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(14),
      O => MD_14_TORGTS
    );
  MD_14_OUTMUX_101 : X_BUF
    port map (
      I => memcontroller_dnout(14),
      O => MD_14_OUTMUX
    );
  MD_14_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(14),
      O => MD_14_OD
    );
  memcontroller_qdout14_IBUF : X_BUF
    port map (
      I => MD(14),
      O => memcontroller_q(14)
    );
  memcontroller_qdout30_OBUFT : X_TRI
    port map (
      I => MD_30_OUTMUX,
      CTL => MD_30_ENABLE,
      O => MD(30)
    );
  MD_30_ENABLEINV : X_INV
    port map (
      I => MD_30_TORGTS,
      O => MD_30_ENABLE
    );
  MD_30_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(30),
      O => MD_30_TORGTS
    );
  MD_30_OUTMUX_102 : X_BUF
    port map (
      I => memcontroller_dnout(30),
      O => MD_30_OUTMUX
    );
  MD_30_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(30),
      O => MD_30_OD
    );
  memcontroller_qdout30_IBUF : X_BUF
    port map (
      I => MD(30),
      O => memcontroller_q(30)
    );
  testrx_macaddrl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_MACADDR_3_IBUF,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACADDR_3_IFF_RST,
      O => testrx_macaddrl(3)
    );
  MACADDR_3_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACADDR_3_IFF_RST
    );
  memcontroller_qdout23_OBUFT : X_TRI
    port map (
      I => MD_23_OUTMUX,
      CTL => MD_23_ENABLE,
      O => MD(23)
    );
  MD_23_ENABLEINV : X_INV
    port map (
      I => MD_23_TORGTS,
      O => MD_23_ENABLE
    );
  MD_23_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(23),
      O => MD_23_TORGTS
    );
  MD_23_OUTMUX_103 : X_BUF
    port map (
      I => memcontroller_dnout(23),
      O => MD_23_OUTMUX
    );
  MD_23_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(23),
      O => MD_23_OD
    );
  memcontroller_qdout23_IBUF : X_BUF
    port map (
      I => MD(23),
      O => memcontroller_q(23)
    );
  memcontroller_qdout15_OBUFT : X_TRI
    port map (
      I => MD_15_OUTMUX,
      CTL => MD_15_ENABLE,
      O => MD(15)
    );
  MD_15_ENABLEINV : X_INV
    port map (
      I => MD_15_TORGTS,
      O => MD_15_ENABLE
    );
  MD_15_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(15),
      O => MD_15_TORGTS
    );
  MD_15_OUTMUX_104 : X_BUF
    port map (
      I => memcontroller_dnout(15),
      O => MD_15_OUTMUX
    );
  MD_15_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(15),
      O => MD_15_OD
    );
  memcontroller_qdout15_IBUF : X_BUF
    port map (
      I => MD(15),
      O => memcontroller_q(15)
    );
  memcontroller_qdout31_OBUFT : X_TRI
    port map (
      I => MD_31_OUTMUX,
      CTL => MD_31_ENABLE,
      O => MD(31)
    );
  MD_31_ENABLEINV : X_INV
    port map (
      I => MD_31_TORGTS,
      O => MD_31_ENABLE
    );
  MD_31_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(31),
      O => MD_31_TORGTS
    );
  MD_31_OUTMUX_105 : X_BUF
    port map (
      I => memcontroller_dnout(31),
      O => MD_31_OUTMUX
    );
  MD_31_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(31),
      O => MD_31_OD
    );
  memcontroller_qdout31_IBUF : X_BUF
    port map (
      I => MD(31),
      O => memcontroller_q(31)
    );
  memcontroller_qdout24_OBUFT : X_TRI
    port map (
      I => MD_24_OUTMUX,
      CTL => MD_24_ENABLE,
      O => MD(24)
    );
  MD_24_ENABLEINV : X_INV
    port map (
      I => MD_24_TORGTS,
      O => MD_24_ENABLE
    );
  MD_24_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(24),
      O => MD_24_TORGTS
    );
  MD_24_OUTMUX_106 : X_BUF
    port map (
      I => memcontroller_dnout(24),
      O => MD_24_OUTMUX
    );
  MD_24_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(24),
      O => MD_24_OD
    );
  memcontroller_qdout24_IBUF : X_BUF
    port map (
      I => MD(24),
      O => memcontroller_q(24)
    );
  memcontroller_qdout16_OBUFT : X_TRI
    port map (
      I => MD_16_OUTMUX,
      CTL => MD_16_ENABLE,
      O => MD(16)
    );
  MD_16_ENABLEINV : X_INV
    port map (
      I => MD_16_TORGTS,
      O => MD_16_ENABLE
    );
  MD_16_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(16),
      O => MD_16_TORGTS
    );
  MD_16_OUTMUX_107 : X_BUF
    port map (
      I => memcontroller_dnout(16),
      O => MD_16_OUTMUX
    );
  MD_16_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(16),
      O => MD_16_OD
    );
  memcontroller_qdout16_IBUF : X_BUF
    port map (
      I => MD(16),
      O => memcontroller_q(16)
    );
  memcontroller_qdout17_OBUFT : X_TRI
    port map (
      I => MD_17_OUTMUX,
      CTL => MD_17_ENABLE,
      O => MD(17)
    );
  MD_17_ENABLEINV : X_INV
    port map (
      I => MD_17_TORGTS,
      O => MD_17_ENABLE
    );
  MD_17_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(17),
      O => MD_17_TORGTS
    );
  MD_17_OUTMUX_108 : X_BUF
    port map (
      I => memcontroller_dnout(17),
      O => MD_17_OUTMUX
    );
  MD_17_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(17),
      O => MD_17_OD
    );
  memcontroller_qdout17_IBUF : X_BUF
    port map (
      I => MD(17),
      O => memcontroller_q(17)
    );
  memcontroller_qdout25_OBUFT : X_TRI
    port map (
      I => MD_25_OUTMUX,
      CTL => MD_25_ENABLE,
      O => MD(25)
    );
  MD_25_ENABLEINV : X_INV
    port map (
      I => MD_25_TORGTS,
      O => MD_25_ENABLE
    );
  MD_25_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(25),
      O => MD_25_TORGTS
    );
  MD_25_OUTMUX_109 : X_BUF
    port map (
      I => memcontroller_dnout(25),
      O => MD_25_OUTMUX
    );
  MD_25_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(25),
      O => MD_25_OD
    );
  memcontroller_qdout25_IBUF : X_BUF
    port map (
      I => MD(25),
      O => memcontroller_q(25)
    );
  memcontroller_qdout18_OBUFT : X_TRI
    port map (
      I => MD_18_OUTMUX,
      CTL => MD_18_ENABLE,
      O => MD(18)
    );
  MD_18_ENABLEINV : X_INV
    port map (
      I => MD_18_TORGTS,
      O => MD_18_ENABLE
    );
  MD_18_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(18),
      O => MD_18_TORGTS
    );
  MD_18_OUTMUX_110 : X_BUF
    port map (
      I => memcontroller_dnout(18),
      O => MD_18_OUTMUX
    );
  MD_18_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(18),
      O => MD_18_OD
    );
  memcontroller_qdout18_IBUF : X_BUF
    port map (
      I => MD(18),
      O => memcontroller_q(18)
    );
  memcontroller_qdout26_OBUFT : X_TRI
    port map (
      I => MD_26_OUTMUX,
      CTL => MD_26_ENABLE,
      O => MD(26)
    );
  MD_26_ENABLEINV : X_INV
    port map (
      I => MD_26_TORGTS,
      O => MD_26_ENABLE
    );
  MD_26_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(26),
      O => MD_26_TORGTS
    );
  MD_26_OUTMUX_111 : X_BUF
    port map (
      I => memcontroller_dnout(26),
      O => MD_26_OUTMUX
    );
  MD_26_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(26),
      O => MD_26_OD
    );
  memcontroller_qdout26_IBUF : X_BUF
    port map (
      I => MD(26),
      O => memcontroller_q(26)
    );
  testrx_macaddrl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_MACADDR_4_IBUF,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACADDR_4_IFF_RST,
      O => testrx_macaddrl(4)
    );
  MACADDR_4_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACADDR_4_IFF_RST
    );
  memcontroller_qdout19_OBUFT : X_TRI
    port map (
      I => MD_19_OUTMUX,
      CTL => MD_19_ENABLE,
      O => MD(19)
    );
  MD_19_ENABLEINV : X_INV
    port map (
      I => MD_19_TORGTS,
      O => MD_19_ENABLE
    );
  MD_19_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(19),
      O => MD_19_TORGTS
    );
  MD_19_OUTMUX_112 : X_BUF
    port map (
      I => memcontroller_dnout(19),
      O => MD_19_OUTMUX
    );
  MD_19_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(19),
      O => MD_19_OD
    );
  memcontroller_qdout19_IBUF : X_BUF
    port map (
      I => MD(19),
      O => memcontroller_q(19)
    );
  memcontroller_qdout27_OBUFT : X_TRI
    port map (
      I => MD_27_OUTMUX,
      CTL => MD_27_ENABLE,
      O => MD(27)
    );
  MD_27_ENABLEINV : X_INV
    port map (
      I => MD_27_TORGTS,
      O => MD_27_ENABLE
    );
  MD_27_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(27),
      O => MD_27_TORGTS
    );
  MD_27_OUTMUX_113 : X_BUF
    port map (
      I => memcontroller_dnout(27),
      O => MD_27_OUTMUX
    );
  MD_27_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(27),
      O => MD_27_OD
    );
  memcontroller_qdout27_IBUF : X_BUF
    port map (
      I => MD(27),
      O => memcontroller_q(27)
    );
  maccontrol_PHYRESET_OBUF_114 : X_TRI
    port map (
      I => PHYRESET_OUTMUX,
      CTL => PHYRESET_ENABLE,
      O => PHYRESET
    );
  PHYRESET_ENABLEINV : X_INV
    port map (
      I => PHYRESET_TORGTS,
      O => PHYRESET_ENABLE
    );
  PHYRESET_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => PHYRESET_TORGTS
    );
  PHYRESET_OUTMUX_115 : X_BUF
    port map (
      I => maccontrol_PHYRESET_OBUF,
      O => PHYRESET_OUTMUX
    );
  PHYRESET_OMUX : X_BUF
    port map (
      I => maccontrol_n0041,
      O => PHYRESET_OD
    );
  memcontroller_qdout28_OBUFT : X_TRI
    port map (
      I => MD_28_OUTMUX,
      CTL => MD_28_ENABLE,
      O => MD(28)
    );
  MD_28_ENABLEINV : X_INV
    port map (
      I => MD_28_TORGTS,
      O => MD_28_ENABLE
    );
  MD_28_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(28),
      O => MD_28_TORGTS
    );
  MD_28_OUTMUX_116 : X_BUF
    port map (
      I => memcontroller_dnout(28),
      O => MD_28_OUTMUX
    );
  MD_28_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(28),
      O => MD_28_OD
    );
  memcontroller_qdout28_IBUF : X_BUF
    port map (
      I => MD(28),
      O => memcontroller_q(28)
    );
  memcontroller_qdout29_OBUFT : X_TRI
    port map (
      I => MD_29_OUTMUX,
      CTL => MD_29_ENABLE,
      O => MD(29)
    );
  MD_29_ENABLEINV : X_INV
    port map (
      I => MD_29_TORGTS,
      O => MD_29_ENABLE
    );
  MD_29_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(29),
      O => MD_29_TORGTS
    );
  MD_29_OUTMUX_117 : X_BUF
    port map (
      I => memcontroller_dnout(29),
      O => MD_29_OUTMUX
    );
  MD_29_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(29),
      O => MD_29_OD
    );
  memcontroller_qdout29_IBUF : X_BUF
    port map (
      I => MD(29),
      O => memcontroller_q(29)
    );
  maccontrol_LED100_OBUF_118 : X_TRI
    port map (
      I => LED100_OUTMUX,
      CTL => LED100_ENABLE,
      O => LED100
    );
  LED100_ENABLEINV : X_INV
    port map (
      I => LED100_TORGTS,
      O => LED100_ENABLE
    );
  LED100_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LED100_TORGTS
    );
  LED100_OUTMUX_119 : X_BUF
    port map (
      I => maccontrol_LED100_OBUF,
      O => LED100_OUTMUX
    );
  LED100_OMUX : X_BUF
    port map (
      I => maccontrol_n0043,
      O => LED100_OD
    );
  NEXTF_IMUX : X_BUF
    port map (
      I => NEXTF_IBUF_0,
      O => NEXTF_IBUF
    );
  NEXTF_IBUF_120 : X_BUF
    port map (
      I => NEXTF,
      O => NEXTF_IBUF_0
    );
  RESET_IMUX : X_BUF
    port map (
      I => RESET_IBUF_1,
      O => RESET_IBUF
    );
  RESET_IBUF_121 : X_BUF
    port map (
      I => RESET,
      O => RESET_IBUF_1
    );
  maccontrol_PHY_status_MII_Interface_iobuffer_OBUFT : X_TRI
    port map (
      I => MDIO_OUTMUX,
      CTL => MDIO_ENABLE,
      O => MDIO
    );
  MDIO_ENABLEINV : X_INV
    port map (
      I => MDIO_TORGTS,
      O => MDIO_ENABLE
    );
  MDIO_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => maccontrol_PHY_status_MII_Interface_sts,
      O => MDIO_TORGTS
    );
  MDIO_OUTMUX_122 : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_sout,
      O => MDIO_OUTMUX
    );
  maccontrol_PHY_status_MII_Interface_iobuffer_IBUF : X_BUF
    port map (
      I => MDIO,
      O => maccontrol_PHY_status_MII_Interface_sin
    );
  testrx_macaddrl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_MACADDR_5_IBUF,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACADDR_5_IFF_RST,
      O => testrx_macaddrl(5)
    );
  MACADDR_5_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACADDR_5_IFF_RST
    );
  MDC_OBUF_123 : X_TRI
    port map (
      I => MDC_OUTMUX,
      CTL => MDC_ENABLE,
      O => MDC
    );
  MDC_ENABLEINV : X_INV
    port map (
      I => MDC_TORGTS,
      O => MDC_ENABLE
    );
  MDC_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MDC_TORGTS
    );
  MDC_OUTMUX_124 : X_BUF
    port map (
      I => MDC_OBUF,
      O => MDC_OUTMUX
    );
  MOE_LOGIC_ZERO_125 : X_ZERO
    port map (
      O => MOE_LOGIC_ZERO
    );
  MOE_OBUF : X_TRI
    port map (
      I => MOE_OUTMUX,
      CTL => MOE_ENABLE,
      O => MOE
    );
  MOE_ENABLEINV : X_INV
    port map (
      I => MOE_TORGTS,
      O => MOE_ENABLE
    );
  MOE_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MOE_TORGTS
    );
  MOE_OUTMUX_126 : X_BUF
    port map (
      I => MOE_LOGIC_ZERO,
      O => MOE_OUTMUX
    );
  testrx_RXD_0_IBUF_127 : X_BUF
    port map (
      I => RXD(0),
      O => testrx_RXD_0_IBUF
    );
  testrx_RXD_1_IBUF_128 : X_BUF
    port map (
      I => RXD(1),
      O => testrx_RXD_1_IBUF
    );
  testrx_RXD_2_IBUF_129 : X_BUF
    port map (
      I => RXD(2),
      O => testrx_RXD_2_IBUF
    );
  testrx_RXD_3_IBUF_130 : X_BUF
    port map (
      I => RXD(3),
      O => testrx_RXD_3_IBUF
    );
  testrx_RXD_4_IBUF_131 : X_BUF
    port map (
      I => RXD(4),
      O => testrx_RXD_4_IBUF
    );
  testrx_RXD_5_IBUF_132 : X_BUF
    port map (
      I => RXD(5),
      O => testrx_RXD_5_IBUF
    );
  memcontroller_MWE_OBUF : X_TRI
    port map (
      I => MWE_OUTMUX,
      CTL => MWE_ENABLE,
      O => MWE
    );
  MWE_ENABLEINV : X_INV
    port map (
      I => MWE_TORGTS,
      O => MWE_ENABLE
    );
  MWE_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MWE_TORGTS
    );
  MWE_OUTMUX_133 : X_BUF
    port map (
      I => memcontroller_WEEXT,
      O => MWE_OUTMUX
    );
  MWE_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MWE_OCEMUXNOT
    );
  MWE_OMUX : X_BUF
    port map (
      I => memcontroller_n0116,
      O => MWE_OD
    );
  testrx_macaddrl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_MACADDR_6_IBUF,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACADDR_6_IFF_RST,
      O => testrx_macaddrl(6)
    );
  MACADDR_6_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACADDR_6_IFF_RST
    );
  testrx_RXD_6_IBUF_134 : X_BUF
    port map (
      I => RXD(6),
      O => testrx_RXD_6_IBUF
    );
  SCS_IMUX : X_BUF
    port map (
      I => SCS_IBUF_2,
      O => SCS_IBUF
    );
  SCS_IBUF_135 : X_BUF
    port map (
      I => SCS,
      O => SCS_IBUF_2
    );
  testrx_RXD_7_IBUF_136 : X_BUF
    port map (
      I => RXD(7),
      O => testrx_RXD_7_IBUF
    );
  SIN_IMUX : X_BUF
    port map (
      I => SIN_IBUF_3,
      O => SIN_IBUF
    );
  SIN_IBUF_137 : X_BUF
    port map (
      I => SIN,
      O => SIN_IBUF_3
    );
  maccontrol_LED1000_OBUF_138 : X_TRI
    port map (
      I => LED1000_OUTMUX,
      CTL => LED1000_ENABLE,
      O => LED1000
    );
  LED1000_ENABLEINV : X_INV
    port map (
      I => LED1000_TORGTS,
      O => LED1000_ENABLE
    );
  LED1000_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LED1000_TORGTS
    );
  LED1000_OUTMUX_139 : X_BUF
    port map (
      I => maccontrol_LED1000_OBUF,
      O => LED1000_OUTMUX
    );
  LED1000_OMUX : X_BUF
    port map (
      I => maccontrol_n0042,
      O => LED1000_OD
    );
  RX_ER_IMUX : X_BUF
    port map (
      I => RX_ER_IBUF_4,
      O => RX_ER_IBUF
    );
  RX_ER_IBUF_140 : X_BUF
    port map (
      I => RX_ER,
      O => RX_ER_IBUF_4
    );
  RX_DV_IMUX : X_BUF
    port map (
      I => RX_DV_IBUF_5,
      O => RX_DV_IBUF
    );
  RX_DV_IBUF_141 : X_BUF
    port map (
      I => RX_DV,
      O => RX_DV_IBUF_5
    );
  testrx_MACDATA_10_OBUF_142 : X_TRI
    port map (
      I => MACDATA_10_OUTMUX,
      CTL => MACDATA_10_ENABLE,
      O => MACDATA(10)
    );
  MACDATA_10_ENABLEINV : X_INV
    port map (
      I => MACDATA_10_TORGTS,
      O => MACDATA_10_ENABLE
    );
  MACDATA_10_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_10_TORGTS
    );
  MACDATA_10_OUTMUX_143 : X_BUF
    port map (
      I => testrx_MACDATA_10_OBUF,
      O => MACDATA_10_OUTMUX
    );
  MACDATA_10_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(10),
      O => MACDATA_10_OD
    );
  testrx_MACDATA_11_OBUF_144 : X_TRI
    port map (
      I => MACDATA_11_OUTMUX,
      CTL => MACDATA_11_ENABLE,
      O => MACDATA(11)
    );
  MACDATA_11_ENABLEINV : X_INV
    port map (
      I => MACDATA_11_TORGTS,
      O => MACDATA_11_ENABLE
    );
  MACDATA_11_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_11_TORGTS
    );
  MACDATA_11_OUTMUX_145 : X_BUF
    port map (
      I => testrx_MACDATA_11_OBUF,
      O => MACDATA_11_OUTMUX
    );
  MACDATA_11_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(11),
      O => MACDATA_11_OD
    );
  testrx_macaddrl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_MACADDR_7_IBUF,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACADDR_7_IFF_RST,
      O => testrx_macaddrl(7)
    );
  MACADDR_7_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACADDR_7_IFF_RST
    );
  testrx_MACDATA_12_OBUF_146 : X_TRI
    port map (
      I => MACDATA_12_OUTMUX,
      CTL => MACDATA_12_ENABLE,
      O => MACDATA(12)
    );
  MACDATA_12_ENABLEINV : X_INV
    port map (
      I => MACDATA_12_TORGTS,
      O => MACDATA_12_ENABLE
    );
  MACDATA_12_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_12_TORGTS
    );
  MACDATA_12_OUTMUX_147 : X_BUF
    port map (
      I => testrx_MACDATA_12_OBUF,
      O => MACDATA_12_OUTMUX
    );
  MACDATA_12_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(12),
      O => MACDATA_12_OD
    );
  testrx_MACDATA_13_OBUF_148 : X_TRI
    port map (
      I => MACDATA_13_OUTMUX,
      CTL => MACDATA_13_ENABLE,
      O => MACDATA(13)
    );
  MACDATA_13_ENABLEINV : X_INV
    port map (
      I => MACDATA_13_TORGTS,
      O => MACDATA_13_ENABLE
    );
  MACDATA_13_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_13_TORGTS
    );
  MACDATA_13_OUTMUX_149 : X_BUF
    port map (
      I => testrx_MACDATA_13_OBUF,
      O => MACDATA_13_OUTMUX
    );
  MACDATA_13_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(13),
      O => MACDATA_13_OD
    );
  TX_ER_LOGIC_ZERO_150 : X_ZERO
    port map (
      O => TX_ER_LOGIC_ZERO
    );
  TX_ER_OBUF : X_TRI
    port map (
      I => TX_ER_OUTMUX,
      CTL => TX_ER_ENABLE,
      O => TX_ER
    );
  TX_ER_ENABLEINV : X_INV
    port map (
      I => TX_ER_TORGTS,
      O => TX_ER_ENABLE
    );
  TX_ER_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TX_ER_TORGTS
    );
  TX_ER_OUTMUX_151 : X_BUF
    port map (
      I => TX_ER_LOGIC_ZERO,
      O => TX_ER_OUTMUX
    );
  testrx_MACDATA_14_OBUF_152 : X_TRI
    port map (
      I => MACDATA_14_OUTMUX,
      CTL => MACDATA_14_ENABLE,
      O => MACDATA(14)
    );
  MACDATA_14_ENABLEINV : X_INV
    port map (
      I => MACDATA_14_TORGTS,
      O => MACDATA_14_ENABLE
    );
  MACDATA_14_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_14_TORGTS
    );
  MACDATA_14_OUTMUX_153 : X_BUF
    port map (
      I => testrx_MACDATA_14_OBUF,
      O => MACDATA_14_OUTMUX
    );
  MACDATA_14_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(14),
      O => MACDATA_14_OD
    );
  testrx_MACDATA_15_OBUF_154 : X_TRI
    port map (
      I => MACDATA_15_OUTMUX,
      CTL => MACDATA_15_ENABLE,
      O => MACDATA(15)
    );
  MACDATA_15_ENABLEINV : X_INV
    port map (
      I => MACDATA_15_TORGTS,
      O => MACDATA_15_ENABLE
    );
  MACDATA_15_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MACDATA_15_TORGTS
    );
  MACDATA_15_OUTMUX_155 : X_BUF
    port map (
      I => testrx_MACDATA_15_OBUF,
      O => MACDATA_15_OUTMUX
    );
  MACDATA_15_OMUX : X_BUF
    port map (
      I => testrx_lmacdata(15),
      O => MACDATA_15_OD
    );
  GTX_CLK_OBUF_156 : X_TRI
    port map (
      I => GTX_CLK_OUTMUX,
      CTL => GTX_CLK_ENABLE,
      O => GTX_CLK
    );
  GTX_CLK_ENABLEINV : X_INV
    port map (
      I => GTX_CLK_TORGTS,
      O => GTX_CLK_ENABLE
    );
  GTX_CLK_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => GTX_CLK_TORGTS
    );
  GTX_CLK_OUTMUX_157 : X_BUF
    port map (
      I => GTX_CLK_OBUF,
      O => GTX_CLK_OUTMUX
    );
  maccontrol_LEDTX_OBUF_158 : X_TRI
    port map (
      I => LEDTX_OUTMUX,
      CTL => LEDTX_ENABLE,
      O => LEDTX
    );
  LEDTX_ENABLEINV : X_INV
    port map (
      I => LEDTX_TORGTS,
      O => LEDTX_ENABLE
    );
  LEDTX_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDTX_TORGTS
    );
  LEDTX_OUTMUX_159 : X_BUF
    port map (
      I => maccontrol_LEDTX_OBUF,
      O => LEDTX_OUTMUX
    );
  LEDTX_OMUX : X_BUF
    port map (
      I => maccontrol_n0045,
      O => LEDTX_OD
    );
  LEDPOWER_OBUF_160 : X_TRI
    port map (
      I => LEDPOWER_OUTMUX,
      CTL => LEDPOWER_ENABLE,
      O => LEDPOWER
    );
  LEDPOWER_ENABLEINV : X_INV
    port map (
      I => LEDPOWER_TORGTS,
      O => LEDPOWER_ENABLE
    );
  LEDPOWER_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDPOWER_TORGTS
    );
  LEDPOWER_OUTMUX_161 : X_BUF
    port map (
      I => LEDPOWER_OBUF,
      O => LEDPOWER_OUTMUX
    );
  LEDPOWER_OMUX : X_BUF
    port map (
      I => Q_n0000(23),
      O => LEDPOWER_OD
    );
  ifclk_DLL : X_CLKDLLE
    generic map(
      CLKDV_DIVIDE => 4.0,
      DUTY_CYCLE_CORRECTION => TRUE,
      MAXPERCLKIN => 40000 ps
    )
    port map (
      CLKIN => IFCLK_IBUFG,
      CLKFB => ifclk_int,
      RST => RESET_IBUF,
      CLK0 => ifclk_to_bufg,
      CLK90 => ifclk_DLL_CLK90,
      CLK180 => ifclk_DLL_CLK180,
      CLK270 => ifclk_DLL_CLK270,
      CLK2X => ifclk_DLL_CLK2X,
      CLK2X180 => ifclk_DLL_CLK2X180,
      CLKDV => ifclk_DLL_CLKDV,
      LOCKED => ifclk_DLL_LOCKED
    );
  clk_DLL : X_CLKDLLE
    generic map(
      CLKDV_DIVIDE => 4.0,
      DUTY_CYCLE_CORRECTION => TRUE,
      MAXPERCLKIN => 40000 ps
    )
    port map (
      CLKIN => CLKIN_IBUFG,
      CLKFB => CLKFB_IBUFG,
      RST => RESET_IBUF,
      CLK0 => clk_to_bufg,
      CLK90 => MCLK_OBUF,
      CLK180 => GTX_CLK_OBUF,
      CLK270 => clk_DLL_CLK270,
      CLK2X => clk_DLL_CLK2X,
      CLK2X180 => clk_DLL_CLK2X180,
      CLKDV => clk_DLL_CLKDV,
      LOCKED => clk_DLL_LOCKED
    );
  rxclk_DLL : X_CLKDLLE
    generic map(
      CLKDV_DIVIDE => 4.0,
      DUTY_CYCLE_CORRECTION => TRUE,
      MAXPERCLKIN => 40000 ps
    )
    port map (
      CLKIN => RX_CLK_IBUFG,
      CLKFB => rx_clk_int,
      RST => NEXTF_IBUF,
      CLK0 => rx_clk_to_bufg,
      CLK90 => rxclk_DLL_CLK90,
      CLK180 => rxclk_DLL_CLK180,
      CLK270 => rxclk_DLL_CLK270,
      CLK2X => rxclk_DLL_CLK2X,
      CLK2X180 => rxclk_DLL_CLK2X180,
      CLKDV => rxclk_DLL_CLKDV,
      LOCKED => rxclk_DLL_LOCKED
    );
  testrx_tempram_LOGIC_ZERO_162 : X_ZERO
    port map (
      O => testrx_tempram_LOGIC_ZERO
    );
  testrx_tempram_LOGIC_ONE_163 : X_ONE
    port map (
      O => testrx_tempram_LOGIC_ONE
    );
  testrx_tempram : X_RAMB4_S8_S16
    generic map(
      INIT_00 => X"00000000000000000000000000000000000000000000000000FEDCBA87654321",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      SETUP_ALL => 3025 ps,
      XON => FALSE
    )
    port map (
      CLKA => rx_clk_int,
      CLKB => ifclk_int,
      ENA => testrx_tempram_LOGIC_ONE,
      ENB => testrx_tempram_LOGIC_ONE,
      RSTA => RESET_IBUF,
      RSTB => RESET_IBUF,
      WEA => testrx_cs_FFd2,
      WEB => testrx_tempram_LOGIC_ZERO,
      GSR => GSR,
      ADDRA(8) => GLOBAL_LOGIC0_64,
      ADDRA(7) => testrx_addr(7),
      ADDRA(6) => testrx_addr(6),
      ADDRA(5) => testrx_addr(5),
      ADDRA(4) => testrx_addr(4),
      ADDRA(3) => testrx_addr(3),
      ADDRA(2) => testrx_addr(2),
      ADDRA(1) => testrx_addr(1),
      ADDRA(0) => testrx_addr(0),
      ADDRB(7) => testrx_macaddrl(7),
      ADDRB(6) => testrx_macaddrl(6),
      ADDRB(5) => testrx_macaddrl(5),
      ADDRB(4) => testrx_macaddrl(4),
      ADDRB(3) => testrx_macaddrl(3),
      ADDRB(2) => testrx_macaddrl(2),
      ADDRB(1) => testrx_macaddrl(1),
      ADDRB(0) => testrx_macaddrl(0),
      DIA(7) => testrx_rxdll(7),
      DIA(6) => testrx_rxdll(6),
      DIA(5) => testrx_rxdll(5),
      DIA(4) => testrx_rxdll(4),
      DIA(3) => testrx_rxdll(3),
      DIA(2) => testrx_rxdll(2),
      DIA(1) => testrx_rxdll(1),
      DIA(0) => testrx_rxdll(0),
      DIB(15) => GLOBAL_LOGIC0_64,
      DIB(14) => GLOBAL_LOGIC0_64,
      DIB(13) => GLOBAL_LOGIC0_64,
      DIB(12) => GLOBAL_LOGIC0_64,
      DIB(11) => GLOBAL_LOGIC0_65,
      DIB(10) => GLOBAL_LOGIC0_64,
      DIB(9) => GLOBAL_LOGIC0_65,
      DIB(8) => GLOBAL_LOGIC0_64,
      DIB(7) => GLOBAL_LOGIC0_64,
      DIB(6) => GLOBAL_LOGIC0_64,
      DIB(5) => GLOBAL_LOGIC0_64,
      DIB(4) => GLOBAL_LOGIC0_64,
      DIB(3) => GLOBAL_LOGIC0_66,
      DIB(2) => GLOBAL_LOGIC0_64,
      DIB(1) => GLOBAL_LOGIC0_65,
      DIB(0) => GLOBAL_LOGIC0_64,
      DOA(7) => testrx_tempram_DOA7,
      DOA(6) => testrx_tempram_DOA6,
      DOA(5) => testrx_tempram_DOA5,
      DOA(4) => testrx_tempram_DOA4,
      DOA(3) => testrx_tempram_DOA3,
      DOA(2) => testrx_tempram_DOA2,
      DOA(1) => testrx_tempram_DOA1,
      DOA(0) => testrx_tempram_DOA0,
      DOB(15) => testrx_lmacdata(15),
      DOB(14) => testrx_lmacdata(14),
      DOB(13) => testrx_lmacdata(13),
      DOB(12) => testrx_lmacdata(12),
      DOB(11) => testrx_lmacdata(11),
      DOB(10) => testrx_lmacdata(10),
      DOB(9) => testrx_lmacdata(9),
      DOB(8) => testrx_lmacdata(8),
      DOB(7) => testrx_lmacdata(7),
      DOB(6) => testrx_lmacdata(6),
      DOB(5) => testrx_lmacdata(5),
      DOB(4) => testrx_lmacdata(4),
      DOB(3) => testrx_lmacdata(3),
      DOB(2) => testrx_lmacdata(2),
      DOB(1) => testrx_lmacdata(1),
      DOB(0) => testrx_lmacdata(0)
    );
  txsim_rom_LOGIC_ZERO_164 : X_ZERO
    port map (
      O => txsim_rom_LOGIC_ZERO
    );
  txsim_rom_LOGIC_ONE_165 : X_ONE
    port map (
      O => txsim_rom_LOGIC_ONE
    );
  txsim_rom : X_RAMB4_S8
    generic map(
      INIT_00 => X"B8014000400000540000450008E38B18E90700FFFFFFFFFFFFD5555555555555",
      INIT_01 => X"0E0D0C0B0A0908000756AF3FB2A2791D2048265EE40008FF00A8C00100A8C058",
      INIT_02 => X"2E2D2C2B2A292827262524232221201F1E1D1C1B1A191817161514131211100F",
      INIT_03 => X"00000000000000000000000000000000000000B26BD4D437363534333231302F",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      XON => FALSE
    )
    port map (
      CLK => clk,
      EN => txsim_rom_LOGIC_ONE,
      RST => RESET_IBUF,
      WE => txsim_rom_LOGIC_ZERO,
      GSR => GSR,
      ADDR(8) => txsim_counter(8),
      ADDR(7) => txsim_counter(7),
      ADDR(6) => txsim_counter(6),
      ADDR(5) => txsim_counter(5),
      ADDR(4) => txsim_counter(4),
      ADDR(3) => txsim_counter(3),
      ADDR(2) => txsim_counter(2),
      ADDR(1) => txsim_counter(1),
      ADDR(0) => txsim_counter(0),
      DI(7) => GLOBAL_LOGIC0_68,
      DI(6) => GLOBAL_LOGIC0_68,
      DI(5) => GLOBAL_LOGIC0_69,
      DI(4) => GLOBAL_LOGIC0_69,
      DI(3) => GLOBAL_LOGIC0_68,
      DI(2) => GLOBAL_LOGIC0_70,
      DI(1) => GLOBAL_LOGIC0_68,
      DI(0) => GLOBAL_LOGIC0_69,
      DO(7) => txsim_ramout(7),
      DO(6) => txsim_ramout(6),
      DO(5) => txsim_ramout(5),
      DO(4) => txsim_ramout(4),
      DO(3) => txsim_ramout(3),
      DO(2) => txsim_ramout(2),
      DO(1) => txsim_ramout(1),
      DO(0) => txsim_ramout(0)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_0111 : X_MUX2
    port map (
      IA => memcontroller_N46780,
      IB => memcontroller_N46782,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_0_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_0111_G : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr4(0),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => addr2(0),
      O => memcontroller_N46782
    );
  memcontroller_Mmux_addrn_inst_mux_f5_0111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr1(0),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N46780
    );
  memcontroller_addrn_0_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_0_F5MUX,
      O => memcontroller_addrn(0)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_2111 : X_MUX2
    port map (
      IA => memcontroller_N46790,
      IB => memcontroller_N46792,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_2_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_2111_G : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => addr2(2),
      ADR3 => addr4(2),
      O => memcontroller_N46792
    );
  memcontroller_Mmux_addrn_inst_mux_f5_2111_F : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => addr1(2),
      O => memcontroller_N46790
    );
  memcontroller_addrn_2_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_2_F5MUX,
      O => memcontroller_addrn(2)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_3111 : X_MUX2
    port map (
      IA => memcontroller_N46795,
      IB => memcontroller_N46797,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_3_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_3111_G : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => addr2(3),
      ADR1 => VCC,
      ADR2 => addr4(3),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N46797
    );
  memcontroller_Mmux_addrn_inst_mux_f5_3111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr1(3),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N46795
    );
  memcontroller_addrn_3_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_3_F5MUX,
      O => memcontroller_addrn(3)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_4111 : X_MUX2
    port map (
      IA => memcontroller_N46800,
      IB => memcontroller_N46802,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_4_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_4111_G : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => addr2(4),
      ADR1 => addr4(4),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N46802
    );
  memcontroller_Mmux_addrn_inst_mux_f5_4111_F : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => addr1(4),
      O => memcontroller_N46800
    );
  memcontroller_addrn_4_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_4_F5MUX,
      O => memcontroller_addrn(4)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_1711 : X_MUX2
    port map (
      IA => memcontroller_N46785,
      IB => memcontroller_N46787,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_1_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_1711_G : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2(1),
      ADR2 => addr4(1),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N46787
    );
  memcontroller_Mmux_addrn_inst_mux_f5_1711_F : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => VCC,
      ADR3 => addr1(1),
      O => memcontroller_N46785
    );
  memcontroller_addrn_1_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_1_F5MUX,
      O => memcontroller_addrn(1)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_5111 : X_MUX2
    port map (
      IA => memcontroller_N46805,
      IB => memcontroller_N46807,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_5_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_5111_G : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => addr2(5),
      ADR1 => addr4(5),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N46807
    );
  memcontroller_Mmux_addrn_inst_mux_f5_5111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr1(5),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N46805
    );
  memcontroller_addrn_5_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_5_F5MUX,
      O => memcontroller_addrn(5)
    );
  memcontroller_addr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_0_OD,
      CE => MA_0_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_0_OFF_RST,
      O => memcontroller_ADDREXT(0)
    );
  MA_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_0_OFF_RST
    );
  memcontroller_Mmux_addrn_inst_mux_f5_6111 : X_MUX2
    port map (
      IA => memcontroller_N46810,
      IB => memcontroller_N46812,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_6_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_6111_G : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr4(6),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => addr2(6),
      O => memcontroller_N46812
    );
  memcontroller_Mmux_addrn_inst_mux_f5_6111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => addr1(6),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N46810
    );
  memcontroller_addrn_6_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_6_F5MUX,
      O => memcontroller_addrn(6)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_7111 : X_MUX2
    port map (
      IA => memcontroller_N46815,
      IB => memcontroller_N46817,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_7_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_7111_G : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => addr2(7),
      ADR3 => addr4(7),
      O => memcontroller_N46817
    );
  memcontroller_Mmux_addrn_inst_mux_f5_7111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => addr1(7),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N46815
    );
  memcontroller_addrn_7_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_7_F5MUX,
      O => memcontroller_addrn(7)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_8111 : X_MUX2
    port map (
      IA => memcontroller_N46820,
      IB => memcontroller_N46822,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_8_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_8111_G : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => addr2(8),
      ADR3 => addr4(8),
      O => memcontroller_N46822
    );
  memcontroller_Mmux_addrn_inst_mux_f5_8111_F : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => addr1(8),
      ADR3 => VCC,
      O => memcontroller_N46820
    );
  memcontroller_addrn_8_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_8_F5MUX,
      O => memcontroller_addrn(8)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_9111 : X_MUX2
    port map (
      IA => memcontroller_N46825,
      IB => memcontroller_N46827,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_9_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_9111_G : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => addr4(9),
      ADR3 => addr2(9),
      O => memcontroller_N46827
    );
  memcontroller_Mmux_addrn_inst_mux_f5_9111_F : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => addr1(9),
      ADR3 => VCC,
      O => memcontroller_N46825
    );
  memcontroller_addrn_9_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_9_F5MUX,
      O => memcontroller_addrn(9)
    );
  maccontrol_PHY_status_MII_Interface_sout414 : X_MUX2
    port map (
      IA => maccontrol_PHY_status_MII_Interface_N46760,
      IB => maccontrol_PHY_status_MII_Interface_N46762,
      SEL => maccontrol_PHY_status_MII_Interface_statecnt(2),
      O => maccontrol_PHY_status_MII_Interface_CHOICE826_F5MUX
    );
  maccontrol_PHY_status_MII_Interface_sout414_G : X_LUT4
    generic map(
      INIT => X"00A0"
    )
    port map (
      ADR0 => maccontrol_PHY_status_din(9),
      ADR1 => VCC,
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      O => maccontrol_PHY_status_MII_Interface_N46762
    );
  maccontrol_PHY_status_MII_Interface_sout414_F : X_LUT4
    generic map(
      INIT => X"008B"
    )
    port map (
      ADR0 => maccontrol_PHY_status_din(13),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR2 => maccontrol_PHY_status_miirw,
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      O => maccontrol_PHY_status_MII_Interface_N46760
    );
  maccontrol_PHY_status_MII_Interface_CHOICE826_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE826_F5MUX,
      O => maccontrol_PHY_status_MII_Interface_CHOICE826
    );
  memcontroller_Mmux_addrn_inst_mux_f5_10111 : X_MUX2
    port map (
      IA => memcontroller_N46830,
      IB => memcontroller_N46832,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_10_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_10111_G : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => addr4(10),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => addr2(10),
      O => memcontroller_N46832
    );
  memcontroller_Mmux_addrn_inst_mux_f5_10111_F : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => VCC,
      ADR3 => addr1(10),
      O => memcontroller_N46830
    );
  memcontroller_addrn_10_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_10_F5MUX,
      O => memcontroller_addrn(10)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_11111 : X_MUX2
    port map (
      IA => memcontroller_N46835,
      IB => memcontroller_N46837,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_11_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_11111_G : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => addr2(11),
      ADR1 => VCC,
      ADR2 => addr4(11),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N46837
    );
  memcontroller_Mmux_addrn_inst_mux_f5_11111_F : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr1(11),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N46835
    );
  memcontroller_addrn_11_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_11_F5MUX,
      O => memcontroller_addrn(11)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_12111 : X_MUX2
    port map (
      IA => memcontroller_N46840,
      IB => memcontroller_N46842,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_12_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_12111_G : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr4(12),
      ADR2 => addr2(12),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N46842
    );
  memcontroller_Mmux_addrn_inst_mux_f5_12111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr1(12),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N46840
    );
  memcontroller_addrn_12_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_12_F5MUX,
      O => memcontroller_addrn(12)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_13111 : X_MUX2
    port map (
      IA => memcontroller_N46845,
      IB => memcontroller_N46847,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_13_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_13111_G : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr4(13),
      ADR2 => addr2(13),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N46847
    );
  memcontroller_Mmux_addrn_inst_mux_f5_13111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr1(13),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N46845
    );
  memcontroller_addrn_13_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_13_F5MUX,
      O => memcontroller_addrn(13)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_14111 : X_MUX2
    port map (
      IA => memcontroller_N46765,
      IB => memcontroller_N46767,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_14_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_14111_G : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => addr2(14),
      ADR2 => VCC,
      ADR3 => addr4(14),
      O => memcontroller_N46767
    );
  memcontroller_Mmux_addrn_inst_mux_f5_14111_F : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => VCC,
      ADR3 => addr1(14),
      O => memcontroller_N46765
    );
  memcontroller_addrn_14_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_14_F5MUX,
      O => memcontroller_addrn(14)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_15111 : X_MUX2
    port map (
      IA => memcontroller_N46770,
      IB => memcontroller_N46772,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_15_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_15111_G : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => addr4(15),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => addr2(15),
      O => memcontroller_N46772
    );
  memcontroller_Mmux_addrn_inst_mux_f5_15111_F : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => addr1(15),
      O => memcontroller_N46770
    );
  memcontroller_addrn_15_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_15_F5MUX,
      O => memcontroller_addrn(15)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_16111 : X_MUX2
    port map (
      IA => memcontroller_N46775,
      IB => memcontroller_clknum_1_2_rt,
      SEL => memcontroller_clknum_0_2,
      O => memcontroller_addrn_16_F5MUX
    );
  memcontroller_clknum_1_2_rt_166 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_clknum_1_2_rt
    );
  memcontroller_Mmux_addrn_inst_mux_f5_16111_F : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N46775
    );
  memcontroller_addrn_16_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_16_F5MUX,
      O => memcontroller_addrn(16)
    );
  maccontrol_ledtx_cnt_123_LOGIC_ZERO_167 : X_ZERO
    port map (
      O => maccontrol_ledtx_cnt_123_LOGIC_ZERO
    );
  maccontrol_ledtx_cnt_123_LOGIC_ONE_168 : X_ONE
    port map (
      O => maccontrol_ledtx_cnt_123_LOGIC_ONE
    );
  maccontrol_ledtx_cnt_inst_cy_224_169 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_123_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_123_LOGIC_ZERO,
      SEL => maccontrol_ledtx_cnt_inst_lut3_155,
      O => maccontrol_ledtx_cnt_inst_cy_224
    );
  maccontrol_ledtx_cnt_inst_lut3_15511 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_ledtx_cnt_123,
      O => maccontrol_ledtx_cnt_inst_lut3_155
    );
  maccontrol_ledtx_cnt_inst_lut3_15611 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => maccontrol_ledtx_cnt_124,
      ADR3 => VCC,
      O => maccontrol_ledtx_cnt_inst_lut3_156
    );
  maccontrol_ledtx_cnt_123_COUTUSED : X_BUF
    port map (
      I => maccontrol_ledtx_cnt_123_CYMUXG,
      O => maccontrol_ledtx_cnt_inst_cy_225
    );
  maccontrol_ledtx_cnt_inst_cy_225_170 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_123_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_inst_cy_224,
      SEL => maccontrol_ledtx_cnt_inst_lut3_156,
      O => maccontrol_ledtx_cnt_123_CYMUXG
    );
  maccontrol_ledtx_cnt_inst_sum_178_171 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_inst_cy_224,
      I1 => maccontrol_ledtx_cnt_inst_lut3_156,
      O => maccontrol_ledtx_cnt_inst_sum_178
    );
  maccontrol_ledtx_cnt_125_LOGIC_ONE_172 : X_ONE
    port map (
      O => maccontrol_ledtx_cnt_125_LOGIC_ONE
    );
  maccontrol_ledtx_cnt_inst_cy_226_173 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_125_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_125_CYINIT,
      SEL => maccontrol_ledtx_cnt_inst_lut3_157,
      O => maccontrol_ledtx_cnt_inst_cy_226
    );
  maccontrol_ledtx_cnt_inst_sum_179_174 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_125_CYINIT,
      I1 => maccontrol_ledtx_cnt_inst_lut3_157,
      O => maccontrol_ledtx_cnt_inst_sum_179
    );
  maccontrol_ledtx_cnt_inst_lut3_15711 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_ledtx_cnt_125,
      O => maccontrol_ledtx_cnt_inst_lut3_157
    );
  maccontrol_ledtx_cnt_inst_lut3_15811 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_ledtx_cnt_126,
      O => maccontrol_ledtx_cnt_inst_lut3_158
    );
  maccontrol_ledtx_cnt_125_COUTUSED : X_BUF
    port map (
      I => maccontrol_ledtx_cnt_125_CYMUXG,
      O => maccontrol_ledtx_cnt_inst_cy_227
    );
  maccontrol_ledtx_cnt_inst_cy_227_175 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_125_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_inst_cy_226,
      SEL => maccontrol_ledtx_cnt_inst_lut3_158,
      O => maccontrol_ledtx_cnt_125_CYMUXG
    );
  maccontrol_ledtx_cnt_inst_sum_180_176 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_inst_cy_226,
      I1 => maccontrol_ledtx_cnt_inst_lut3_158,
      O => maccontrol_ledtx_cnt_inst_sum_180
    );
  maccontrol_ledtx_cnt_125_CYINIT_177 : X_BUF
    port map (
      I => maccontrol_ledtx_cnt_inst_cy_225,
      O => maccontrol_ledtx_cnt_125_CYINIT
    );
  maccontrol_ledtx_cnt_127_LOGIC_ONE_178 : X_ONE
    port map (
      O => maccontrol_ledtx_cnt_127_LOGIC_ONE
    );
  maccontrol_ledtx_cnt_inst_cy_228_179 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_127_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_127_CYINIT,
      SEL => maccontrol_ledtx_cnt_inst_lut3_159,
      O => maccontrol_ledtx_cnt_inst_cy_228
    );
  maccontrol_ledtx_cnt_inst_sum_181_180 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_127_CYINIT,
      I1 => maccontrol_ledtx_cnt_inst_lut3_159,
      O => maccontrol_ledtx_cnt_inst_sum_181
    );
  maccontrol_ledtx_cnt_inst_lut3_15911 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_ledtx_cnt_127,
      O => maccontrol_ledtx_cnt_inst_lut3_159
    );
  maccontrol_ledtx_cnt_inst_lut3_16011 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => maccontrol_ledtx_cnt_128,
      ADR3 => VCC,
      O => maccontrol_ledtx_cnt_inst_lut3_160
    );
  maccontrol_ledtx_cnt_127_COUTUSED : X_BUF
    port map (
      I => maccontrol_ledtx_cnt_127_CYMUXG,
      O => maccontrol_ledtx_cnt_inst_cy_229
    );
  maccontrol_ledtx_cnt_inst_cy_229_181 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_127_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_inst_cy_228,
      SEL => maccontrol_ledtx_cnt_inst_lut3_160,
      O => maccontrol_ledtx_cnt_127_CYMUXG
    );
  maccontrol_ledtx_cnt_inst_sum_182_182 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_inst_cy_228,
      I1 => maccontrol_ledtx_cnt_inst_lut3_160,
      O => maccontrol_ledtx_cnt_inst_sum_182
    );
  maccontrol_ledtx_cnt_127_CYINIT_183 : X_BUF
    port map (
      I => maccontrol_ledtx_cnt_inst_cy_227,
      O => maccontrol_ledtx_cnt_127_CYINIT
    );
  maccontrol_ledtx_cnt_129_LOGIC_ONE_184 : X_ONE
    port map (
      O => maccontrol_ledtx_cnt_129_LOGIC_ONE
    );
  maccontrol_ledtx_cnt_inst_cy_230_185 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_129_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_129_CYINIT,
      SEL => maccontrol_ledtx_cnt_inst_lut3_161,
      O => maccontrol_ledtx_cnt_inst_cy_230
    );
  maccontrol_ledtx_cnt_inst_sum_183_186 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_129_CYINIT,
      I1 => maccontrol_ledtx_cnt_inst_lut3_161,
      O => maccontrol_ledtx_cnt_inst_sum_183
    );
  maccontrol_ledtx_cnt_inst_lut3_16111 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_ledtx_cnt_129,
      O => maccontrol_ledtx_cnt_inst_lut3_161
    );
  maccontrol_ledtx_cnt_inst_lut3_16211 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_ledtx_cnt_130,
      O => maccontrol_ledtx_cnt_inst_lut3_162
    );
  maccontrol_ledtx_cnt_129_COUTUSED : X_BUF
    port map (
      I => maccontrol_ledtx_cnt_129_CYMUXG,
      O => maccontrol_ledtx_cnt_inst_cy_231
    );
  maccontrol_ledtx_cnt_inst_cy_231_187 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_129_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_inst_cy_230,
      SEL => maccontrol_ledtx_cnt_inst_lut3_162,
      O => maccontrol_ledtx_cnt_129_CYMUXG
    );
  maccontrol_ledtx_cnt_inst_sum_184_188 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_inst_cy_230,
      I1 => maccontrol_ledtx_cnt_inst_lut3_162,
      O => maccontrol_ledtx_cnt_inst_sum_184
    );
  maccontrol_ledtx_cnt_129_CYINIT_189 : X_BUF
    port map (
      I => maccontrol_ledtx_cnt_inst_cy_229,
      O => maccontrol_ledtx_cnt_129_CYINIT
    );
  maccontrol_ledtx_cnt_131_LOGIC_ONE_190 : X_ONE
    port map (
      O => maccontrol_ledtx_cnt_131_LOGIC_ONE
    );
  maccontrol_ledtx_cnt_inst_cy_232_191 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_131_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_131_CYINIT,
      SEL => maccontrol_ledtx_cnt_inst_lut3_163,
      O => maccontrol_ledtx_cnt_inst_cy_232
    );
  maccontrol_ledtx_cnt_inst_sum_185_192 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_131_CYINIT,
      I1 => maccontrol_ledtx_cnt_inst_lut3_163,
      O => maccontrol_ledtx_cnt_inst_sum_185
    );
  maccontrol_ledtx_cnt_inst_lut3_16311 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_ledtx_cnt_131,
      O => maccontrol_ledtx_cnt_inst_lut3_163
    );
  maccontrol_ledtx_cnt_inst_lut3_16411 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_ledtx_cnt_132,
      O => maccontrol_ledtx_cnt_inst_lut3_164
    );
  maccontrol_ledtx_cnt_131_COUTUSED : X_BUF
    port map (
      I => maccontrol_ledtx_cnt_131_CYMUXG,
      O => maccontrol_ledtx_cnt_inst_cy_233
    );
  maccontrol_ledtx_cnt_inst_cy_233_193 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_131_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_inst_cy_232,
      SEL => maccontrol_ledtx_cnt_inst_lut3_164,
      O => maccontrol_ledtx_cnt_131_CYMUXG
    );
  maccontrol_ledtx_cnt_inst_sum_186_194 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_inst_cy_232,
      I1 => maccontrol_ledtx_cnt_inst_lut3_164,
      O => maccontrol_ledtx_cnt_inst_sum_186
    );
  maccontrol_ledtx_cnt_131_CYINIT_195 : X_BUF
    port map (
      I => maccontrol_ledtx_cnt_inst_cy_231,
      O => maccontrol_ledtx_cnt_131_CYINIT
    );
  maccontrol_ledtx_cnt_133_LOGIC_ONE_196 : X_ONE
    port map (
      O => maccontrol_ledtx_cnt_133_LOGIC_ONE
    );
  maccontrol_ledtx_cnt_inst_cy_234_197 : X_MUX2
    port map (
      IA => maccontrol_ledtx_cnt_133_LOGIC_ONE,
      IB => maccontrol_ledtx_cnt_133_CYINIT,
      SEL => maccontrol_ledtx_cnt_inst_lut3_165,
      O => maccontrol_ledtx_cnt_inst_cy_234
    );
  maccontrol_ledtx_cnt_inst_sum_187_198 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_133_CYINIT,
      I1 => maccontrol_ledtx_cnt_inst_lut3_165,
      O => maccontrol_ledtx_cnt_inst_sum_187
    );
  maccontrol_ledtx_cnt_inst_lut3_16511 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_ledtx_cnt_133,
      O => maccontrol_ledtx_cnt_inst_lut3_165
    );
  maccontrol_ledtx_cnt_inst_lut3_16611 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_ledtx_cnt_134,
      O => maccontrol_ledtx_cnt_inst_lut3_166
    );
  maccontrol_ledtx_cnt_inst_sum_188_199 : X_XOR2
    port map (
      I0 => maccontrol_ledtx_cnt_inst_cy_234,
      I1 => maccontrol_ledtx_cnt_inst_lut3_166,
      O => maccontrol_ledtx_cnt_inst_sum_188
    );
  maccontrol_ledtx_cnt_133_CYINIT_200 : X_BUF
    port map (
      I => maccontrol_ledtx_cnt_inst_cy_233,
      O => maccontrol_ledtx_cnt_133_CYINIT
    );
  maccontrol_bitcnt_85_LOGIC_ZERO_201 : X_ZERO
    port map (
      O => maccontrol_bitcnt_85_LOGIC_ZERO
    );
  maccontrol_bitcnt_inst_cy_183_202 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_6,
      IB => maccontrol_bitcnt_85_LOGIC_ZERO,
      SEL => maccontrol_Mshreg_scslll_84_rt,
      O => maccontrol_bitcnt_inst_cy_183
    );
  maccontrol_Mshreg_scslll_84_rt_203 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_6,
      ADR1 => maccontrol_Mshreg_scslll_84,
      ADR2 => VCC,
      ADR3 => VCC,
      O => maccontrol_Mshreg_scslll_84_rt
    );
  maccontrol_bitcnt_inst_lut3_1171 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_57,
      ADR1 => maccontrol_Mshreg_scslll_84,
      ADR2 => VCC,
      ADR3 => maccontrol_bitcnt_85,
      O => maccontrol_bitcnt_inst_lut3_117
    );
  maccontrol_bitcnt_85_COUTUSED : X_BUF
    port map (
      I => maccontrol_bitcnt_85_CYMUXG,
      O => maccontrol_bitcnt_inst_cy_184
    );
  maccontrol_bitcnt_inst_cy_184_204 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_57,
      IB => maccontrol_bitcnt_inst_cy_183,
      SEL => maccontrol_bitcnt_inst_lut3_117,
      O => maccontrol_bitcnt_85_CYMUXG
    );
  maccontrol_bitcnt_inst_sum_139_205 : X_XOR2
    port map (
      I0 => maccontrol_bitcnt_inst_cy_183,
      I1 => maccontrol_bitcnt_inst_lut3_117,
      O => maccontrol_bitcnt_inst_sum_139
    );
  memcontroller_addr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_1_OD,
      CE => MA_1_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_1_OFF_RST,
      O => memcontroller_ADDREXT(1)
    );
  MA_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_1_OFF_RST
    );
  maccontrol_bitcnt_86_LOGIC_ZERO_206 : X_ZERO
    port map (
      O => maccontrol_bitcnt_86_LOGIC_ZERO
    );
  maccontrol_bitcnt_inst_cy_185_207 : X_MUX2
    port map (
      IA => maccontrol_bitcnt_86_LOGIC_ZERO,
      IB => maccontrol_bitcnt_86_CYINIT,
      SEL => maccontrol_bitcnt_inst_lut3_118,
      O => maccontrol_bitcnt_inst_cy_185
    );
  maccontrol_bitcnt_inst_sum_140_208 : X_XOR2
    port map (
      I0 => maccontrol_bitcnt_86_CYINIT,
      I1 => maccontrol_bitcnt_inst_lut3_118,
      O => maccontrol_bitcnt_inst_sum_140
    );
  maccontrol_bitcnt_inst_lut3_1181 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => maccontrol_Mshreg_scslll_84,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_bitcnt_86,
      O => maccontrol_bitcnt_inst_lut3_118
    );
  maccontrol_bitcnt_inst_lut3_1191 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => maccontrol_Mshreg_scslll_84,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_bitcnt_87,
      O => maccontrol_bitcnt_inst_lut3_119
    );
  maccontrol_bitcnt_86_COUTUSED : X_BUF
    port map (
      I => maccontrol_bitcnt_86_CYMUXG,
      O => maccontrol_bitcnt_inst_cy_186
    );
  maccontrol_bitcnt_inst_cy_186_209 : X_MUX2
    port map (
      IA => maccontrol_bitcnt_86_LOGIC_ZERO,
      IB => maccontrol_bitcnt_inst_cy_185,
      SEL => maccontrol_bitcnt_inst_lut3_119,
      O => maccontrol_bitcnt_86_CYMUXG
    );
  maccontrol_bitcnt_inst_sum_141_210 : X_XOR2
    port map (
      I0 => maccontrol_bitcnt_inst_cy_185,
      I1 => maccontrol_bitcnt_inst_lut3_119,
      O => maccontrol_bitcnt_inst_sum_141
    );
  maccontrol_bitcnt_86_CYINIT_211 : X_BUF
    port map (
      I => maccontrol_bitcnt_inst_cy_184,
      O => maccontrol_bitcnt_86_CYINIT
    );
  maccontrol_bitcnt_88_LOGIC_ZERO_212 : X_ZERO
    port map (
      O => maccontrol_bitcnt_88_LOGIC_ZERO
    );
  maccontrol_bitcnt_inst_cy_187_213 : X_MUX2
    port map (
      IA => maccontrol_bitcnt_88_LOGIC_ZERO,
      IB => maccontrol_bitcnt_88_CYINIT,
      SEL => maccontrol_bitcnt_inst_lut3_120,
      O => maccontrol_bitcnt_inst_cy_187
    );
  maccontrol_bitcnt_inst_sum_142_214 : X_XOR2
    port map (
      I0 => maccontrol_bitcnt_88_CYINIT,
      I1 => maccontrol_bitcnt_inst_lut3_120,
      O => maccontrol_bitcnt_inst_sum_142
    );
  maccontrol_bitcnt_inst_lut3_1201 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_bitcnt_88,
      ADR2 => maccontrol_Mshreg_scslll_84,
      ADR3 => VCC,
      O => maccontrol_bitcnt_inst_lut3_120
    );
  maccontrol_bitcnt_inst_lut3_1211 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => maccontrol_Mshreg_scslll_84,
      ADR1 => VCC,
      ADR2 => maccontrol_bitcnt_89,
      ADR3 => VCC,
      O => maccontrol_bitcnt_inst_lut3_121
    );
  maccontrol_bitcnt_88_COUTUSED : X_BUF
    port map (
      I => maccontrol_bitcnt_88_CYMUXG,
      O => maccontrol_bitcnt_inst_cy_188
    );
  maccontrol_bitcnt_inst_cy_188_215 : X_MUX2
    port map (
      IA => maccontrol_bitcnt_88_LOGIC_ZERO,
      IB => maccontrol_bitcnt_inst_cy_187,
      SEL => maccontrol_bitcnt_inst_lut3_121,
      O => maccontrol_bitcnt_88_CYMUXG
    );
  maccontrol_bitcnt_inst_sum_143_216 : X_XOR2
    port map (
      I0 => maccontrol_bitcnt_inst_cy_187,
      I1 => maccontrol_bitcnt_inst_lut3_121,
      O => maccontrol_bitcnt_inst_sum_143
    );
  maccontrol_bitcnt_88_CYINIT_217 : X_BUF
    port map (
      I => maccontrol_bitcnt_inst_cy_186,
      O => maccontrol_bitcnt_88_CYINIT
    );
  maccontrol_bitcnt_inst_sum_144_218 : X_XOR2
    port map (
      I0 => maccontrol_bitcnt_90_CYINIT,
      I1 => maccontrol_bitcnt_inst_lut3_122,
      O => maccontrol_bitcnt_inst_sum_144
    );
  maccontrol_bitcnt_inst_lut3_1221 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => maccontrol_Mshreg_scslll_84,
      ADR3 => maccontrol_bitcnt_90,
      O => maccontrol_bitcnt_inst_lut3_122
    );
  maccontrol_n00541_1_219 : X_LUT4
    generic map(
      INIT => X"0C00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_sclkdeltall,
      ADR2 => maccontrol_bitcnt_90,
      ADR3 => maccontrol_N30218,
      O => maccontrol_bitcnt_90_GROM
    );
  maccontrol_bitcnt_90_YUSED : X_BUF
    port map (
      I => maccontrol_bitcnt_90_GROM,
      O => maccontrol_n00541_1
    );
  maccontrol_bitcnt_90_CYINIT_220 : X_BUF
    port map (
      I => maccontrol_bitcnt_inst_cy_188,
      O => maccontrol_bitcnt_90_CYINIT
    );
  maccontrol_phyrstcnt_91_LOGIC_ONE_221 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_91_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_190_222 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_59,
      IB => maccontrol_phyrstcnt_91_LOGIC_ONE,
      SEL => maccontrol_N30228_rt,
      O => maccontrol_phyrstcnt_inst_cy_190
    );
  maccontrol_N30228_rt_223 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_59,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_N30228,
      O => maccontrol_N30228_rt
    );
  maccontrol_phyrstcnt_91_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_3,
      ADR1 => VCC,
      ADR2 => maccontrol_phyrstcnt_inst_lut3_1231_O,
      ADR3 => VCC,
      O => maccontrol_phyrstcnt_91_GROM
    );
  maccontrol_phyrstcnt_91_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_91_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_191
    );
  maccontrol_phyrstcnt_inst_cy_191_224 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_3,
      IB => maccontrol_phyrstcnt_inst_cy_190,
      SEL => maccontrol_phyrstcnt_91_GROM,
      O => maccontrol_phyrstcnt_91_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_145_225 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_190,
      I1 => maccontrol_phyrstcnt_91_GROM,
      O => maccontrol_phyrstcnt_inst_sum_145
    );
  maccontrol_phyrstcnt_92_LOGIC_ONE_226 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_92_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_192_227 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_92_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_92_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1241_O,
      O => maccontrol_phyrstcnt_inst_cy_192
    );
  maccontrol_phyrstcnt_inst_sum_146_228 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_92_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1241_O,
      O => maccontrol_phyrstcnt_inst_sum_146
    );
  maccontrol_phyrstcnt_inst_lut3_1241 : X_LUT4
    generic map(
      INIT => X"80FF"
    )
    port map (
      ADR0 => maccontrol_Ker303141_1,
      ADR1 => maccontrol_N46337,
      ADR2 => maccontrol_N30199,
      ADR3 => maccontrol_phyrstcnt_92,
      O => maccontrol_phyrstcnt_inst_lut3_1241_O
    );
  maccontrol_phyrstcnt_inst_lut3_1251 : X_LUT4
    generic map(
      INIT => X"B333"
    )
    port map (
      ADR0 => maccontrol_Ker303141_1,
      ADR1 => maccontrol_phyrstcnt_93,
      ADR2 => maccontrol_N30199,
      ADR3 => maccontrol_N46337,
      O => maccontrol_phyrstcnt_inst_lut3_1251_O
    );
  maccontrol_phyrstcnt_92_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_92_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_193
    );
  maccontrol_phyrstcnt_inst_cy_193_229 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_92_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_192,
      SEL => maccontrol_phyrstcnt_inst_lut3_1251_O,
      O => maccontrol_phyrstcnt_92_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_147_230 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_192,
      I1 => maccontrol_phyrstcnt_inst_lut3_1251_O,
      O => maccontrol_phyrstcnt_inst_sum_147
    );
  maccontrol_phyrstcnt_92_CYINIT_231 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_191,
      O => maccontrol_phyrstcnt_92_CYINIT
    );
  maccontrol_phyrstcnt_94_LOGIC_ONE_232 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_94_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_194_233 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_94_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_94_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1261_O,
      O => maccontrol_phyrstcnt_inst_cy_194
    );
  maccontrol_phyrstcnt_inst_sum_148_234 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_94_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1261_O,
      O => maccontrol_phyrstcnt_inst_sum_148
    );
  maccontrol_phyrstcnt_inst_lut3_1261 : X_LUT4
    generic map(
      INIT => X"B333"
    )
    port map (
      ADR0 => maccontrol_Ker303141_1,
      ADR1 => maccontrol_phyrstcnt_94,
      ADR2 => maccontrol_N30199,
      ADR3 => maccontrol_N46337,
      O => maccontrol_phyrstcnt_inst_lut3_1261_O
    );
  maccontrol_phyrstcnt_inst_lut3_1271 : X_LUT4
    generic map(
      INIT => X"1333"
    )
    port map (
      ADR0 => maccontrol_N46337,
      ADR1 => maccontrol_phyrstcnt_95,
      ADR2 => maccontrol_N30199,
      ADR3 => maccontrol_Ker303141_1,
      O => maccontrol_phyrstcnt_inst_lut3_1271_O
    );
  maccontrol_phyrstcnt_94_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_94_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_195
    );
  maccontrol_phyrstcnt_inst_cy_195_235 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_94_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_194,
      SEL => maccontrol_phyrstcnt_inst_lut3_1271_O,
      O => maccontrol_phyrstcnt_94_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_149_236 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_194,
      I1 => maccontrol_phyrstcnt_inst_lut3_1271_O,
      O => maccontrol_phyrstcnt_inst_sum_149
    );
  maccontrol_phyrstcnt_94_CYINIT_237 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_193,
      O => maccontrol_phyrstcnt_94_CYINIT
    );
  maccontrol_phyrstcnt_96_LOGIC_ONE_238 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_96_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_196_239 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_96_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_96_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1281_O,
      O => maccontrol_phyrstcnt_inst_cy_196
    );
  maccontrol_phyrstcnt_inst_sum_150_240 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_96_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1281_O,
      O => maccontrol_phyrstcnt_inst_sum_150
    );
  maccontrol_phyrstcnt_inst_lut3_1281 : X_LUT4
    generic map(
      INIT => X"B333"
    )
    port map (
      ADR0 => maccontrol_N46337,
      ADR1 => maccontrol_phyrstcnt_96,
      ADR2 => maccontrol_Ker303141_1,
      ADR3 => maccontrol_N30199,
      O => maccontrol_phyrstcnt_inst_lut3_1281_O
    );
  maccontrol_phyrstcnt_inst_lut3_1291 : X_LUT4
    generic map(
      INIT => X"1333"
    )
    port map (
      ADR0 => maccontrol_N46337,
      ADR1 => maccontrol_phyrstcnt_97,
      ADR2 => maccontrol_Ker303141_1,
      ADR3 => maccontrol_N30199,
      O => maccontrol_phyrstcnt_inst_lut3_1291_O
    );
  maccontrol_phyrstcnt_96_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_96_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_197
    );
  maccontrol_phyrstcnt_inst_cy_197_241 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_96_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_196,
      SEL => maccontrol_phyrstcnt_inst_lut3_1291_O,
      O => maccontrol_phyrstcnt_96_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_151_242 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_196,
      I1 => maccontrol_phyrstcnt_inst_lut3_1291_O,
      O => maccontrol_phyrstcnt_inst_sum_151
    );
  maccontrol_phyrstcnt_96_CYINIT_243 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_195,
      O => maccontrol_phyrstcnt_96_CYINIT
    );
  maccontrol_phyrstcnt_98_LOGIC_ONE_244 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_98_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_198_245 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_98_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_98_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1301_O,
      O => maccontrol_phyrstcnt_inst_cy_198
    );
  maccontrol_phyrstcnt_inst_sum_152_246 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_98_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1301_O,
      O => maccontrol_phyrstcnt_inst_sum_152
    );
  maccontrol_phyrstcnt_inst_lut3_1301 : X_LUT4
    generic map(
      INIT => X"007F"
    )
    port map (
      ADR0 => maccontrol_N46337,
      ADR1 => maccontrol_N30199,
      ADR2 => maccontrol_Ker303141_1,
      ADR3 => maccontrol_phyrstcnt_98,
      O => maccontrol_phyrstcnt_inst_lut3_1301_O
    );
  maccontrol_phyrstcnt_inst_lut3_1311 : X_LUT4
    generic map(
      INIT => X"1555"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_99,
      ADR1 => maccontrol_N46337,
      ADR2 => maccontrol_Ker303141_1,
      ADR3 => maccontrol_N30199,
      O => maccontrol_phyrstcnt_inst_lut3_1311_O
    );
  maccontrol_phyrstcnt_98_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_98_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_199
    );
  maccontrol_phyrstcnt_inst_cy_199_247 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_98_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_198,
      SEL => maccontrol_phyrstcnt_inst_lut3_1311_O,
      O => maccontrol_phyrstcnt_98_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_153_248 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_198,
      I1 => maccontrol_phyrstcnt_inst_lut3_1311_O,
      O => maccontrol_phyrstcnt_inst_sum_153
    );
  maccontrol_phyrstcnt_98_CYINIT_249 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_197,
      O => maccontrol_phyrstcnt_98_CYINIT
    );
  maccontrol_phyrstcnt_100_LOGIC_ONE_250 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_100_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_200_251 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_100_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_100_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1321_O,
      O => maccontrol_phyrstcnt_inst_cy_200
    );
  maccontrol_phyrstcnt_inst_sum_154_252 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_100_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1321_O,
      O => maccontrol_phyrstcnt_inst_sum_154
    );
  maccontrol_phyrstcnt_inst_lut3_1321 : X_LUT4
    generic map(
      INIT => X"007F"
    )
    port map (
      ADR0 => maccontrol_N46337,
      ADR1 => maccontrol_N30199,
      ADR2 => maccontrol_Ker303141_1,
      ADR3 => maccontrol_phyrstcnt_100,
      O => maccontrol_phyrstcnt_inst_lut3_1321_O
    );
  maccontrol_phyrstcnt_inst_lut3_1331 : X_LUT4
    generic map(
      INIT => X"070F"
    )
    port map (
      ADR0 => maccontrol_N46337,
      ADR1 => maccontrol_N30199,
      ADR2 => maccontrol_phyrstcnt_101,
      ADR3 => maccontrol_Ker303141_1,
      O => maccontrol_phyrstcnt_inst_lut3_1331_O
    );
  maccontrol_phyrstcnt_100_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_100_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_201
    );
  maccontrol_phyrstcnt_inst_cy_201_253 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_100_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_200,
      SEL => maccontrol_phyrstcnt_inst_lut3_1331_O,
      O => maccontrol_phyrstcnt_100_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_155_254 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_200,
      I1 => maccontrol_phyrstcnt_inst_lut3_1331_O,
      O => maccontrol_phyrstcnt_inst_sum_155
    );
  maccontrol_phyrstcnt_100_CYINIT_255 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_199,
      O => maccontrol_phyrstcnt_100_CYINIT
    );
  maccontrol_phyrstcnt_102_LOGIC_ONE_256 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_102_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_202_257 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_102_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_102_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1341_O,
      O => maccontrol_phyrstcnt_inst_cy_202
    );
  maccontrol_phyrstcnt_inst_sum_156_258 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_102_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1341_O,
      O => maccontrol_phyrstcnt_inst_sum_156
    );
  maccontrol_phyrstcnt_inst_lut3_1341 : X_LUT4
    generic map(
      INIT => X"B333"
    )
    port map (
      ADR0 => maccontrol_N46337,
      ADR1 => maccontrol_phyrstcnt_102,
      ADR2 => maccontrol_N30199,
      ADR3 => maccontrol_Ker303141_2,
      O => maccontrol_phyrstcnt_inst_lut3_1341_O
    );
  maccontrol_phyrstcnt_inst_lut3_1351 : X_LUT4
    generic map(
      INIT => X"80FF"
    )
    port map (
      ADR0 => maccontrol_N46337,
      ADR1 => maccontrol_Ker303141_2,
      ADR2 => maccontrol_N30199,
      ADR3 => maccontrol_phyrstcnt_103,
      O => maccontrol_phyrstcnt_inst_lut3_1351_O
    );
  maccontrol_phyrstcnt_102_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_102_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_203
    );
  maccontrol_phyrstcnt_inst_cy_203_259 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_102_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_202,
      SEL => maccontrol_phyrstcnt_inst_lut3_1351_O,
      O => maccontrol_phyrstcnt_102_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_157_260 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_202,
      I1 => maccontrol_phyrstcnt_inst_lut3_1351_O,
      O => maccontrol_phyrstcnt_inst_sum_157
    );
  maccontrol_phyrstcnt_102_CYINIT_261 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_201,
      O => maccontrol_phyrstcnt_102_CYINIT
    );
  maccontrol_phyrstcnt_104_LOGIC_ONE_262 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_104_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_204_263 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_104_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_104_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1361_O,
      O => maccontrol_phyrstcnt_inst_cy_204
    );
  maccontrol_phyrstcnt_inst_sum_158_264 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_104_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1361_O,
      O => maccontrol_phyrstcnt_inst_sum_158
    );
  maccontrol_phyrstcnt_inst_lut3_1361 : X_LUT4
    generic map(
      INIT => X"D555"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_104,
      ADR1 => maccontrol_N30285,
      ADR2 => maccontrol_Ker303141_2,
      ADR3 => maccontrol_N46356,
      O => maccontrol_phyrstcnt_inst_lut3_1361_O
    );
  maccontrol_phyrstcnt_inst_lut3_1371 : X_LUT4
    generic map(
      INIT => X"D555"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_105,
      ADR1 => maccontrol_N30285,
      ADR2 => maccontrol_Ker303141_2,
      ADR3 => maccontrol_N46356,
      O => maccontrol_phyrstcnt_inst_lut3_1371_O
    );
  maccontrol_phyrstcnt_104_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_104_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_205
    );
  maccontrol_phyrstcnt_inst_cy_205_265 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_104_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_204,
      SEL => maccontrol_phyrstcnt_inst_lut3_1371_O,
      O => maccontrol_phyrstcnt_104_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_159_266 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_204,
      I1 => maccontrol_phyrstcnt_inst_lut3_1371_O,
      O => maccontrol_phyrstcnt_inst_sum_159
    );
  maccontrol_phyrstcnt_104_CYINIT_267 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_203,
      O => maccontrol_phyrstcnt_104_CYINIT
    );
  maccontrol_phyrstcnt_106_LOGIC_ONE_268 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_106_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_206_269 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_106_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_106_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1381_O,
      O => maccontrol_phyrstcnt_inst_cy_206
    );
  maccontrol_phyrstcnt_inst_sum_160_270 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_106_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1381_O,
      O => maccontrol_phyrstcnt_inst_sum_160
    );
  maccontrol_phyrstcnt_inst_lut3_1381 : X_LUT4
    generic map(
      INIT => X"80FF"
    )
    port map (
      ADR0 => maccontrol_Ker303141_2,
      ADR1 => maccontrol_N30285,
      ADR2 => maccontrol_N46356,
      ADR3 => maccontrol_phyrstcnt_106,
      O => maccontrol_phyrstcnt_inst_lut3_1381_O
    );
  maccontrol_phyrstcnt_inst_lut3_1391 : X_LUT4
    generic map(
      INIT => X"D555"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_107,
      ADR1 => maccontrol_N30285,
      ADR2 => maccontrol_Ker303141_2,
      ADR3 => maccontrol_N46356,
      O => maccontrol_phyrstcnt_inst_lut3_1391_O
    );
  maccontrol_phyrstcnt_106_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_106_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_207
    );
  maccontrol_phyrstcnt_inst_cy_207_271 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_106_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_206,
      SEL => maccontrol_phyrstcnt_inst_lut3_1391_O,
      O => maccontrol_phyrstcnt_106_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_161_272 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_206,
      I1 => maccontrol_phyrstcnt_inst_lut3_1391_O,
      O => maccontrol_phyrstcnt_inst_sum_161
    );
  maccontrol_phyrstcnt_106_CYINIT_273 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_205,
      O => maccontrol_phyrstcnt_106_CYINIT
    );
  maccontrol_phyrstcnt_108_LOGIC_ONE_274 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_108_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_208_275 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_108_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_108_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1401_O,
      O => maccontrol_phyrstcnt_inst_cy_208
    );
  maccontrol_phyrstcnt_inst_sum_162_276 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_108_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1401_O,
      O => maccontrol_phyrstcnt_inst_sum_162
    );
  maccontrol_phyrstcnt_inst_lut3_1401 : X_LUT4
    generic map(
      INIT => X"D555"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_108,
      ADR1 => maccontrol_N30285,
      ADR2 => maccontrol_N46356,
      ADR3 => maccontrol_Ker303141_2,
      O => maccontrol_phyrstcnt_inst_lut3_1401_O
    );
  maccontrol_phyrstcnt_inst_lut3_1411 : X_LUT4
    generic map(
      INIT => X"B333"
    )
    port map (
      ADR0 => maccontrol_N46356,
      ADR1 => maccontrol_phyrstcnt_109,
      ADR2 => maccontrol_N30285,
      ADR3 => maccontrol_Ker303141_2,
      O => maccontrol_phyrstcnt_inst_lut3_1411_O
    );
  maccontrol_phyrstcnt_108_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_108_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_209
    );
  maccontrol_phyrstcnt_inst_cy_209_277 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_108_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_208,
      SEL => maccontrol_phyrstcnt_inst_lut3_1411_O,
      O => maccontrol_phyrstcnt_108_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_163_278 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_208,
      I1 => maccontrol_phyrstcnt_inst_lut3_1411_O,
      O => maccontrol_phyrstcnt_inst_sum_163
    );
  maccontrol_phyrstcnt_108_CYINIT_279 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_207,
      O => maccontrol_phyrstcnt_108_CYINIT
    );
  maccontrol_phyrstcnt_110_LOGIC_ONE_280 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_110_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_210_281 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_110_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_110_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1421_O,
      O => maccontrol_phyrstcnt_inst_cy_210
    );
  maccontrol_phyrstcnt_inst_sum_164_282 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_110_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1421_O,
      O => maccontrol_phyrstcnt_inst_sum_164
    );
  maccontrol_phyrstcnt_inst_lut3_1421 : X_LUT4
    generic map(
      INIT => X"F3F3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_phyrstcnt_110,
      ADR2 => maccontrol_N30228,
      ADR3 => VCC,
      O => maccontrol_phyrstcnt_inst_lut3_1421_O
    );
  maccontrol_phyrstcnt_inst_lut3_1431 : X_LUT4
    generic map(
      INIT => X"FF0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => maccontrol_phyrstcnt_111,
      ADR3 => maccontrol_N30228,
      O => maccontrol_phyrstcnt_inst_lut3_1431_O
    );
  maccontrol_phyrstcnt_110_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_110_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_211
    );
  maccontrol_phyrstcnt_inst_cy_211_283 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_110_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_210,
      SEL => maccontrol_phyrstcnt_inst_lut3_1431_O,
      O => maccontrol_phyrstcnt_110_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_165_284 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_210,
      I1 => maccontrol_phyrstcnt_inst_lut3_1431_O,
      O => maccontrol_phyrstcnt_inst_sum_165
    );
  maccontrol_phyrstcnt_110_CYINIT_285 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_209,
      O => maccontrol_phyrstcnt_110_CYINIT
    );
  maccontrol_phyrstcnt_112_LOGIC_ONE_286 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_112_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_212_287 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_112_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_112_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1441_O,
      O => maccontrol_phyrstcnt_inst_cy_212
    );
  maccontrol_phyrstcnt_inst_sum_166_288 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_112_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1441_O,
      O => maccontrol_phyrstcnt_inst_sum_166
    );
  maccontrol_phyrstcnt_inst_lut3_1441 : X_LUT4
    generic map(
      INIT => X"DDDD"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_112,
      ADR1 => maccontrol_N30228,
      ADR2 => VCC,
      ADR3 => VCC,
      O => maccontrol_phyrstcnt_inst_lut3_1441_O
    );
  maccontrol_phyrstcnt_inst_lut3_1451 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => maccontrol_N30228,
      ADR1 => VCC,
      ADR2 => maccontrol_phyrstcnt_113,
      ADR3 => VCC,
      O => maccontrol_phyrstcnt_inst_lut3_1451_O
    );
  maccontrol_phyrstcnt_112_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_112_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_213
    );
  maccontrol_phyrstcnt_inst_cy_213_289 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_112_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_212,
      SEL => maccontrol_phyrstcnt_inst_lut3_1451_O,
      O => maccontrol_phyrstcnt_112_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_167_290 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_212,
      I1 => maccontrol_phyrstcnt_inst_lut3_1451_O,
      O => maccontrol_phyrstcnt_inst_sum_167
    );
  maccontrol_phyrstcnt_112_CYINIT_291 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_211,
      O => maccontrol_phyrstcnt_112_CYINIT
    );
  maccontrol_phyrstcnt_114_LOGIC_ONE_292 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_114_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_214_293 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_114_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_114_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1461_O,
      O => maccontrol_phyrstcnt_inst_cy_214
    );
  maccontrol_phyrstcnt_inst_sum_168_294 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_114_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1461_O,
      O => maccontrol_phyrstcnt_inst_sum_168
    );
  maccontrol_phyrstcnt_inst_lut3_1461 : X_LUT4
    generic map(
      INIT => X"CCFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_N30228,
      ADR2 => VCC,
      ADR3 => maccontrol_phyrstcnt_114,
      O => maccontrol_phyrstcnt_inst_lut3_1461_O
    );
  maccontrol_phyrstcnt_inst_lut3_1471 : X_LUT4
    generic map(
      INIT => X"AAFF"
    )
    port map (
      ADR0 => maccontrol_N30228,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_phyrstcnt_115,
      O => maccontrol_phyrstcnt_inst_lut3_1471_O
    );
  maccontrol_phyrstcnt_114_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_114_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_215
    );
  maccontrol_phyrstcnt_inst_cy_215_295 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_114_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_214,
      SEL => maccontrol_phyrstcnt_inst_lut3_1471_O,
      O => maccontrol_phyrstcnt_114_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_169_296 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_214,
      I1 => maccontrol_phyrstcnt_inst_lut3_1471_O,
      O => maccontrol_phyrstcnt_inst_sum_169
    );
  maccontrol_phyrstcnt_114_CYINIT_297 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_213,
      O => maccontrol_phyrstcnt_114_CYINIT
    );
  maccontrol_phyrstcnt_116_LOGIC_ONE_298 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_116_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_216_299 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_116_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_116_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1481_O,
      O => maccontrol_phyrstcnt_inst_cy_216
    );
  maccontrol_phyrstcnt_inst_sum_170_300 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_116_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1481_O,
      O => maccontrol_phyrstcnt_inst_sum_170
    );
  maccontrol_phyrstcnt_inst_lut3_1481 : X_LUT4
    generic map(
      INIT => X"CCFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_N30228,
      ADR2 => VCC,
      ADR3 => maccontrol_phyrstcnt_116,
      O => maccontrol_phyrstcnt_inst_lut3_1481_O
    );
  maccontrol_phyrstcnt_inst_lut3_1491 : X_LUT4
    generic map(
      INIT => X"CCFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_N30228,
      ADR2 => VCC,
      ADR3 => maccontrol_phyrstcnt_117,
      O => maccontrol_phyrstcnt_inst_lut3_1491_O
    );
  maccontrol_phyrstcnt_116_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_116_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_217
    );
  maccontrol_phyrstcnt_inst_cy_217_301 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_116_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_216,
      SEL => maccontrol_phyrstcnt_inst_lut3_1491_O,
      O => maccontrol_phyrstcnt_116_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_171_302 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_216,
      I1 => maccontrol_phyrstcnt_inst_lut3_1491_O,
      O => maccontrol_phyrstcnt_inst_sum_171
    );
  maccontrol_phyrstcnt_116_CYINIT_303 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_215,
      O => maccontrol_phyrstcnt_116_CYINIT
    );
  maccontrol_phyrstcnt_118_LOGIC_ONE_304 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_118_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_218_305 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_118_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_118_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1501_O,
      O => maccontrol_phyrstcnt_inst_cy_218
    );
  maccontrol_phyrstcnt_inst_sum_172_306 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_118_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1501_O,
      O => maccontrol_phyrstcnt_inst_sum_172
    );
  maccontrol_phyrstcnt_inst_lut3_1501 : X_LUT4
    generic map(
      INIT => X"FF33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_phyrstcnt_118,
      ADR2 => VCC,
      ADR3 => maccontrol_N30228,
      O => maccontrol_phyrstcnt_inst_lut3_1501_O
    );
  maccontrol_phyrstcnt_inst_lut3_1511 : X_LUT4
    generic map(
      INIT => X"FF0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => maccontrol_phyrstcnt_119,
      ADR3 => maccontrol_N30228,
      O => maccontrol_phyrstcnt_inst_lut3_1511_O
    );
  maccontrol_phyrstcnt_118_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_118_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_219
    );
  maccontrol_phyrstcnt_inst_cy_219_307 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_118_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_218,
      SEL => maccontrol_phyrstcnt_inst_lut3_1511_O,
      O => maccontrol_phyrstcnt_118_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_173_308 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_218,
      I1 => maccontrol_phyrstcnt_inst_lut3_1511_O,
      O => maccontrol_phyrstcnt_inst_sum_173
    );
  maccontrol_phyrstcnt_118_CYINIT_309 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_217,
      O => maccontrol_phyrstcnt_118_CYINIT
    );
  maccontrol_phyrstcnt_120_LOGIC_ONE_310 : X_ONE
    port map (
      O => maccontrol_phyrstcnt_120_LOGIC_ONE
    );
  maccontrol_phyrstcnt_inst_cy_220_311 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_120_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_120_CYINIT,
      SEL => maccontrol_phyrstcnt_inst_lut3_1521_O,
      O => maccontrol_phyrstcnt_inst_cy_220
    );
  maccontrol_phyrstcnt_inst_sum_174_312 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_120_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1521_O,
      O => maccontrol_phyrstcnt_inst_sum_174
    );
  maccontrol_phyrstcnt_inst_lut3_1521 : X_LUT4
    generic map(
      INIT => X"BBBB"
    )
    port map (
      ADR0 => maccontrol_N30228,
      ADR1 => maccontrol_phyrstcnt_120,
      ADR2 => VCC,
      ADR3 => VCC,
      O => maccontrol_phyrstcnt_inst_lut3_1521_O
    );
  maccontrol_phyrstcnt_inst_lut3_1531 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => maccontrol_N30228,
      ADR1 => VCC,
      ADR2 => maccontrol_phyrstcnt_121,
      ADR3 => VCC,
      O => maccontrol_phyrstcnt_inst_lut3_1531_O
    );
  maccontrol_phyrstcnt_120_COUTUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_120_CYMUXG,
      O => maccontrol_phyrstcnt_inst_cy_221
    );
  maccontrol_phyrstcnt_inst_cy_221_313 : X_MUX2
    port map (
      IA => maccontrol_phyrstcnt_120_LOGIC_ONE,
      IB => maccontrol_phyrstcnt_inst_cy_220,
      SEL => maccontrol_phyrstcnt_inst_lut3_1531_O,
      O => maccontrol_phyrstcnt_120_CYMUXG
    );
  maccontrol_phyrstcnt_inst_sum_175_314 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_inst_cy_220,
      I1 => maccontrol_phyrstcnt_inst_lut3_1531_O,
      O => maccontrol_phyrstcnt_inst_sum_175
    );
  maccontrol_phyrstcnt_120_CYINIT_315 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_219,
      O => maccontrol_phyrstcnt_120_CYINIT
    );
  memcontroller_addr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_2_OD,
      CE => MA_2_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_2_OFF_RST,
      O => memcontroller_ADDREXT(2)
    );
  MA_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_2_OFF_RST
    );
  maccontrol_phyrstcnt_inst_sum_176_316 : X_XOR2
    port map (
      I0 => maccontrol_phyrstcnt_122_CYINIT,
      I1 => maccontrol_phyrstcnt_inst_lut3_1541_O,
      O => maccontrol_phyrstcnt_inst_sum_176
    );
  maccontrol_phyrstcnt_inst_lut3_1541 : X_LUT4
    generic map(
      INIT => X"BBBB"
    )
    port map (
      ADR0 => maccontrol_N30228,
      ADR1 => maccontrol_phyrstcnt_122,
      ADR2 => VCC,
      ADR3 => VCC,
      O => maccontrol_phyrstcnt_inst_lut3_1541_O
    );
  maccontrol_n0039124_1_317 : X_LUT4
    generic map(
      INIT => X"00A8"
    )
    port map (
      ADR0 => clkslen,
      ADR1 => maccontrol_N30228,
      ADR2 => maccontrol_CHOICE1608,
      ADR3 => RESET_IBUF,
      O => maccontrol_phyrstcnt_122_GROM
    );
  maccontrol_phyrstcnt_122_YUSED : X_BUF
    port map (
      I => maccontrol_phyrstcnt_122_GROM,
      O => maccontrol_n0039124_1
    );
  maccontrol_phyrstcnt_122_CYINIT_318 : X_BUF
    port map (
      I => maccontrol_phyrstcnt_inst_cy_221,
      O => maccontrol_phyrstcnt_122_CYINIT
    );
  cnt0_0_LOGIC_ZERO_319 : X_ZERO
    port map (
      O => cnt0_0_LOGIC_ZERO
    );
  cnt0_Madd_n0000_inst_cy_24_320 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_30,
      IB => cnt0_0_LOGIC_ZERO,
      SEL => cnt0_Madd_n0000_inst_lut2_24,
      O => cnt0_Madd_n0000_inst_cy_24
    );
  cnt0_Madd_n0000_inst_lut2_241 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_30,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => cnt0(0),
      O => cnt0_Madd_n0000_inst_lut2_24
    );
  cnt0_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_38,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => cnt0(1),
      O => cnt0_0_GROM
    );
  cnt0_0_COUTUSED : X_BUF
    port map (
      I => cnt0_0_CYMUXG,
      O => cnt0_Madd_n0000_inst_cy_25
    );
  cnt0_Madd_n0000_inst_cy_25_321 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_38,
      IB => cnt0_Madd_n0000_inst_cy_24,
      SEL => cnt0_0_GROM,
      O => cnt0_0_CYMUXG
    );
  cnt0_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => cnt0_Madd_n0000_inst_cy_24,
      I1 => cnt0_0_GROM,
      O => cnt0_n0000(1)
    );
  cnt0_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => cnt0_n0000(3),
      CE => Q_n0034,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => err,
      O => cnt0(3)
    );
  cnt0_2_LOGIC_ZERO_322 : X_ZERO
    port map (
      O => cnt0_2_LOGIC_ZERO
    );
  cnt0_Madd_n0000_inst_cy_26_323 : X_MUX2
    port map (
      IA => cnt0_2_LOGIC_ZERO,
      IB => cnt0_2_CYINIT,
      SEL => cnt0_2_FROM,
      O => cnt0_Madd_n0000_inst_cy_26
    );
  cnt0_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => cnt0_2_CYINIT,
      I1 => cnt0_2_FROM,
      O => cnt0_n0000(2)
    );
  cnt0_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => cnt0(2),
      O => cnt0_2_FROM
    );
  cnt0_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt0(3),
      ADR3 => VCC,
      O => cnt0_2_GROM
    );
  cnt0_2_COUTUSED : X_BUF
    port map (
      I => cnt0_2_CYMUXG,
      O => cnt0_Madd_n0000_inst_cy_27
    );
  cnt0_Madd_n0000_inst_cy_27_324 : X_MUX2
    port map (
      IA => cnt0_2_LOGIC_ZERO,
      IB => cnt0_Madd_n0000_inst_cy_26,
      SEL => cnt0_2_GROM,
      O => cnt0_2_CYMUXG
    );
  cnt0_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => cnt0_Madd_n0000_inst_cy_26,
      I1 => cnt0_2_GROM,
      O => cnt0_n0000(3)
    );
  cnt0_2_CYINIT_325 : X_BUF
    port map (
      I => cnt0_Madd_n0000_inst_cy_25,
      O => cnt0_2_CYINIT
    );
  cnt0_4_LOGIC_ZERO_326 : X_ZERO
    port map (
      O => cnt0_4_LOGIC_ZERO
    );
  cnt0_Madd_n0000_inst_cy_28_327 : X_MUX2
    port map (
      IA => cnt0_4_LOGIC_ZERO,
      IB => cnt0_4_CYINIT,
      SEL => cnt0_4_FROM,
      O => cnt0_Madd_n0000_inst_cy_28
    );
  cnt0_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => cnt0_4_CYINIT,
      I1 => cnt0_4_FROM,
      O => cnt0_n0000(4)
    );
  cnt0_4_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => cnt0(4),
      O => cnt0_4_FROM
    );
  cnt0_5_rt_328 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt0(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt0_5_rt
    );
  cnt0_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => cnt0_Madd_n0000_inst_cy_28,
      I1 => cnt0_5_rt,
      O => cnt0_n0000(5)
    );
  cnt0_4_CYINIT_329 : X_BUF
    port map (
      I => cnt0_Madd_n0000_inst_cy_27,
      O => cnt0_4_CYINIT
    );
  memtest2_Mcompar_n0020_inst_cy_167_LOGIC_ONE_330 : X_ONE
    port map (
      O => memtest2_Mcompar_n0020_inst_cy_167_LOGIC_ONE
    );
  memtest2_Mcompar_n0020_inst_cy_167_LOGIC_ZERO_331 : X_ZERO
    port map (
      O => memtest2_Mcompar_n0020_inst_cy_167_LOGIC_ZERO
    );
  memtest2_Mcompar_n0020_inst_cy_166_332 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0020_inst_cy_167_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0020_inst_cy_167_LOGIC_ONE,
      SEL => memtest2_Mcompar_n0020_inst_lut4_25,
      O => memtest2_Mcompar_n0020_inst_cy_166
    );
  memtest2_Mcompar_n0020_inst_lut4_251 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest2_Mshreg_data4_24_45,
      ADR1 => memtest2_datain(25),
      ADR2 => memtest2_Mshreg_data4_25_44,
      ADR3 => memtest2_datain(24),
      O => memtest2_Mcompar_n0020_inst_lut4_25
    );
  memtest2_Mcompar_n0020_inst_lut4_261 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest2_datain(26),
      ADR1 => memtest2_datain(27),
      ADR2 => memtest2_Mshreg_data4_27_42,
      ADR3 => memtest2_Mshreg_data4_26_43,
      O => memtest2_Mcompar_n0020_inst_lut4_26
    );
  memtest2_Mcompar_n0020_inst_cy_167_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0020_inst_cy_167_CYMUXG,
      O => memtest2_Mcompar_n0020_inst_cy_167
    );
  memtest2_Mcompar_n0020_inst_cy_167_333 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0020_inst_cy_167_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0020_inst_cy_166,
      SEL => memtest2_Mcompar_n0020_inst_lut4_26,
      O => memtest2_Mcompar_n0020_inst_cy_167_CYMUXG
    );
  memtest2_deq_3_LOGIC_ZERO_334 : X_ZERO
    port map (
      O => memtest2_deq_3_LOGIC_ZERO
    );
  memtest2_Mcompar_n0020_inst_cy_168_335 : X_MUX2
    port map (
      IA => memtest2_deq_3_LOGIC_ZERO,
      IB => memtest2_deq_3_CYINIT,
      SEL => memtest2_Mcompar_n0020_inst_lut4_27,
      O => memtest2_Mcompar_n0020_inst_cy_168
    );
  memtest2_Mcompar_n0020_inst_lut4_271 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest2_datain(28),
      ADR1 => memtest2_datain(29),
      ADR2 => memtest2_Mshreg_data4_29_40,
      ADR3 => memtest2_Mshreg_data4_28_41,
      O => memtest2_Mcompar_n0020_inst_lut4_27
    );
  memtest2_Mcompar_n0020_inst_lut4_281 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest2_Mshreg_data4_30_39,
      ADR1 => memtest2_datain(31),
      ADR2 => memtest2_Mshreg_data4_31_38,
      ADR3 => memtest2_datain(30),
      O => memtest2_Mcompar_n0020_inst_lut4_28
    );
  memtest2_deq_3_COUTUSED : X_BUF
    port map (
      I => memtest2_deq_3_CYMUXG,
      O => memtest2_deq(3)
    );
  memtest2_Mcompar_n0020_inst_cy_169 : X_MUX2
    port map (
      IA => memtest2_deq_3_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0020_inst_cy_168,
      SEL => memtest2_Mcompar_n0020_inst_lut4_28,
      O => memtest2_deq_3_CYMUXG
    );
  memtest2_deq_3_CYINIT_336 : X_BUF
    port map (
      I => memtest2_Mcompar_n0020_inst_cy_167,
      O => memtest2_deq_3_CYINIT
    );
  cnt_0_LOGIC_ZERO_337 : X_ZERO
    port map (
      O => cnt_0_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_0_338 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_8,
      IB => cnt_0_LOGIC_ZERO,
      SEL => Madd_n0000_inst_lut2_0,
      O => Madd_n0000_inst_cy_0
    );
  Madd_n0000_inst_lut2_01 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_8,
      ADR1 => cnt(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => Madd_n0000_inst_lut2_0
    );
  cnt_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_54,
      ADR1 => VCC,
      ADR2 => cnt(1),
      ADR3 => VCC,
      O => cnt_0_GROM
    );
  cnt_0_COUTUSED : X_BUF
    port map (
      I => cnt_0_CYMUXG,
      O => Madd_n0000_inst_cy_1
    );
  Madd_n0000_inst_cy_1_339 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_54,
      IB => Madd_n0000_inst_cy_0,
      SEL => cnt_0_GROM,
      O => cnt_0_CYMUXG
    );
  Madd_n0000_inst_sum_1 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_0,
      I1 => cnt_0_GROM,
      O => Q_n0000(1)
    );
  cnt_2_LOGIC_ZERO_340 : X_ZERO
    port map (
      O => cnt_2_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_2_341 : X_MUX2
    port map (
      IA => cnt_2_LOGIC_ZERO,
      IB => cnt_2_CYINIT,
      SEL => cnt_2_FROM,
      O => Madd_n0000_inst_cy_2
    );
  Madd_n0000_inst_sum_2 : X_XOR2
    port map (
      I0 => cnt_2_CYINIT,
      I1 => cnt_2_FROM,
      O => Q_n0000(2)
    );
  cnt_2_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_2_FROM
    );
  cnt_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(3),
      ADR3 => VCC,
      O => cnt_2_GROM
    );
  cnt_2_COUTUSED : X_BUF
    port map (
      I => cnt_2_CYMUXG,
      O => Madd_n0000_inst_cy_3
    );
  Madd_n0000_inst_cy_3_342 : X_MUX2
    port map (
      IA => cnt_2_LOGIC_ZERO,
      IB => Madd_n0000_inst_cy_2,
      SEL => cnt_2_GROM,
      O => cnt_2_CYMUXG
    );
  Madd_n0000_inst_sum_3 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_2,
      I1 => cnt_2_GROM,
      O => Q_n0000(3)
    );
  cnt_2_CYINIT_343 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_1,
      O => cnt_2_CYINIT
    );
  cnt_4_LOGIC_ZERO_344 : X_ZERO
    port map (
      O => cnt_4_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_4_345 : X_MUX2
    port map (
      IA => cnt_4_LOGIC_ZERO,
      IB => cnt_4_CYINIT,
      SEL => cnt_4_FROM,
      O => Madd_n0000_inst_cy_4
    );
  Madd_n0000_inst_sum_4 : X_XOR2
    port map (
      I0 => cnt_4_CYINIT,
      I1 => cnt_4_FROM,
      O => Q_n0000(4)
    );
  cnt_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_4_FROM
    );
  cnt_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(5),
      ADR3 => VCC,
      O => cnt_4_GROM
    );
  cnt_4_COUTUSED : X_BUF
    port map (
      I => cnt_4_CYMUXG,
      O => Madd_n0000_inst_cy_5
    );
  Madd_n0000_inst_cy_5_346 : X_MUX2
    port map (
      IA => cnt_4_LOGIC_ZERO,
      IB => Madd_n0000_inst_cy_4,
      SEL => cnt_4_GROM,
      O => cnt_4_CYMUXG
    );
  Madd_n0000_inst_sum_5 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_4,
      I1 => cnt_4_GROM,
      O => Q_n0000(5)
    );
  cnt_4_CYINIT_347 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_3,
      O => cnt_4_CYINIT
    );
  cnt_6_LOGIC_ZERO_348 : X_ZERO
    port map (
      O => cnt_6_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_6_349 : X_MUX2
    port map (
      IA => cnt_6_LOGIC_ZERO,
      IB => cnt_6_CYINIT,
      SEL => cnt_6_FROM,
      O => Madd_n0000_inst_cy_6
    );
  Madd_n0000_inst_sum_6 : X_XOR2
    port map (
      I0 => cnt_6_CYINIT,
      I1 => cnt_6_FROM,
      O => Q_n0000(6)
    );
  cnt_6_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_6_FROM
    );
  cnt_6_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(7),
      ADR3 => VCC,
      O => cnt_6_GROM
    );
  cnt_6_COUTUSED : X_BUF
    port map (
      I => cnt_6_CYMUXG,
      O => Madd_n0000_inst_cy_7
    );
  Madd_n0000_inst_cy_7_350 : X_MUX2
    port map (
      IA => cnt_6_LOGIC_ZERO,
      IB => Madd_n0000_inst_cy_6,
      SEL => cnt_6_GROM,
      O => cnt_6_CYMUXG
    );
  Madd_n0000_inst_sum_7 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_6,
      I1 => cnt_6_GROM,
      O => Q_n0000(7)
    );
  cnt_6_CYINIT_351 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_5,
      O => cnt_6_CYINIT
    );
  cnt_8_LOGIC_ZERO_352 : X_ZERO
    port map (
      O => cnt_8_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_8_353 : X_MUX2
    port map (
      IA => cnt_8_LOGIC_ZERO,
      IB => cnt_8_CYINIT,
      SEL => cnt_8_FROM,
      O => Madd_n0000_inst_cy_8
    );
  Madd_n0000_inst_sum_8 : X_XOR2
    port map (
      I0 => cnt_8_CYINIT,
      I1 => cnt_8_FROM,
      O => Q_n0000(8)
    );
  cnt_8_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_8_FROM
    );
  cnt_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(9),
      ADR3 => VCC,
      O => cnt_8_GROM
    );
  cnt_8_COUTUSED : X_BUF
    port map (
      I => cnt_8_CYMUXG,
      O => Madd_n0000_inst_cy_9
    );
  Madd_n0000_inst_cy_9_354 : X_MUX2
    port map (
      IA => cnt_8_LOGIC_ZERO,
      IB => Madd_n0000_inst_cy_8,
      SEL => cnt_8_GROM,
      O => cnt_8_CYMUXG
    );
  Madd_n0000_inst_sum_9 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_8,
      I1 => cnt_8_GROM,
      O => Q_n0000(9)
    );
  cnt_8_CYINIT_355 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_7,
      O => cnt_8_CYINIT
    );
  cnt_10_LOGIC_ZERO_356 : X_ZERO
    port map (
      O => cnt_10_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_10_357 : X_MUX2
    port map (
      IA => cnt_10_LOGIC_ZERO,
      IB => cnt_10_CYINIT,
      SEL => cnt_10_FROM,
      O => Madd_n0000_inst_cy_10
    );
  Madd_n0000_inst_sum_10 : X_XOR2
    port map (
      I0 => cnt_10_CYINIT,
      I1 => cnt_10_FROM,
      O => Q_n0000(10)
    );
  cnt_10_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_10_FROM
    );
  cnt_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(11),
      ADR3 => VCC,
      O => cnt_10_GROM
    );
  cnt_10_COUTUSED : X_BUF
    port map (
      I => cnt_10_CYMUXG,
      O => Madd_n0000_inst_cy_11
    );
  Madd_n0000_inst_cy_11_358 : X_MUX2
    port map (
      IA => cnt_10_LOGIC_ZERO,
      IB => Madd_n0000_inst_cy_10,
      SEL => cnt_10_GROM,
      O => cnt_10_CYMUXG
    );
  Madd_n0000_inst_sum_11 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_10,
      I1 => cnt_10_GROM,
      O => Q_n0000(11)
    );
  cnt_10_CYINIT_359 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_9,
      O => cnt_10_CYINIT
    );
  cnt_12_LOGIC_ZERO_360 : X_ZERO
    port map (
      O => cnt_12_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_12_361 : X_MUX2
    port map (
      IA => cnt_12_LOGIC_ZERO,
      IB => cnt_12_CYINIT,
      SEL => cnt_12_FROM,
      O => Madd_n0000_inst_cy_12
    );
  Madd_n0000_inst_sum_12 : X_XOR2
    port map (
      I0 => cnt_12_CYINIT,
      I1 => cnt_12_FROM,
      O => Q_n0000(12)
    );
  cnt_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_12_FROM
    );
  cnt_12_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(13),
      ADR3 => VCC,
      O => cnt_12_GROM
    );
  cnt_12_COUTUSED : X_BUF
    port map (
      I => cnt_12_CYMUXG,
      O => Madd_n0000_inst_cy_13
    );
  Madd_n0000_inst_cy_13_362 : X_MUX2
    port map (
      IA => cnt_12_LOGIC_ZERO,
      IB => Madd_n0000_inst_cy_12,
      SEL => cnt_12_GROM,
      O => cnt_12_CYMUXG
    );
  Madd_n0000_inst_sum_13 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_12,
      I1 => cnt_12_GROM,
      O => Q_n0000(13)
    );
  cnt_12_CYINIT_363 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_11,
      O => cnt_12_CYINIT
    );
  cnt_14_LOGIC_ZERO_364 : X_ZERO
    port map (
      O => cnt_14_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_14_365 : X_MUX2
    port map (
      IA => cnt_14_LOGIC_ZERO,
      IB => cnt_14_CYINIT,
      SEL => cnt_14_FROM,
      O => Madd_n0000_inst_cy_14
    );
  Madd_n0000_inst_sum_14 : X_XOR2
    port map (
      I0 => cnt_14_CYINIT,
      I1 => cnt_14_FROM,
      O => Q_n0000(14)
    );
  cnt_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_14_FROM
    );
  cnt_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(15),
      ADR3 => VCC,
      O => cnt_14_GROM
    );
  cnt_14_COUTUSED : X_BUF
    port map (
      I => cnt_14_CYMUXG,
      O => Madd_n0000_inst_cy_15
    );
  Madd_n0000_inst_cy_15_366 : X_MUX2
    port map (
      IA => cnt_14_LOGIC_ZERO,
      IB => Madd_n0000_inst_cy_14,
      SEL => cnt_14_GROM,
      O => cnt_14_CYMUXG
    );
  Madd_n0000_inst_sum_15 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_14,
      I1 => cnt_14_GROM,
      O => Q_n0000(15)
    );
  cnt_14_CYINIT_367 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_13,
      O => cnt_14_CYINIT
    );
  cnt_16_LOGIC_ZERO_368 : X_ZERO
    port map (
      O => cnt_16_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_16_369 : X_MUX2
    port map (
      IA => cnt_16_LOGIC_ZERO,
      IB => cnt_16_CYINIT,
      SEL => cnt_16_FROM,
      O => Madd_n0000_inst_cy_16
    );
  Madd_n0000_inst_sum_16 : X_XOR2
    port map (
      I0 => cnt_16_CYINIT,
      I1 => cnt_16_FROM,
      O => Q_n0000(16)
    );
  cnt_16_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_16_FROM
    );
  cnt_16_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(17),
      ADR3 => VCC,
      O => cnt_16_GROM
    );
  cnt_16_COUTUSED : X_BUF
    port map (
      I => cnt_16_CYMUXG,
      O => Madd_n0000_inst_cy_17
    );
  Madd_n0000_inst_cy_17_370 : X_MUX2
    port map (
      IA => cnt_16_LOGIC_ZERO,
      IB => Madd_n0000_inst_cy_16,
      SEL => cnt_16_GROM,
      O => cnt_16_CYMUXG
    );
  Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_16,
      I1 => cnt_16_GROM,
      O => Q_n0000(17)
    );
  cnt_16_CYINIT_371 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_15,
      O => cnt_16_CYINIT
    );
  cnt_18_LOGIC_ZERO_372 : X_ZERO
    port map (
      O => cnt_18_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_18_373 : X_MUX2
    port map (
      IA => cnt_18_LOGIC_ZERO,
      IB => cnt_18_CYINIT,
      SEL => cnt_18_FROM,
      O => Madd_n0000_inst_cy_18
    );
  Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => cnt_18_CYINIT,
      I1 => cnt_18_FROM,
      O => Q_n0000(18)
    );
  cnt_18_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_18_FROM
    );
  cnt_18_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(19),
      ADR3 => VCC,
      O => cnt_18_GROM
    );
  cnt_18_COUTUSED : X_BUF
    port map (
      I => cnt_18_CYMUXG,
      O => Madd_n0000_inst_cy_19
    );
  Madd_n0000_inst_cy_19_374 : X_MUX2
    port map (
      IA => cnt_18_LOGIC_ZERO,
      IB => Madd_n0000_inst_cy_18,
      SEL => cnt_18_GROM,
      O => cnt_18_CYMUXG
    );
  Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_18,
      I1 => cnt_18_GROM,
      O => Q_n0000(19)
    );
  cnt_18_CYINIT_375 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_17,
      O => cnt_18_CYINIT
    );
  cnt_20_LOGIC_ZERO_376 : X_ZERO
    port map (
      O => cnt_20_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_20_377 : X_MUX2
    port map (
      IA => cnt_20_LOGIC_ZERO,
      IB => cnt_20_CYINIT,
      SEL => cnt_20_FROM,
      O => Madd_n0000_inst_cy_20
    );
  Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => cnt_20_CYINIT,
      I1 => cnt_20_FROM,
      O => Q_n0000(20)
    );
  cnt_20_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(20),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_20_FROM
    );
  cnt_20_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(21),
      ADR3 => VCC,
      O => cnt_20_GROM
    );
  cnt_20_COUTUSED : X_BUF
    port map (
      I => cnt_20_CYMUXG,
      O => Madd_n0000_inst_cy_21
    );
  Madd_n0000_inst_cy_21_378 : X_MUX2
    port map (
      IA => cnt_20_LOGIC_ZERO,
      IB => Madd_n0000_inst_cy_20,
      SEL => cnt_20_GROM,
      O => cnt_20_CYMUXG
    );
  Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_20,
      I1 => cnt_20_GROM,
      O => Q_n0000(21)
    );
  cnt_20_CYINIT_379 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_19,
      O => cnt_20_CYINIT
    );
  cnt_22_LOGIC_ZERO_380 : X_ZERO
    port map (
      O => cnt_22_LOGIC_ZERO
    );
  Madd_n0000_inst_cy_22_381 : X_MUX2
    port map (
      IA => cnt_22_LOGIC_ZERO,
      IB => cnt_22_CYINIT,
      SEL => cnt_22_FROM,
      O => Madd_n0000_inst_cy_22
    );
  Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => cnt_22_CYINIT,
      I1 => cnt_22_FROM,
      O => Q_n0000(22)
    );
  cnt_22_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => cnt(22),
      ADR2 => VCC,
      ADR3 => VCC,
      O => cnt_22_FROM
    );
  cnt_23_rt_382 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => cnt(23),
      ADR3 => VCC,
      O => cnt_23_rt
    );
  cnt_22_YUSED : X_BUF
    port map (
      I => cnt_22_XORG,
      O => Q_n0000(23)
    );
  Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => Madd_n0000_inst_cy_22,
      I1 => cnt_23_rt,
      O => cnt_22_XORG
    );
  cnt_22_CYINIT_383 : X_BUF
    port map (
      I => Madd_n0000_inst_cy_21,
      O => cnt_22_CYINIT
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_0_LOGIC_ZERO_384 : X_ZERO
    port map (
      O => maccontrol_PHY_status_MII_Interface_mdccnt_0_LOGIC_ZERO
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_121_385 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_1,
      IB => maccontrol_PHY_status_MII_Interface_mdccnt_0_LOGIC_ZERO,
      SEL => maccontrol_PHY_status_MII_Interface_cs_FFd5_rt,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_121
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd5_rt_386 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd5_rt
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_01 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_61,
      ADR1 => VCC,
      ADR2 => maccontrol_PHY_status_MII_Interface_mdccnt(0),
      ADR3 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_0
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_0_COUTUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_0_CYMUXG,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_122
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_122_387 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_61,
      IB => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_121,
      SEL => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_0,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_0_CYMUXG
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_121_388 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_121,
      I1 => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_0,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_121
    );
  memcontroller_addr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_3_OD,
      CE => MA_3_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_3_OFF_RST,
      O => memcontroller_ADDREXT(3)
    );
  MA_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_3_OFF_RST
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_1_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_123,
      CE => maccontrol_PHY_status_MII_Interface_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_mdccnt_1_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_mdccnt(2)
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_1_LOGIC_ZERO_389 : X_ZERO
    port map (
      O => maccontrol_PHY_status_MII_Interface_mdccnt_1_LOGIC_ZERO
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_123_390 : X_MUX2
    port map (
      IA => maccontrol_PHY_status_MII_Interface_mdccnt_1_LOGIC_ZERO,
      IB => maccontrol_PHY_status_MII_Interface_mdccnt_1_CYINIT,
      SEL => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_1,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_123
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_122_391 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_mdccnt_1_CYINIT,
      I1 => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_1,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_122
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_11 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_MII_Interface_mdccnt(1),
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_1
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_21 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => VCC,
      ADR2 => maccontrol_PHY_status_MII_Interface_mdccnt(2),
      ADR3 => VCC,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_2
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_1_COUTUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_1_CYMUXG,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_124
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_124_392 : X_MUX2
    port map (
      IA => maccontrol_PHY_status_MII_Interface_mdccnt_1_LOGIC_ZERO,
      IB => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_123,
      SEL => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_2,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_1_CYMUXG
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_123_393 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_123,
      I1 => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_2,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_123
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_1_CYINIT_394 : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_122,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_1_CYINIT
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_3_LOGIC_ZERO_395 : X_ZERO
    port map (
      O => maccontrol_PHY_status_MII_Interface_mdccnt_3_LOGIC_ZERO
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_125_396 : X_MUX2
    port map (
      IA => maccontrol_PHY_status_MII_Interface_mdccnt_3_LOGIC_ZERO,
      IB => maccontrol_PHY_status_MII_Interface_mdccnt_3_CYINIT,
      SEL => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_3,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_125
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_124_397 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_mdccnt_3_CYINIT,
      I1 => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_3,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_124
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_31 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_mdccnt(3),
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_3
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_41 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => VCC,
      ADR2 => maccontrol_PHY_status_MII_Interface_mdccnt(4),
      ADR3 => VCC,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_4
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_3_COUTUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_3_CYMUXG,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_126
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_126_398 : X_MUX2
    port map (
      IA => maccontrol_PHY_status_MII_Interface_mdccnt_3_LOGIC_ZERO,
      IB => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_125,
      SEL => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_4,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_3_CYMUXG
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_125_399 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_125,
      I1 => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_4,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_125
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_3_CYINIT_400 : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_124,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_3_CYINIT
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_126_401 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_mdccnt_5_CYINIT,
      I1 => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_5,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_126
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_51 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_mdccnt(5),
      O => maccontrol_PHY_status_MII_Interface_mdccnt_inst_lut3_5
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd3_In_SW0 : X_LUT4
    generic map(
      INIT => X"CCFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_MII_Interface_mdccnt(5),
      ADR2 => VCC,
      ADR3 => MDC_OBUF,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_5_GROM
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_5_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_5_GROM,
      O => maccontrol_PHY_status_MII_Interface_N41734
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_5_CYINIT_402 : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_inst_cy_126,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_5_CYINIT
    );
  memtest_Mcompar_n0002_inst_cy_129_LOGIC_ONE_403 : X_ONE
    port map (
      O => memtest_Mcompar_n0002_inst_cy_129_LOGIC_ONE
    );
  memtest_Mcompar_n0002_inst_cy_129_LOGIC_ZERO_404 : X_ZERO
    port map (
      O => memtest_Mcompar_n0002_inst_cy_129_LOGIC_ZERO
    );
  memtest_Mcompar_n0002_inst_cy_128_405 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_129_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_129_LOGIC_ONE,
      SEL => memtest_Mcompar_n0002_inst_lut4_0,
      O => memtest_Mcompar_n0002_inst_cy_128
    );
  memtest_Mcompar_n0002_inst_lut4_01 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => q4(0),
      ADR1 => q4(1),
      ADR2 => memtest_Mshreg_dataw4_0_37,
      ADR3 => memtest_Mshreg_dataw4_1_36,
      O => memtest_Mcompar_n0002_inst_lut4_0
    );
  memtest_Mcompar_n0002_inst_lut4_16 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest_Mshreg_dataw4_3_34,
      ADR1 => q4(2),
      ADR2 => memtest_Mshreg_dataw4_2_35,
      ADR3 => q4(3),
      O => memtest_Mcompar_n0002_inst_lut4_1
    );
  memtest_Mcompar_n0002_inst_cy_129_COUTUSED : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_129_CYMUXG,
      O => memtest_Mcompar_n0002_inst_cy_129
    );
  memtest_Mcompar_n0002_inst_cy_129_406 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_129_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_128,
      SEL => memtest_Mcompar_n0002_inst_lut4_1,
      O => memtest_Mcompar_n0002_inst_cy_129_CYMUXG
    );
  memtest_Mcompar_n0002_inst_cy_131_LOGIC_ZERO_407 : X_ZERO
    port map (
      O => memtest_Mcompar_n0002_inst_cy_131_LOGIC_ZERO
    );
  memtest_Mcompar_n0002_inst_cy_130_408 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_131_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_131_CYINIT,
      SEL => memtest_Mcompar_n0002_inst_lut4_2,
      O => memtest_Mcompar_n0002_inst_cy_130
    );
  memtest_Mcompar_n0002_inst_lut4_21 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => memtest_Mshreg_dataw4_5_32,
      ADR1 => q4(5),
      ADR2 => q4(4),
      ADR3 => memtest_Mshreg_dataw4_4_33,
      O => memtest_Mcompar_n0002_inst_lut4_2
    );
  memtest_Mcompar_n0002_inst_lut4_31 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => q4(7),
      ADR1 => q4(6),
      ADR2 => memtest_Mshreg_dataw4_6_31,
      ADR3 => memtest_Mshreg_dataw4_7_30,
      O => memtest_Mcompar_n0002_inst_lut4_3
    );
  memtest_Mcompar_n0002_inst_cy_131_COUTUSED : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_131_CYMUXG,
      O => memtest_Mcompar_n0002_inst_cy_131
    );
  memtest_Mcompar_n0002_inst_cy_131_409 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_131_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_130,
      SEL => memtest_Mcompar_n0002_inst_lut4_3,
      O => memtest_Mcompar_n0002_inst_cy_131_CYMUXG
    );
  memtest_Mcompar_n0002_inst_cy_131_CYINIT_410 : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_129,
      O => memtest_Mcompar_n0002_inst_cy_131_CYINIT
    );
  memtest_Mcompar_n0002_inst_cy_133_LOGIC_ZERO_411 : X_ZERO
    port map (
      O => memtest_Mcompar_n0002_inst_cy_133_LOGIC_ZERO
    );
  memtest_Mcompar_n0002_inst_cy_132_412 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_133_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_133_CYINIT,
      SEL => memtest_Mcompar_n0002_inst_lut4_4,
      O => memtest_Mcompar_n0002_inst_cy_132
    );
  memtest_Mcompar_n0002_inst_lut4_41 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => q4(8),
      ADR1 => memtest_Mshreg_dataw4_9_28,
      ADR2 => q4(9),
      ADR3 => memtest_Mshreg_dataw4_8_29,
      O => memtest_Mcompar_n0002_inst_lut4_4
    );
  memtest_Mcompar_n0002_inst_lut4_51 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => q4(10),
      ADR1 => memtest_Mshreg_dataw4_11_26,
      ADR2 => memtest_Mshreg_dataw4_10_27,
      ADR3 => q4(11),
      O => memtest_Mcompar_n0002_inst_lut4_5
    );
  memtest_Mcompar_n0002_inst_cy_133_COUTUSED : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_133_CYMUXG,
      O => memtest_Mcompar_n0002_inst_cy_133
    );
  memtest_Mcompar_n0002_inst_cy_133_413 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_133_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_132,
      SEL => memtest_Mcompar_n0002_inst_lut4_5,
      O => memtest_Mcompar_n0002_inst_cy_133_CYMUXG
    );
  memtest_Mcompar_n0002_inst_cy_133_CYINIT_414 : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_131,
      O => memtest_Mcompar_n0002_inst_cy_133_CYINIT
    );
  memtest_Mcompar_n0002_inst_cy_135_LOGIC_ZERO_415 : X_ZERO
    port map (
      O => memtest_Mcompar_n0002_inst_cy_135_LOGIC_ZERO
    );
  memtest_Mcompar_n0002_inst_cy_134_416 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_135_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_135_CYINIT,
      SEL => memtest_Mcompar_n0002_inst_lut4_6,
      O => memtest_Mcompar_n0002_inst_cy_134
    );
  memtest_Mcompar_n0002_inst_lut4_61 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => q4(13),
      ADR1 => memtest_Mshreg_dataw4_12_25,
      ADR2 => q4(12),
      ADR3 => memtest_Mshreg_dataw4_13_24,
      O => memtest_Mcompar_n0002_inst_lut4_6
    );
  memtest_Mcompar_n0002_inst_lut4_71 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => memtest_Mshreg_dataw4_14_23,
      ADR1 => memtest_Mshreg_dataw4_15_22,
      ADR2 => q4(14),
      ADR3 => q4(15),
      O => memtest_Mcompar_n0002_inst_lut4_7
    );
  memtest_Mcompar_n0002_inst_cy_135_COUTUSED : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_135_CYMUXG,
      O => memtest_Mcompar_n0002_inst_cy_135
    );
  memtest_Mcompar_n0002_inst_cy_135_417 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_135_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_134,
      SEL => memtest_Mcompar_n0002_inst_lut4_7,
      O => memtest_Mcompar_n0002_inst_cy_135_CYMUXG
    );
  memtest_Mcompar_n0002_inst_cy_135_CYINIT_418 : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_133,
      O => memtest_Mcompar_n0002_inst_cy_135_CYINIT
    );
  memtest_Mcompar_n0002_inst_cy_137_LOGIC_ZERO_419 : X_ZERO
    port map (
      O => memtest_Mcompar_n0002_inst_cy_137_LOGIC_ZERO
    );
  memtest_Mcompar_n0002_inst_cy_136_420 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_137_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_137_CYINIT,
      SEL => memtest_Mcompar_n0002_inst_lut4_8,
      O => memtest_Mcompar_n0002_inst_cy_136
    );
  memtest_Mcompar_n0002_inst_lut4_81 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest_Mshreg_dataw4_16_21,
      ADR1 => memtest_Mshreg_dataw4_17_20,
      ADR2 => q4(17),
      ADR3 => q4(16),
      O => memtest_Mcompar_n0002_inst_lut4_8
    );
  memtest_Mcompar_n0002_inst_lut4_91 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => memtest_Mshreg_dataw4_19_18,
      ADR1 => q4(19),
      ADR2 => memtest_Mshreg_dataw4_18_19,
      ADR3 => q4(18),
      O => memtest_Mcompar_n0002_inst_lut4_9
    );
  memtest_Mcompar_n0002_inst_cy_137_COUTUSED : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_137_CYMUXG,
      O => memtest_Mcompar_n0002_inst_cy_137
    );
  memtest_Mcompar_n0002_inst_cy_137_421 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_137_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_136,
      SEL => memtest_Mcompar_n0002_inst_lut4_9,
      O => memtest_Mcompar_n0002_inst_cy_137_CYMUXG
    );
  memtest_Mcompar_n0002_inst_cy_137_CYINIT_422 : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_135,
      O => memtest_Mcompar_n0002_inst_cy_137_CYINIT
    );
  memtest_Mcompar_n0002_inst_cy_139_LOGIC_ZERO_423 : X_ZERO
    port map (
      O => memtest_Mcompar_n0002_inst_cy_139_LOGIC_ZERO
    );
  memtest_Mcompar_n0002_inst_cy_138_424 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_139_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_139_CYINIT,
      SEL => memtest_Mcompar_n0002_inst_lut4_10,
      O => memtest_Mcompar_n0002_inst_cy_138
    );
  memtest_Mcompar_n0002_inst_lut4_101 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => q4(20),
      ADR1 => memtest_Mshreg_dataw4_20_17,
      ADR2 => memtest_Mshreg_dataw4_21_16,
      ADR3 => q4(21),
      O => memtest_Mcompar_n0002_inst_lut4_10
    );
  memtest_Mcompar_n0002_inst_lut4_111 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => q4(22),
      ADR1 => memtest_Mshreg_dataw4_22_15,
      ADR2 => q4(23),
      ADR3 => memtest_Mshreg_dataw4_23_14,
      O => memtest_Mcompar_n0002_inst_lut4_11
    );
  memtest_Mcompar_n0002_inst_cy_139_COUTUSED : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_139_CYMUXG,
      O => memtest_Mcompar_n0002_inst_cy_139
    );
  memtest_Mcompar_n0002_inst_cy_139_425 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_139_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_138,
      SEL => memtest_Mcompar_n0002_inst_lut4_11,
      O => memtest_Mcompar_n0002_inst_cy_139_CYMUXG
    );
  memtest_Mcompar_n0002_inst_cy_139_CYINIT_426 : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_137,
      O => memtest_Mcompar_n0002_inst_cy_139_CYINIT
    );
  memtest_Mcompar_n0002_inst_cy_141_LOGIC_ZERO_427 : X_ZERO
    port map (
      O => memtest_Mcompar_n0002_inst_cy_141_LOGIC_ZERO
    );
  memtest_Mcompar_n0002_inst_cy_140_428 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_141_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_141_CYINIT,
      SEL => memtest_Mcompar_n0002_inst_lut4_12,
      O => memtest_Mcompar_n0002_inst_cy_140
    );
  memtest_Mcompar_n0002_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest_Mshreg_dataw4_24_13,
      ADR1 => memtest_Mshreg_dataw4_25_12,
      ADR2 => q4(25),
      ADR3 => q4(24),
      O => memtest_Mcompar_n0002_inst_lut4_12
    );
  memtest_Mcompar_n0002_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => memtest_Mshreg_dataw4_27_10,
      ADR1 => memtest_Mshreg_dataw4_26_11,
      ADR2 => q4(27),
      ADR3 => q4(26),
      O => memtest_Mcompar_n0002_inst_lut4_13
    );
  memtest_Mcompar_n0002_inst_cy_141_COUTUSED : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_141_CYMUXG,
      O => memtest_Mcompar_n0002_inst_cy_141
    );
  memtest_Mcompar_n0002_inst_cy_141_429 : X_MUX2
    port map (
      IA => memtest_Mcompar_n0002_inst_cy_141_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_140,
      SEL => memtest_Mcompar_n0002_inst_lut4_13,
      O => memtest_Mcompar_n0002_inst_cy_141_CYMUXG
    );
  memtest_Mcompar_n0002_inst_cy_141_CYINIT_430 : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_139,
      O => memtest_Mcompar_n0002_inst_cy_141_CYINIT
    );
  memtest_n0002_LOGIC_ZERO_431 : X_ZERO
    port map (
      O => memtest_n0002_LOGIC_ZERO
    );
  memtest_Mcompar_n0002_inst_cy_142_432 : X_MUX2
    port map (
      IA => memtest_n0002_LOGIC_ZERO,
      IB => memtest_n0002_CYINIT,
      SEL => memtest_Mcompar_n0002_inst_lut4_14,
      O => memtest_Mcompar_n0002_inst_cy_142
    );
  memtest_Mcompar_n0002_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => q4(28),
      ADR1 => memtest_Mshreg_dataw4_28_9,
      ADR2 => q4(29),
      ADR3 => memtest_Mshreg_dataw4_29_8,
      O => memtest_Mcompar_n0002_inst_lut4_14
    );
  memtest_Mcompar_n0002_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => q4(31),
      ADR1 => memtest_Mshreg_dataw4_31_6,
      ADR2 => q4(30),
      ADR3 => memtest_Mshreg_dataw4_30_7,
      O => memtest_Mcompar_n0002_inst_lut4_15
    );
  memtest_n0002_COUTUSED : X_BUF
    port map (
      I => memtest_n0002_CYMUXG,
      O => memtest_n0002
    );
  memtest_Mcompar_n0002_inst_cy_143 : X_MUX2
    port map (
      IA => memtest_n0002_LOGIC_ZERO,
      IB => memtest_Mcompar_n0002_inst_cy_142,
      SEL => memtest_Mcompar_n0002_inst_lut4_15,
      O => memtest_n0002_CYMUXG
    );
  memtest_n0002_CYINIT_433 : X_BUF
    port map (
      I => memtest_Mcompar_n0002_inst_cy_141,
      O => memtest_n0002_CYINIT
    );
  testrx_addr_0_LOGIC_ZERO_434 : X_ZERO
    port map (
      O => testrx_addr_0_LOGIC_ZERO
    );
  testrx_addr_Madd_n0000_inst_cy_30_435 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1,
      IB => testrx_addr_0_LOGIC_ZERO,
      SEL => testrx_addr_Madd_n0000_inst_lut2_30,
      O => testrx_addr_Madd_n0000_inst_cy_30
    );
  testrx_addr_Madd_n0000_inst_lut2_301 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1,
      ADR1 => VCC,
      ADR2 => testrx_addr(0),
      ADR3 => VCC,
      O => testrx_addr_Madd_n0000_inst_lut2_30
    );
  testrx_addr_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_67,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => testrx_addr(1),
      O => testrx_addr_0_GROM
    );
  testrx_addr_0_COUTUSED : X_BUF
    port map (
      I => testrx_addr_0_CYMUXG,
      O => testrx_addr_Madd_n0000_inst_cy_31
    );
  testrx_addr_Madd_n0000_inst_cy_31_436 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_67,
      IB => testrx_addr_Madd_n0000_inst_cy_30,
      SEL => testrx_addr_0_GROM,
      O => testrx_addr_0_CYMUXG
    );
  testrx_addr_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => testrx_addr_Madd_n0000_inst_cy_30,
      I1 => testrx_addr_0_GROM,
      O => testrx_addr_n0000(1)
    );
  testrx_addr_2_LOGIC_ZERO_437 : X_ZERO
    port map (
      O => testrx_addr_2_LOGIC_ZERO
    );
  testrx_addr_Madd_n0000_inst_cy_32_438 : X_MUX2
    port map (
      IA => testrx_addr_2_LOGIC_ZERO,
      IB => testrx_addr_2_CYINIT,
      SEL => testrx_addr_2_FROM,
      O => testrx_addr_Madd_n0000_inst_cy_32
    );
  testrx_addr_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => testrx_addr_2_CYINIT,
      I1 => testrx_addr_2_FROM,
      O => testrx_addr_n0000(2)
    );
  testrx_addr_2_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => testrx_addr(2),
      ADR3 => VCC,
      O => testrx_addr_2_FROM
    );
  testrx_addr_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => testrx_addr(3),
      O => testrx_addr_2_GROM
    );
  testrx_addr_2_COUTUSED : X_BUF
    port map (
      I => testrx_addr_2_CYMUXG,
      O => testrx_addr_Madd_n0000_inst_cy_33
    );
  testrx_addr_Madd_n0000_inst_cy_33_439 : X_MUX2
    port map (
      IA => testrx_addr_2_LOGIC_ZERO,
      IB => testrx_addr_Madd_n0000_inst_cy_32,
      SEL => testrx_addr_2_GROM,
      O => testrx_addr_2_CYMUXG
    );
  testrx_addr_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => testrx_addr_Madd_n0000_inst_cy_32,
      I1 => testrx_addr_2_GROM,
      O => testrx_addr_n0000(3)
    );
  testrx_addr_2_CYINIT_440 : X_BUF
    port map (
      I => testrx_addr_Madd_n0000_inst_cy_31,
      O => testrx_addr_2_CYINIT
    );
  testrx_addr_4_LOGIC_ZERO_441 : X_ZERO
    port map (
      O => testrx_addr_4_LOGIC_ZERO
    );
  testrx_addr_Madd_n0000_inst_cy_34_442 : X_MUX2
    port map (
      IA => testrx_addr_4_LOGIC_ZERO,
      IB => testrx_addr_4_CYINIT,
      SEL => testrx_addr_4_FROM,
      O => testrx_addr_Madd_n0000_inst_cy_34
    );
  testrx_addr_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => testrx_addr_4_CYINIT,
      I1 => testrx_addr_4_FROM,
      O => testrx_addr_n0000(4)
    );
  testrx_addr_4_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => testrx_addr(4),
      O => testrx_addr_4_FROM
    );
  testrx_addr_4_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => testrx_addr(5),
      O => testrx_addr_4_GROM
    );
  testrx_addr_4_COUTUSED : X_BUF
    port map (
      I => testrx_addr_4_CYMUXG,
      O => testrx_addr_Madd_n0000_inst_cy_35
    );
  testrx_addr_Madd_n0000_inst_cy_35_443 : X_MUX2
    port map (
      IA => testrx_addr_4_LOGIC_ZERO,
      IB => testrx_addr_Madd_n0000_inst_cy_34,
      SEL => testrx_addr_4_GROM,
      O => testrx_addr_4_CYMUXG
    );
  testrx_addr_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => testrx_addr_Madd_n0000_inst_cy_34,
      I1 => testrx_addr_4_GROM,
      O => testrx_addr_n0000(5)
    );
  testrx_addr_4_CYINIT_444 : X_BUF
    port map (
      I => testrx_addr_Madd_n0000_inst_cy_33,
      O => testrx_addr_4_CYINIT
    );
  testrx_addr_6_LOGIC_ZERO_445 : X_ZERO
    port map (
      O => testrx_addr_6_LOGIC_ZERO
    );
  testrx_addr_Madd_n0000_inst_cy_36_446 : X_MUX2
    port map (
      IA => testrx_addr_6_LOGIC_ZERO,
      IB => testrx_addr_6_CYINIT,
      SEL => testrx_addr_6_FROM,
      O => testrx_addr_Madd_n0000_inst_cy_36
    );
  testrx_addr_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => testrx_addr_6_CYINIT,
      I1 => testrx_addr_6_FROM,
      O => testrx_addr_n0000(6)
    );
  testrx_addr_6_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => testrx_addr(6),
      ADR3 => VCC,
      O => testrx_addr_6_FROM
    );
  testrx_addr_7_rt_447 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => testrx_addr(7),
      O => testrx_addr_7_rt
    );
  testrx_addr_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => testrx_addr_Madd_n0000_inst_cy_36,
      I1 => testrx_addr_7_rt,
      O => testrx_addr_n0000(7)
    );
  testrx_addr_6_CYINIT_448 : X_BUF
    port map (
      I => testrx_addr_Madd_n0000_inst_cy_35,
      O => testrx_addr_6_CYINIT
    );
  memtest2_cnt_0_LOGIC_ZERO_449 : X_ZERO
    port map (
      O => memtest2_cnt_0_LOGIC_ZERO
    );
  memtest2_cnt_Madd_n0000_inst_cy_86_450 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_16,
      IB => memtest2_cnt_0_LOGIC_ZERO,
      SEL => memtest2_cnt_Madd_n0000_inst_lut2_86,
      O => memtest2_cnt_Madd_n0000_inst_cy_86
    );
  memtest2_cnt_Madd_n0000_inst_lut2_861 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_16,
      ADR1 => memtest2_cnt(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_cnt_Madd_n0000_inst_lut2_86
    );
  memtest2_cnt_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_52,
      ADR1 => VCC,
      ADR2 => memtest2_cnt(1),
      ADR3 => VCC,
      O => memtest2_cnt_0_GROM
    );
  memtest2_cnt_0_COUTUSED : X_BUF
    port map (
      I => memtest2_cnt_0_CYMUXG,
      O => memtest2_cnt_Madd_n0000_inst_cy_87
    );
  memtest2_cnt_Madd_n0000_inst_cy_87_451 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_52,
      IB => memtest2_cnt_Madd_n0000_inst_cy_86,
      SEL => memtest2_cnt_0_GROM,
      O => memtest2_cnt_0_CYMUXG
    );
  memtest2_cnt_Madd_n0000_inst_sum_87 : X_XOR2
    port map (
      I0 => memtest2_cnt_Madd_n0000_inst_cy_86,
      I1 => memtest2_cnt_0_GROM,
      O => memtest2_cnt_n0000(1)
    );
  memtest2_cnt_2_LOGIC_ZERO_452 : X_ZERO
    port map (
      O => memtest2_cnt_2_LOGIC_ZERO
    );
  memtest2_cnt_Madd_n0000_inst_cy_88_453 : X_MUX2
    port map (
      IA => memtest2_cnt_2_LOGIC_ZERO,
      IB => memtest2_cnt_2_CYINIT,
      SEL => memtest2_cnt_2_FROM,
      O => memtest2_cnt_Madd_n0000_inst_cy_88
    );
  memtest2_cnt_Madd_n0000_inst_sum_88 : X_XOR2
    port map (
      I0 => memtest2_cnt_2_CYINIT,
      I1 => memtest2_cnt_2_FROM,
      O => memtest2_cnt_n0000(2)
    );
  memtest2_cnt_2_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memtest2_cnt(2),
      ADR3 => VCC,
      O => memtest2_cnt_2_FROM
    );
  memtest2_cnt_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memtest2_cnt(3),
      ADR3 => VCC,
      O => memtest2_cnt_2_GROM
    );
  memtest2_cnt_2_COUTUSED : X_BUF
    port map (
      I => memtest2_cnt_2_CYMUXG,
      O => memtest2_cnt_Madd_n0000_inst_cy_89
    );
  memtest2_cnt_Madd_n0000_inst_cy_89_454 : X_MUX2
    port map (
      IA => memtest2_cnt_2_LOGIC_ZERO,
      IB => memtest2_cnt_Madd_n0000_inst_cy_88,
      SEL => memtest2_cnt_2_GROM,
      O => memtest2_cnt_2_CYMUXG
    );
  memtest2_cnt_Madd_n0000_inst_sum_89 : X_XOR2
    port map (
      I0 => memtest2_cnt_Madd_n0000_inst_cy_88,
      I1 => memtest2_cnt_2_GROM,
      O => memtest2_cnt_n0000(3)
    );
  memtest2_cnt_2_CYINIT_455 : X_BUF
    port map (
      I => memtest2_cnt_Madd_n0000_inst_cy_87,
      O => memtest2_cnt_2_CYINIT
    );
  memtest2_cnt_4_LOGIC_ZERO_456 : X_ZERO
    port map (
      O => memtest2_cnt_4_LOGIC_ZERO
    );
  memtest2_cnt_Madd_n0000_inst_cy_90_457 : X_MUX2
    port map (
      IA => memtest2_cnt_4_LOGIC_ZERO,
      IB => memtest2_cnt_4_CYINIT,
      SEL => memtest2_cnt_4_FROM,
      O => memtest2_cnt_Madd_n0000_inst_cy_90
    );
  memtest2_cnt_Madd_n0000_inst_sum_90 : X_XOR2
    port map (
      I0 => memtest2_cnt_4_CYINIT,
      I1 => memtest2_cnt_4_FROM,
      O => memtest2_cnt_n0000(4)
    );
  memtest2_cnt_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_cnt_4_FROM
    );
  memtest2_cnt_4_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => memtest2_cnt(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_cnt_4_GROM
    );
  memtest2_cnt_4_COUTUSED : X_BUF
    port map (
      I => memtest2_cnt_4_CYMUXG,
      O => memtest2_cnt_Madd_n0000_inst_cy_91
    );
  memtest2_cnt_Madd_n0000_inst_cy_91_458 : X_MUX2
    port map (
      IA => memtest2_cnt_4_LOGIC_ZERO,
      IB => memtest2_cnt_Madd_n0000_inst_cy_90,
      SEL => memtest2_cnt_4_GROM,
      O => memtest2_cnt_4_CYMUXG
    );
  memtest2_cnt_Madd_n0000_inst_sum_91 : X_XOR2
    port map (
      I0 => memtest2_cnt_Madd_n0000_inst_cy_90,
      I1 => memtest2_cnt_4_GROM,
      O => memtest2_cnt_n0000(5)
    );
  memtest2_cnt_4_CYINIT_459 : X_BUF
    port map (
      I => memtest2_cnt_Madd_n0000_inst_cy_89,
      O => memtest2_cnt_4_CYINIT
    );
  memtest2_cnt_6_LOGIC_ZERO_460 : X_ZERO
    port map (
      O => memtest2_cnt_6_LOGIC_ZERO
    );
  memtest2_cnt_Madd_n0000_inst_cy_92_461 : X_MUX2
    port map (
      IA => memtest2_cnt_6_LOGIC_ZERO,
      IB => memtest2_cnt_6_CYINIT,
      SEL => memtest2_cnt_6_FROM,
      O => memtest2_cnt_Madd_n0000_inst_cy_92
    );
  memtest2_cnt_Madd_n0000_inst_sum_92 : X_XOR2
    port map (
      I0 => memtest2_cnt_6_CYINIT,
      I1 => memtest2_cnt_6_FROM,
      O => memtest2_cnt_n0000(6)
    );
  memtest2_cnt_6_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => memtest2_cnt(6),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_cnt_6_FROM
    );
  memtest2_cnt_6_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memtest2_cnt(7),
      ADR3 => VCC,
      O => memtest2_cnt_6_GROM
    );
  memtest2_cnt_6_COUTUSED : X_BUF
    port map (
      I => memtest2_cnt_6_CYMUXG,
      O => memtest2_cnt_Madd_n0000_inst_cy_93
    );
  memtest2_cnt_Madd_n0000_inst_cy_93_462 : X_MUX2
    port map (
      IA => memtest2_cnt_6_LOGIC_ZERO,
      IB => memtest2_cnt_Madd_n0000_inst_cy_92,
      SEL => memtest2_cnt_6_GROM,
      O => memtest2_cnt_6_CYMUXG
    );
  memtest2_cnt_Madd_n0000_inst_sum_93 : X_XOR2
    port map (
      I0 => memtest2_cnt_Madd_n0000_inst_cy_92,
      I1 => memtest2_cnt_6_GROM,
      O => memtest2_cnt_n0000(7)
    );
  memtest2_cnt_6_CYINIT_463 : X_BUF
    port map (
      I => memtest2_cnt_Madd_n0000_inst_cy_91,
      O => memtest2_cnt_6_CYINIT
    );
  memcontroller_addr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_4_OD,
      CE => MA_4_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_4_OFF_RST,
      O => memcontroller_ADDREXT(4)
    );
  MA_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_4_OFF_RST
    );
  memtest2_cnt_8_LOGIC_ZERO_464 : X_ZERO
    port map (
      O => memtest2_cnt_8_LOGIC_ZERO
    );
  memtest2_cnt_Madd_n0000_inst_cy_94_465 : X_MUX2
    port map (
      IA => memtest2_cnt_8_LOGIC_ZERO,
      IB => memtest2_cnt_8_CYINIT,
      SEL => memtest2_cnt_8_FROM,
      O => memtest2_cnt_Madd_n0000_inst_cy_94
    );
  memtest2_cnt_Madd_n0000_inst_sum_94 : X_XOR2
    port map (
      I0 => memtest2_cnt_8_CYINIT,
      I1 => memtest2_cnt_8_FROM,
      O => memtest2_cnt_n0000(8)
    );
  memtest2_cnt_8_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_cnt_8_FROM
    );
  memtest2_cnt_8_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memtest2_cnt(9),
      O => memtest2_cnt_8_GROM
    );
  memtest2_cnt_8_COUTUSED : X_BUF
    port map (
      I => memtest2_cnt_8_CYMUXG,
      O => memtest2_cnt_Madd_n0000_inst_cy_95
    );
  memtest2_cnt_Madd_n0000_inst_cy_95_466 : X_MUX2
    port map (
      IA => memtest2_cnt_8_LOGIC_ZERO,
      IB => memtest2_cnt_Madd_n0000_inst_cy_94,
      SEL => memtest2_cnt_8_GROM,
      O => memtest2_cnt_8_CYMUXG
    );
  memtest2_cnt_Madd_n0000_inst_sum_95 : X_XOR2
    port map (
      I0 => memtest2_cnt_Madd_n0000_inst_cy_94,
      I1 => memtest2_cnt_8_GROM,
      O => memtest2_cnt_n0000(9)
    );
  memtest2_cnt_8_CYINIT_467 : X_BUF
    port map (
      I => memtest2_cnt_Madd_n0000_inst_cy_93,
      O => memtest2_cnt_8_CYINIT
    );
  memtest2_cnt_10_LOGIC_ZERO_468 : X_ZERO
    port map (
      O => memtest2_cnt_10_LOGIC_ZERO
    );
  memtest2_cnt_Madd_n0000_inst_cy_96_469 : X_MUX2
    port map (
      IA => memtest2_cnt_10_LOGIC_ZERO,
      IB => memtest2_cnt_10_CYINIT,
      SEL => memtest2_cnt_10_FROM,
      O => memtest2_cnt_Madd_n0000_inst_cy_96
    );
  memtest2_cnt_Madd_n0000_inst_sum_96 : X_XOR2
    port map (
      I0 => memtest2_cnt_10_CYINIT,
      I1 => memtest2_cnt_10_FROM,
      O => memtest2_cnt_n0000(10)
    );
  memtest2_cnt_10_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_cnt_10_FROM
    );
  memtest2_cnt_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memtest2_cnt(11),
      O => memtest2_cnt_10_GROM
    );
  memtest2_cnt_10_COUTUSED : X_BUF
    port map (
      I => memtest2_cnt_10_CYMUXG,
      O => memtest2_cnt_Madd_n0000_inst_cy_97
    );
  memtest2_cnt_Madd_n0000_inst_cy_97_470 : X_MUX2
    port map (
      IA => memtest2_cnt_10_LOGIC_ZERO,
      IB => memtest2_cnt_Madd_n0000_inst_cy_96,
      SEL => memtest2_cnt_10_GROM,
      O => memtest2_cnt_10_CYMUXG
    );
  memtest2_cnt_Madd_n0000_inst_sum_97 : X_XOR2
    port map (
      I0 => memtest2_cnt_Madd_n0000_inst_cy_96,
      I1 => memtest2_cnt_10_GROM,
      O => memtest2_cnt_n0000(11)
    );
  memtest2_cnt_10_CYINIT_471 : X_BUF
    port map (
      I => memtest2_cnt_Madd_n0000_inst_cy_95,
      O => memtest2_cnt_10_CYINIT
    );
  memtest2_cnt_12_LOGIC_ZERO_472 : X_ZERO
    port map (
      O => memtest2_cnt_12_LOGIC_ZERO
    );
  memtest2_cnt_Madd_n0000_inst_cy_98_473 : X_MUX2
    port map (
      IA => memtest2_cnt_12_LOGIC_ZERO,
      IB => memtest2_cnt_12_CYINIT,
      SEL => memtest2_cnt_12_FROM,
      O => memtest2_cnt_Madd_n0000_inst_cy_98
    );
  memtest2_cnt_Madd_n0000_inst_sum_98 : X_XOR2
    port map (
      I0 => memtest2_cnt_12_CYINIT,
      I1 => memtest2_cnt_12_FROM,
      O => memtest2_cnt_n0000(12)
    );
  memtest2_cnt_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_cnt_12_FROM
    );
  memtest2_cnt_12_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memtest2_cnt(13),
      O => memtest2_cnt_12_GROM
    );
  memtest2_cnt_12_COUTUSED : X_BUF
    port map (
      I => memtest2_cnt_12_CYMUXG,
      O => memtest2_cnt_Madd_n0000_inst_cy_99
    );
  memtest2_cnt_Madd_n0000_inst_cy_99_474 : X_MUX2
    port map (
      IA => memtest2_cnt_12_LOGIC_ZERO,
      IB => memtest2_cnt_Madd_n0000_inst_cy_98,
      SEL => memtest2_cnt_12_GROM,
      O => memtest2_cnt_12_CYMUXG
    );
  memtest2_cnt_Madd_n0000_inst_sum_99 : X_XOR2
    port map (
      I0 => memtest2_cnt_Madd_n0000_inst_cy_98,
      I1 => memtest2_cnt_12_GROM,
      O => memtest2_cnt_n0000(13)
    );
  memtest2_cnt_12_CYINIT_475 : X_BUF
    port map (
      I => memtest2_cnt_Madd_n0000_inst_cy_97,
      O => memtest2_cnt_12_CYINIT
    );
  memtest2_cnt_14_LOGIC_ZERO_476 : X_ZERO
    port map (
      O => memtest2_cnt_14_LOGIC_ZERO
    );
  memtest2_cnt_Madd_n0000_inst_cy_100_477 : X_MUX2
    port map (
      IA => memtest2_cnt_14_LOGIC_ZERO,
      IB => memtest2_cnt_14_CYINIT,
      SEL => memtest2_cnt_14_FROM,
      O => memtest2_cnt_Madd_n0000_inst_cy_100
    );
  memtest2_cnt_Madd_n0000_inst_sum_100 : X_XOR2
    port map (
      I0 => memtest2_cnt_14_CYINIT,
      I1 => memtest2_cnt_14_FROM,
      O => memtest2_cnt_n0000(14)
    );
  memtest2_cnt_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_cnt_14_FROM
    );
  memtest2_cnt_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memtest2_cnt(15),
      ADR3 => VCC,
      O => memtest2_cnt_14_GROM
    );
  memtest2_cnt_14_COUTUSED : X_BUF
    port map (
      I => memtest2_cnt_14_CYMUXG,
      O => memtest2_cnt_Madd_n0000_inst_cy_101
    );
  memtest2_cnt_Madd_n0000_inst_cy_101_478 : X_MUX2
    port map (
      IA => memtest2_cnt_14_LOGIC_ZERO,
      IB => memtest2_cnt_Madd_n0000_inst_cy_100,
      SEL => memtest2_cnt_14_GROM,
      O => memtest2_cnt_14_CYMUXG
    );
  memtest2_cnt_Madd_n0000_inst_sum_101 : X_XOR2
    port map (
      I0 => memtest2_cnt_Madd_n0000_inst_cy_100,
      I1 => memtest2_cnt_14_GROM,
      O => memtest2_cnt_n0000(15)
    );
  memtest2_cnt_14_CYINIT_479 : X_BUF
    port map (
      I => memtest2_cnt_Madd_n0000_inst_cy_99,
      O => memtest2_cnt_14_CYINIT
    );
  memtest2_cnt_Madd_n0000_inst_sum_102 : X_XOR2
    port map (
      I0 => memtest2_cnt_16_CYINIT,
      I1 => memtest2_cnt_16_rt,
      O => memtest2_cnt_n0000(16)
    );
  memtest2_cnt_16_rt_480 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_cnt_16_rt
    );
  memtest2_cnt_16_CYINIT_481 : X_BUF
    port map (
      I => memtest2_cnt_Madd_n0000_inst_cy_101,
      O => memtest2_cnt_16_CYINIT
    );
  memtest2_Mcompar_n0025_inst_cy_161_LOGIC_ONE_482 : X_ONE
    port map (
      O => memtest2_Mcompar_n0025_inst_cy_161_LOGIC_ONE
    );
  memtest2_Mcompar_n0025_inst_cy_161_LOGIC_ZERO_483 : X_ZERO
    port map (
      O => memtest2_Mcompar_n0025_inst_cy_161_LOGIC_ZERO
    );
  memtest2_Mcompar_n0025_inst_cy_160_484 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0025_inst_cy_161_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0025_inst_cy_161_LOGIC_ONE,
      SEL => memtest2_Mcompar_n0025_inst_lut4_22,
      O => memtest2_Mcompar_n0025_inst_cy_160
    );
  memtest2_Mcompar_n0025_inst_lut4_221 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(4),
      ADR1 => memtest2_cnt(3),
      ADR2 => memtest2_cnt(1),
      ADR3 => memtest2_cnt(2),
      O => memtest2_Mcompar_n0025_inst_lut4_22
    );
  memtest2_Mcompar_n0025_inst_lut4_231 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(7),
      ADR1 => memtest2_cnt(5),
      ADR2 => memtest2_cnt(6),
      ADR3 => memtest2_cnt(8),
      O => memtest2_Mcompar_n0025_inst_lut4_23
    );
  memtest2_Mcompar_n0025_inst_cy_161_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0025_inst_cy_161_CYMUXG,
      O => memtest2_Mcompar_n0025_inst_cy_161
    );
  memtest2_Mcompar_n0025_inst_cy_161_485 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0025_inst_cy_161_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0025_inst_cy_160,
      SEL => memtest2_Mcompar_n0025_inst_lut4_23,
      O => memtest2_Mcompar_n0025_inst_cy_161_CYMUXG
    );
  memtest2_Mcompar_n0025_inst_cy_163_LOGIC_ZERO_486 : X_ZERO
    port map (
      O => memtest2_Mcompar_n0025_inst_cy_163_LOGIC_ZERO
    );
  memtest2_Mcompar_n0025_inst_cy_162_487 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0025_inst_cy_163_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0025_inst_cy_163_CYINIT,
      SEL => memtest2_Mcompar_n0025_inst_lut4_24,
      O => memtest2_Mcompar_n0025_inst_cy_162
    );
  memtest2_Mcompar_n0025_inst_lut4_241 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(10),
      ADR1 => memtest2_cnt(12),
      ADR2 => memtest2_cnt(9),
      ADR3 => memtest2_cnt(11),
      O => memtest2_Mcompar_n0025_inst_lut4_24
    );
  memtest2_Mcompar_n0025_inst_lut3_61 : X_LUT4
    generic map(
      INIT => X"0003"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(14),
      ADR2 => memtest2_cnt(15),
      ADR3 => memtest2_cnt(13),
      O => memtest2_Mcompar_n0025_inst_lut3_6
    );
  memtest2_Mcompar_n0025_inst_cy_163_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0025_inst_cy_163_CYMUXG,
      O => memtest2_Mcompar_n0025_inst_cy_163
    );
  memtest2_Mcompar_n0025_inst_cy_163_488 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0025_inst_cy_163_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0025_inst_cy_162,
      SEL => memtest2_Mcompar_n0025_inst_lut3_6,
      O => memtest2_Mcompar_n0025_inst_cy_163_CYMUXG
    );
  memtest2_Mcompar_n0025_inst_cy_163_CYINIT_489 : X_BUF
    port map (
      I => memtest2_Mcompar_n0025_inst_cy_161,
      O => memtest2_Mcompar_n0025_inst_cy_163_CYINIT
    );
  memtest2_n0025_LOGIC_ONE_490 : X_ONE
    port map (
      O => memtest2_n0025_LOGIC_ONE
    );
  memtest2_Mcompar_n0025_inst_cy_164_491 : X_MUX2
    port map (
      IA => memtest2_n0025_LOGIC_ONE,
      IB => memtest2_n0025_CYINIT,
      SEL => memtest2_SIG_0,
      O => memtest2_Mcompar_n0025_inst_cy_164
    );
  memtest2_BEL_0 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memtest2_cnt(16),
      O => memtest2_SIG_0
    );
  memtest2_BEL_1 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_SIG_1
    );
  memtest2_n0025_COUTUSED : X_BUF
    port map (
      I => memtest2_n0025_CYMUXG,
      O => memtest2_n0025
    );
  memtest2_Mcompar_n0025_inst_cy_165 : X_MUX2
    port map (
      IA => memtest2_n0025_LOGIC_ONE,
      IB => memtest2_Mcompar_n0025_inst_cy_164,
      SEL => memtest2_SIG_1,
      O => memtest2_n0025_CYMUXG
    );
  memtest2_n0025_CYINIT_492 : X_BUF
    port map (
      I => memtest2_Mcompar_n0025_inst_cy_163,
      O => memtest2_n0025_CYINIT
    );
  memtest2_Mcompar_n0017_inst_cy_167_LOGIC_ONE_493 : X_ONE
    port map (
      O => memtest2_Mcompar_n0017_inst_cy_167_LOGIC_ONE
    );
  memtest2_Mcompar_n0017_inst_cy_167_LOGIC_ZERO_494 : X_ZERO
    port map (
      O => memtest2_Mcompar_n0017_inst_cy_167_LOGIC_ZERO
    );
  memtest2_Mcompar_n0017_inst_cy_166_495 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0017_inst_cy_167_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0017_inst_cy_167_LOGIC_ONE,
      SEL => memtest2_Mcompar_n0017_inst_lut4_25,
      O => memtest2_Mcompar_n0017_inst_cy_166
    );
  memtest2_Mcompar_n0017_inst_lut4_251 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => memtest2_Mshreg_data4_1_68,
      ADR1 => memtest2_datain(0),
      ADR2 => memtest2_datain(1),
      ADR3 => memtest2_Mshreg_data4_0_69,
      O => memtest2_Mcompar_n0017_inst_lut4_25
    );
  memtest2_Mcompar_n0017_inst_lut4_261 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest2_Mshreg_data4_2_67,
      ADR1 => memtest2_Mshreg_data4_3_66,
      ADR2 => memtest2_datain(3),
      ADR3 => memtest2_datain(2),
      O => memtest2_Mcompar_n0017_inst_lut4_26
    );
  memtest2_Mcompar_n0017_inst_cy_167_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0017_inst_cy_167_CYMUXG,
      O => memtest2_Mcompar_n0017_inst_cy_167
    );
  memtest2_Mcompar_n0017_inst_cy_167_496 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0017_inst_cy_167_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0017_inst_cy_166,
      SEL => memtest2_Mcompar_n0017_inst_lut4_26,
      O => memtest2_Mcompar_n0017_inst_cy_167_CYMUXG
    );
  memtest2_deq_0_LOGIC_ZERO_497 : X_ZERO
    port map (
      O => memtest2_deq_0_LOGIC_ZERO
    );
  memtest2_Mcompar_n0017_inst_cy_168_498 : X_MUX2
    port map (
      IA => memtest2_deq_0_LOGIC_ZERO,
      IB => memtest2_deq_0_CYINIT,
      SEL => memtest2_Mcompar_n0017_inst_lut4_27,
      O => memtest2_Mcompar_n0017_inst_cy_168
    );
  memtest2_Mcompar_n0017_inst_lut4_271 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => memtest2_Mshreg_data4_4_65,
      ADR1 => memtest2_Mshreg_data4_5_64,
      ADR2 => memtest2_datain(4),
      ADR3 => memtest2_datain(5),
      O => memtest2_Mcompar_n0017_inst_lut4_27
    );
  memtest2_Mcompar_n0017_inst_lut4_281 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest2_Mshreg_data4_6_63,
      ADR1 => memtest2_Mshreg_data4_7_62,
      ADR2 => memtest2_datain(7),
      ADR3 => memtest2_datain(6),
      O => memtest2_Mcompar_n0017_inst_lut4_28
    );
  memtest2_deq_0_COUTUSED : X_BUF
    port map (
      I => memtest2_deq_0_CYMUXG,
      O => memtest2_deq(0)
    );
  memtest2_Mcompar_n0017_inst_cy_169 : X_MUX2
    port map (
      IA => memtest2_deq_0_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0017_inst_cy_168,
      SEL => memtest2_Mcompar_n0017_inst_lut4_28,
      O => memtest2_deq_0_CYMUXG
    );
  memtest2_deq_0_CYINIT_499 : X_BUF
    port map (
      I => memtest2_Mcompar_n0017_inst_cy_167,
      O => memtest2_deq_0_CYINIT
    );
  maccontrol_PHY_status_MII_Interface_n0078_1_LOGIC_ZERO_500 : X_ZERO
    port map (
      O => maccontrol_PHY_status_MII_Interface_n0078_1_LOGIC_ZERO
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_24_501 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_2,
      IB => maccontrol_PHY_status_MII_Interface_n0078_1_LOGIC_ZERO,
      SEL => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_lut2_24,
      O => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_24
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_lut2_241 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(0),
      O => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_lut2_24
    );
  maccontrol_PHY_status_MII_Interface_n0078_1_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_60,
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => maccontrol_PHY_status_MII_Interface_n0078_1_GROM
    );
  maccontrol_PHY_status_MII_Interface_n0078_1_COUTUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0078_1_CYMUXG,
      O => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_25
    );
  maccontrol_PHY_status_MII_Interface_n0078_1_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0078_1_XORG,
      O => maccontrol_PHY_status_MII_Interface_n0078(1)
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_25_502 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_60,
      IB => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_24,
      SEL => maccontrol_PHY_status_MII_Interface_n0078_1_GROM,
      O => maccontrol_PHY_status_MII_Interface_n0078_1_CYMUXG
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_sum_25 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_24,
      I1 => maccontrol_PHY_status_MII_Interface_n0078_1_GROM,
      O => maccontrol_PHY_status_MII_Interface_n0078_1_XORG
    );
  maccontrol_PHY_status_MII_Interface_n0078_2_LOGIC_ZERO_503 : X_ZERO
    port map (
      O => maccontrol_PHY_status_MII_Interface_n0078_2_LOGIC_ZERO
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_26_504 : X_MUX2
    port map (
      IA => maccontrol_PHY_status_MII_Interface_n0078_2_LOGIC_ZERO,
      IB => maccontrol_PHY_status_MII_Interface_n0078_2_CYINIT,
      SEL => maccontrol_PHY_status_MII_Interface_n0078_2_FROM,
      O => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_26
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_sum_26 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_n0078_2_CYINIT,
      I1 => maccontrol_PHY_status_MII_Interface_n0078_2_FROM,
      O => maccontrol_PHY_status_MII_Interface_n0078_2_XORF
    );
  maccontrol_PHY_status_MII_Interface_n0078_2_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => maccontrol_PHY_status_MII_Interface_n0078_2_FROM
    );
  maccontrol_PHY_status_MII_Interface_n0078_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      O => maccontrol_PHY_status_MII_Interface_n0078_2_GROM
    );
  maccontrol_PHY_status_MII_Interface_n0078_2_COUTUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0078_2_CYMUXG,
      O => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_27
    );
  maccontrol_PHY_status_MII_Interface_n0078_2_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0078_2_XORF,
      O => maccontrol_PHY_status_MII_Interface_n0078(2)
    );
  maccontrol_PHY_status_MII_Interface_n0078_2_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0078_2_XORG,
      O => maccontrol_PHY_status_MII_Interface_n0078(3)
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_27_505 : X_MUX2
    port map (
      IA => maccontrol_PHY_status_MII_Interface_n0078_2_LOGIC_ZERO,
      IB => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_26,
      SEL => maccontrol_PHY_status_MII_Interface_n0078_2_GROM,
      O => maccontrol_PHY_status_MII_Interface_n0078_2_CYMUXG
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_sum_27 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_26,
      I1 => maccontrol_PHY_status_MII_Interface_n0078_2_GROM,
      O => maccontrol_PHY_status_MII_Interface_n0078_2_XORG
    );
  maccontrol_PHY_status_MII_Interface_n0078_2_CYINIT_506 : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_25,
      O => maccontrol_PHY_status_MII_Interface_n0078_2_CYINIT
    );
  maccontrol_PHY_status_MII_Interface_n0078_4_LOGIC_ZERO_507 : X_ZERO
    port map (
      O => maccontrol_PHY_status_MII_Interface_n0078_4_LOGIC_ZERO
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_28_508 : X_MUX2
    port map (
      IA => maccontrol_PHY_status_MII_Interface_n0078_4_LOGIC_ZERO,
      IB => maccontrol_PHY_status_MII_Interface_n0078_4_CYINIT,
      SEL => maccontrol_PHY_status_MII_Interface_n0078_4_FROM,
      O => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_28
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_sum_28 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_n0078_4_CYINIT,
      I1 => maccontrol_PHY_status_MII_Interface_n0078_4_FROM,
      O => maccontrol_PHY_status_MII_Interface_n0078_4_XORF
    );
  maccontrol_PHY_status_MII_Interface_n0078_4_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR3 => VCC,
      O => maccontrol_PHY_status_MII_Interface_n0078_4_FROM
    );
  maccontrol_PHY_status_MII_Interface_statecnt_5_rt_509 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(5),
      O => maccontrol_PHY_status_MII_Interface_statecnt_5_rt
    );
  maccontrol_PHY_status_MII_Interface_n0078_4_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0078_4_XORF,
      O => maccontrol_PHY_status_MII_Interface_n0078(4)
    );
  maccontrol_PHY_status_MII_Interface_n0078_4_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0078_4_XORG,
      O => maccontrol_PHY_status_MII_Interface_n0078(5)
    );
  maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_sum_29 : X_XOR2
    port map (
      I0 => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_28,
      I1 => maccontrol_PHY_status_MII_Interface_statecnt_5_rt,
      O => maccontrol_PHY_status_MII_Interface_n0078_4_XORG
    );
  maccontrol_PHY_status_MII_Interface_n0078_4_CYINIT_510 : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_Madd_n0078_inst_cy_27,
      O => maccontrol_PHY_status_MII_Interface_n0078_4_CYINIT
    );
  memtest2_Mcompar_n0018_inst_cy_167_LOGIC_ONE_511 : X_ONE
    port map (
      O => memtest2_Mcompar_n0018_inst_cy_167_LOGIC_ONE
    );
  memtest2_Mcompar_n0018_inst_cy_167_LOGIC_ZERO_512 : X_ZERO
    port map (
      O => memtest2_Mcompar_n0018_inst_cy_167_LOGIC_ZERO
    );
  memtest2_Mcompar_n0018_inst_cy_166_513 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0018_inst_cy_167_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0018_inst_cy_167_LOGIC_ONE,
      SEL => memtest2_Mcompar_n0018_inst_lut4_25,
      O => memtest2_Mcompar_n0018_inst_cy_166
    );
  memtest2_Mcompar_n0018_inst_lut4_251 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest2_datain(8),
      ADR1 => memtest2_Mshreg_data4_9_60,
      ADR2 => memtest2_datain(9),
      ADR3 => memtest2_Mshreg_data4_8_61,
      O => memtest2_Mcompar_n0018_inst_lut4_25
    );
  memtest2_Mcompar_n0018_inst_lut4_261 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => memtest2_datain(10),
      ADR1 => memtest2_datain(11),
      ADR2 => memtest2_Mshreg_data4_11_58,
      ADR3 => memtest2_Mshreg_data4_10_59,
      O => memtest2_Mcompar_n0018_inst_lut4_26
    );
  memtest2_Mcompar_n0018_inst_cy_167_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0018_inst_cy_167_CYMUXG,
      O => memtest2_Mcompar_n0018_inst_cy_167
    );
  memtest2_Mcompar_n0018_inst_cy_167_514 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0018_inst_cy_167_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0018_inst_cy_166,
      SEL => memtest2_Mcompar_n0018_inst_lut4_26,
      O => memtest2_Mcompar_n0018_inst_cy_167_CYMUXG
    );
  memtest2_deq_1_LOGIC_ZERO_515 : X_ZERO
    port map (
      O => memtest2_deq_1_LOGIC_ZERO
    );
  memtest2_Mcompar_n0018_inst_cy_168_516 : X_MUX2
    port map (
      IA => memtest2_deq_1_LOGIC_ZERO,
      IB => memtest2_deq_1_CYINIT,
      SEL => memtest2_Mcompar_n0018_inst_lut4_27,
      O => memtest2_Mcompar_n0018_inst_cy_168
    );
  memtest2_Mcompar_n0018_inst_lut4_271 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => memtest2_Mshreg_data4_12_57,
      ADR1 => memtest2_datain(13),
      ADR2 => memtest2_datain(12),
      ADR3 => memtest2_Mshreg_data4_13_56,
      O => memtest2_Mcompar_n0018_inst_lut4_27
    );
  memtest2_Mcompar_n0018_inst_lut4_281 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => memtest2_Mshreg_data4_15_54,
      ADR1 => memtest2_Mshreg_data4_14_55,
      ADR2 => memtest2_datain(15),
      ADR3 => memtest2_datain(14),
      O => memtest2_Mcompar_n0018_inst_lut4_28
    );
  memtest2_deq_1_COUTUSED : X_BUF
    port map (
      I => memtest2_deq_1_CYMUXG,
      O => memtest2_deq(1)
    );
  memtest2_Mcompar_n0018_inst_cy_169 : X_MUX2
    port map (
      IA => memtest2_deq_1_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0018_inst_cy_168,
      SEL => memtest2_Mcompar_n0018_inst_lut4_28,
      O => memtest2_deq_1_CYMUXG
    );
  memtest2_deq_1_CYINIT_517 : X_BUF
    port map (
      I => memtest2_Mcompar_n0018_inst_cy_167,
      O => memtest2_deq_1_CYINIT
    );
  memtest2_Mcompar_n0027_inst_cy_153_LOGIC_ONE_518 : X_ONE
    port map (
      O => memtest2_Mcompar_n0027_inst_cy_153_LOGIC_ONE
    );
  memtest2_Mcompar_n0027_inst_cy_153_LOGIC_ZERO_519 : X_ZERO
    port map (
      O => memtest2_Mcompar_n0027_inst_cy_153_LOGIC_ZERO
    );
  memtest2_Mcompar_n0027_inst_cy_152_520 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0027_inst_cy_153_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0027_inst_cy_153_LOGIC_ONE,
      SEL => memtest2_SIG_2,
      O => memtest2_Mcompar_n0027_inst_cy_152
    );
  memtest2_BEL_2 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memtest2_cnt(1),
      ADR3 => VCC,
      O => memtest2_SIG_2
    );
  memtest2_BEL_3 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memtest2_cnt(1),
      ADR3 => VCC,
      O => memtest2_SIG_3
    );
  memtest2_Mcompar_n0027_inst_cy_153_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0027_inst_cy_153_CYMUXG,
      O => memtest2_Mcompar_n0027_inst_cy_153
    );
  memtest2_Mcompar_n0027_inst_cy_153_521 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0027_inst_cy_153_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0027_inst_cy_152,
      SEL => memtest2_SIG_3,
      O => memtest2_Mcompar_n0027_inst_cy_153_CYMUXG
    );
  memtest2_Mcompar_n0027_inst_cy_155_LOGIC_ONE_522 : X_ONE
    port map (
      O => memtest2_Mcompar_n0027_inst_cy_155_LOGIC_ONE
    );
  memtest2_Mcompar_n0027_inst_cy_154_523 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0027_inst_cy_155_LOGIC_ONE,
      IB => memtest2_Mcompar_n0027_inst_cy_155_CYINIT,
      SEL => memtest2_Mcompar_n0027_inst_lut4_19,
      O => memtest2_Mcompar_n0027_inst_cy_154
    );
  memtest2_Mcompar_n0027_inst_lut4_191 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(5),
      ADR1 => memtest2_cnt(4),
      ADR2 => memtest2_cnt(2),
      ADR3 => memtest2_cnt(3),
      O => memtest2_Mcompar_n0027_inst_lut4_19
    );
  memtest2_Mcompar_n0027_inst_lut4_201 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(8),
      ADR1 => memtest2_cnt(6),
      ADR2 => memtest2_cnt(7),
      ADR3 => memtest2_cnt(9),
      O => memtest2_Mcompar_n0027_inst_lut4_20
    );
  memtest2_Mcompar_n0027_inst_cy_155_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0027_inst_cy_155_CYMUXG,
      O => memtest2_Mcompar_n0027_inst_cy_155
    );
  memtest2_Mcompar_n0027_inst_cy_155_524 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0027_inst_cy_155_LOGIC_ONE,
      IB => memtest2_Mcompar_n0027_inst_cy_154,
      SEL => memtest2_Mcompar_n0027_inst_lut4_20,
      O => memtest2_Mcompar_n0027_inst_cy_155_CYMUXG
    );
  memtest2_Mcompar_n0027_inst_cy_155_CYINIT_525 : X_BUF
    port map (
      I => memtest2_Mcompar_n0027_inst_cy_153,
      O => memtest2_Mcompar_n0027_inst_cy_155_CYINIT
    );
  memtest2_Mcompar_n0027_inst_cy_157_LOGIC_ONE_526 : X_ONE
    port map (
      O => memtest2_Mcompar_n0027_inst_cy_157_LOGIC_ONE
    );
  memtest2_Mcompar_n0027_inst_cy_156_527 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0027_inst_cy_157_LOGIC_ONE,
      IB => memtest2_Mcompar_n0027_inst_cy_157_CYINIT,
      SEL => memtest2_Mcompar_n0027_inst_lut4_21,
      O => memtest2_Mcompar_n0027_inst_cy_156
    );
  memtest2_Mcompar_n0027_inst_lut4_211 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(12),
      ADR1 => memtest2_cnt(10),
      ADR2 => memtest2_cnt(13),
      ADR3 => memtest2_cnt(11),
      O => memtest2_Mcompar_n0027_inst_lut4_21
    );
  memtest2_Mcompar_n0027_inst_lut2_1241 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(15),
      ADR2 => memtest2_cnt(14),
      ADR3 => VCC,
      O => memtest2_Mcompar_n0027_inst_lut2_124
    );
  memtest2_Mcompar_n0027_inst_cy_157_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0027_inst_cy_157_CYMUXG,
      O => memtest2_Mcompar_n0027_inst_cy_157
    );
  memtest2_Mcompar_n0027_inst_cy_157_528 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0027_inst_cy_157_LOGIC_ONE,
      IB => memtest2_Mcompar_n0027_inst_cy_156,
      SEL => memtest2_Mcompar_n0027_inst_lut2_124,
      O => memtest2_Mcompar_n0027_inst_cy_157_CYMUXG
    );
  memtest2_Mcompar_n0027_inst_cy_157_CYINIT_529 : X_BUF
    port map (
      I => memtest2_Mcompar_n0027_inst_cy_155,
      O => memtest2_Mcompar_n0027_inst_cy_157_CYINIT
    );
  memtest2_n0027_LOGIC_ZERO_530 : X_ZERO
    port map (
      O => memtest2_n0027_LOGIC_ZERO
    );
  memtest2_Mcompar_n0027_inst_cy_158_531 : X_MUX2
    port map (
      IA => memtest2_n0027_LOGIC_ZERO,
      IB => memtest2_n0027_CYINIT,
      SEL => memtest2_SIG_4,
      O => memtest2_Mcompar_n0027_inst_cy_158
    );
  memtest2_BEL_4 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_SIG_4
    );
  memtest2_BEL_5 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_SIG_5
    );
  memtest2_n0027_COUTUSED : X_BUF
    port map (
      I => memtest2_n0027_CYMUXG,
      O => memtest2_n0027
    );
  memtest2_Mcompar_n0027_inst_cy_159 : X_MUX2
    port map (
      IA => memtest2_n0027_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0027_inst_cy_158,
      SEL => memtest2_SIG_5,
      O => memtest2_n0027_CYMUXG
    );
  memtest2_n0027_CYINIT_532 : X_BUF
    port map (
      I => memtest2_Mcompar_n0027_inst_cy_157,
      O => memtest2_n0027_CYINIT
    );
  memcontroller_addr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_5_OD,
      CE => MA_5_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_5_OFF_RST,
      O => memcontroller_ADDREXT(5)
    );
  MA_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_5_OFF_RST
    );
  memtest2_Mcompar_n0019_inst_cy_167_LOGIC_ONE_533 : X_ONE
    port map (
      O => memtest2_Mcompar_n0019_inst_cy_167_LOGIC_ONE
    );
  memtest2_Mcompar_n0019_inst_cy_167_LOGIC_ZERO_534 : X_ZERO
    port map (
      O => memtest2_Mcompar_n0019_inst_cy_167_LOGIC_ZERO
    );
  memtest2_Mcompar_n0019_inst_cy_166_535 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0019_inst_cy_167_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0019_inst_cy_167_LOGIC_ONE,
      SEL => memtest2_Mcompar_n0019_inst_lut4_25,
      O => memtest2_Mcompar_n0019_inst_cy_166
    );
  memtest2_Mcompar_n0019_inst_lut4_251 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => memtest2_Mshreg_data4_16_53,
      ADR1 => memtest2_Mshreg_data4_17_52,
      ADR2 => memtest2_datain(16),
      ADR3 => memtest2_datain(17),
      O => memtest2_Mcompar_n0019_inst_lut4_25
    );
  memtest2_Mcompar_n0019_inst_lut4_261 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => memtest2_Mshreg_data4_18_51,
      ADR1 => memtest2_Mshreg_data4_19_50,
      ADR2 => memtest2_datain(18),
      ADR3 => memtest2_datain(19),
      O => memtest2_Mcompar_n0019_inst_lut4_26
    );
  memtest2_Mcompar_n0019_inst_cy_167_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0019_inst_cy_167_CYMUXG,
      O => memtest2_Mcompar_n0019_inst_cy_167
    );
  memtest2_Mcompar_n0019_inst_cy_167_536 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0019_inst_cy_167_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0019_inst_cy_166,
      SEL => memtest2_Mcompar_n0019_inst_lut4_26,
      O => memtest2_Mcompar_n0019_inst_cy_167_CYMUXG
    );
  memtest2_deq_2_LOGIC_ZERO_537 : X_ZERO
    port map (
      O => memtest2_deq_2_LOGIC_ZERO
    );
  memtest2_Mcompar_n0019_inst_cy_168_538 : X_MUX2
    port map (
      IA => memtest2_deq_2_LOGIC_ZERO,
      IB => memtest2_deq_2_CYINIT,
      SEL => memtest2_Mcompar_n0019_inst_lut4_27,
      O => memtest2_Mcompar_n0019_inst_cy_168
    );
  memtest2_Mcompar_n0019_inst_lut4_271 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => memtest2_datain(20),
      ADR1 => memtest2_Mshreg_data4_21_48,
      ADR2 => memtest2_Mshreg_data4_20_49,
      ADR3 => memtest2_datain(21),
      O => memtest2_Mcompar_n0019_inst_lut4_27
    );
  memtest2_Mcompar_n0019_inst_lut4_281 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => memtest2_datain(22),
      ADR1 => memtest2_Mshreg_data4_22_47,
      ADR2 => memtest2_Mshreg_data4_23_46,
      ADR3 => memtest2_datain(23),
      O => memtest2_Mcompar_n0019_inst_lut4_28
    );
  memtest2_deq_2_COUTUSED : X_BUF
    port map (
      I => memtest2_deq_2_CYMUXG,
      O => memtest2_deq(2)
    );
  memtest2_Mcompar_n0019_inst_cy_169 : X_MUX2
    port map (
      IA => memtest2_deq_2_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0019_inst_cy_168,
      SEL => memtest2_Mcompar_n0019_inst_lut4_28,
      O => memtest2_deq_2_CYMUXG
    );
  memtest2_deq_2_CYINIT_539 : X_BUF
    port map (
      I => memtest2_Mcompar_n0019_inst_cy_167,
      O => memtest2_deq_2_CYINIT
    );
  txsim_counter_0_LOGIC_ZERO_540 : X_ZERO
    port map (
      O => txsim_counter_0_LOGIC_ZERO
    );
  txsim_counter_Madd_n0000_inst_cy_103_541 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_4,
      IB => txsim_counter_0_LOGIC_ZERO,
      SEL => txsim_counter_Madd_n0000_inst_lut2_103,
      O => txsim_counter_Madd_n0000_inst_cy_103
    );
  txsim_counter_Madd_n0000_inst_lut2_1031 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_4,
      ADR1 => txsim_counter(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => txsim_counter_Madd_n0000_inst_lut2_103
    );
  txsim_counter_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_58,
      ADR1 => VCC,
      ADR2 => txsim_counter(1),
      ADR3 => VCC,
      O => txsim_counter_0_GROM
    );
  txsim_counter_0_COUTUSED : X_BUF
    port map (
      I => txsim_counter_0_CYMUXG,
      O => txsim_counter_Madd_n0000_inst_cy_104
    );
  txsim_counter_Madd_n0000_inst_cy_104_542 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_58,
      IB => txsim_counter_Madd_n0000_inst_cy_103,
      SEL => txsim_counter_0_GROM,
      O => txsim_counter_0_CYMUXG
    );
  txsim_counter_Madd_n0000_inst_sum_104 : X_XOR2
    port map (
      I0 => txsim_counter_Madd_n0000_inst_cy_103,
      I1 => txsim_counter_0_GROM,
      O => txsim_counter_n0000(1)
    );
  txsim_counter_2_LOGIC_ZERO_543 : X_ZERO
    port map (
      O => txsim_counter_2_LOGIC_ZERO
    );
  txsim_counter_Madd_n0000_inst_cy_105_544 : X_MUX2
    port map (
      IA => txsim_counter_2_LOGIC_ZERO,
      IB => txsim_counter_2_CYINIT,
      SEL => txsim_counter_2_FROM,
      O => txsim_counter_Madd_n0000_inst_cy_105
    );
  txsim_counter_Madd_n0000_inst_sum_105 : X_XOR2
    port map (
      I0 => txsim_counter_2_CYINIT,
      I1 => txsim_counter_2_FROM,
      O => txsim_counter_n0000(2)
    );
  txsim_counter_2_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => txsim_counter(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => txsim_counter_2_FROM
    );
  txsim_counter_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => txsim_counter(3),
      ADR3 => VCC,
      O => txsim_counter_2_GROM
    );
  txsim_counter_2_COUTUSED : X_BUF
    port map (
      I => txsim_counter_2_CYMUXG,
      O => txsim_counter_Madd_n0000_inst_cy_106
    );
  txsim_counter_Madd_n0000_inst_cy_106_545 : X_MUX2
    port map (
      IA => txsim_counter_2_LOGIC_ZERO,
      IB => txsim_counter_Madd_n0000_inst_cy_105,
      SEL => txsim_counter_2_GROM,
      O => txsim_counter_2_CYMUXG
    );
  txsim_counter_Madd_n0000_inst_sum_106 : X_XOR2
    port map (
      I0 => txsim_counter_Madd_n0000_inst_cy_105,
      I1 => txsim_counter_2_GROM,
      O => txsim_counter_n0000(3)
    );
  txsim_counter_2_CYINIT_546 : X_BUF
    port map (
      I => txsim_counter_Madd_n0000_inst_cy_104,
      O => txsim_counter_2_CYINIT
    );
  txsim_counter_4_LOGIC_ZERO_547 : X_ZERO
    port map (
      O => txsim_counter_4_LOGIC_ZERO
    );
  txsim_counter_Madd_n0000_inst_cy_107_548 : X_MUX2
    port map (
      IA => txsim_counter_4_LOGIC_ZERO,
      IB => txsim_counter_4_CYINIT,
      SEL => txsim_counter_4_FROM,
      O => txsim_counter_Madd_n0000_inst_cy_107
    );
  txsim_counter_Madd_n0000_inst_sum_107 : X_XOR2
    port map (
      I0 => txsim_counter_4_CYINIT,
      I1 => txsim_counter_4_FROM,
      O => txsim_counter_n0000(4)
    );
  txsim_counter_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => txsim_counter(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => txsim_counter_4_FROM
    );
  txsim_counter_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => txsim_counter(5),
      ADR3 => VCC,
      O => txsim_counter_4_GROM
    );
  txsim_counter_4_COUTUSED : X_BUF
    port map (
      I => txsim_counter_4_CYMUXG,
      O => txsim_counter_Madd_n0000_inst_cy_108
    );
  txsim_counter_Madd_n0000_inst_cy_108_549 : X_MUX2
    port map (
      IA => txsim_counter_4_LOGIC_ZERO,
      IB => txsim_counter_Madd_n0000_inst_cy_107,
      SEL => txsim_counter_4_GROM,
      O => txsim_counter_4_CYMUXG
    );
  txsim_counter_Madd_n0000_inst_sum_108 : X_XOR2
    port map (
      I0 => txsim_counter_Madd_n0000_inst_cy_107,
      I1 => txsim_counter_4_GROM,
      O => txsim_counter_n0000(5)
    );
  txsim_counter_4_CYINIT_550 : X_BUF
    port map (
      I => txsim_counter_Madd_n0000_inst_cy_106,
      O => txsim_counter_4_CYINIT
    );
  txsim_counter_6_LOGIC_ZERO_551 : X_ZERO
    port map (
      O => txsim_counter_6_LOGIC_ZERO
    );
  txsim_counter_Madd_n0000_inst_cy_109_552 : X_MUX2
    port map (
      IA => txsim_counter_6_LOGIC_ZERO,
      IB => txsim_counter_6_CYINIT,
      SEL => txsim_counter_6_FROM,
      O => txsim_counter_Madd_n0000_inst_cy_109
    );
  txsim_counter_Madd_n0000_inst_sum_109 : X_XOR2
    port map (
      I0 => txsim_counter_6_CYINIT,
      I1 => txsim_counter_6_FROM,
      O => txsim_counter_n0000(6)
    );
  txsim_counter_6_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => txsim_counter(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => txsim_counter_6_FROM
    );
  txsim_counter_6_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => txsim_counter(7),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => txsim_counter_6_GROM
    );
  txsim_counter_6_COUTUSED : X_BUF
    port map (
      I => txsim_counter_6_CYMUXG,
      O => txsim_counter_Madd_n0000_inst_cy_110
    );
  txsim_counter_Madd_n0000_inst_cy_110_553 : X_MUX2
    port map (
      IA => txsim_counter_6_LOGIC_ZERO,
      IB => txsim_counter_Madd_n0000_inst_cy_109,
      SEL => txsim_counter_6_GROM,
      O => txsim_counter_6_CYMUXG
    );
  txsim_counter_Madd_n0000_inst_sum_110 : X_XOR2
    port map (
      I0 => txsim_counter_Madd_n0000_inst_cy_109,
      I1 => txsim_counter_6_GROM,
      O => txsim_counter_n0000(7)
    );
  txsim_counter_6_CYINIT_554 : X_BUF
    port map (
      I => txsim_counter_Madd_n0000_inst_cy_108,
      O => txsim_counter_6_CYINIT
    );
  txsim_counter_8_LOGIC_ZERO_555 : X_ZERO
    port map (
      O => txsim_counter_8_LOGIC_ZERO
    );
  txsim_counter_Madd_n0000_inst_cy_111_556 : X_MUX2
    port map (
      IA => txsim_counter_8_LOGIC_ZERO,
      IB => txsim_counter_8_CYINIT,
      SEL => txsim_counter_8_FROM,
      O => txsim_counter_Madd_n0000_inst_cy_111
    );
  txsim_counter_Madd_n0000_inst_sum_111 : X_XOR2
    port map (
      I0 => txsim_counter_8_CYINIT,
      I1 => txsim_counter_8_FROM,
      O => txsim_counter_n0000(8)
    );
  txsim_counter_8_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => txsim_counter(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => txsim_counter_8_FROM
    );
  txsim_counter_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => txsim_counter(9),
      ADR3 => VCC,
      O => txsim_counter_8_GROM
    );
  txsim_counter_8_COUTUSED : X_BUF
    port map (
      I => txsim_counter_8_CYMUXG,
      O => txsim_counter_Madd_n0000_inst_cy_112
    );
  txsim_counter_Madd_n0000_inst_cy_112_557 : X_MUX2
    port map (
      IA => txsim_counter_8_LOGIC_ZERO,
      IB => txsim_counter_Madd_n0000_inst_cy_111,
      SEL => txsim_counter_8_GROM,
      O => txsim_counter_8_CYMUXG
    );
  txsim_counter_Madd_n0000_inst_sum_112 : X_XOR2
    port map (
      I0 => txsim_counter_Madd_n0000_inst_cy_111,
      I1 => txsim_counter_8_GROM,
      O => txsim_counter_n0000(9)
    );
  txsim_counter_8_CYINIT_558 : X_BUF
    port map (
      I => txsim_counter_Madd_n0000_inst_cy_110,
      O => txsim_counter_8_CYINIT
    );
  txsim_counter_10_LOGIC_ZERO_559 : X_ZERO
    port map (
      O => txsim_counter_10_LOGIC_ZERO
    );
  txsim_counter_Madd_n0000_inst_cy_113_560 : X_MUX2
    port map (
      IA => txsim_counter_10_LOGIC_ZERO,
      IB => txsim_counter_10_CYINIT,
      SEL => txsim_counter_10_FROM,
      O => txsim_counter_Madd_n0000_inst_cy_113
    );
  txsim_counter_Madd_n0000_inst_sum_113 : X_XOR2
    port map (
      I0 => txsim_counter_10_CYINIT,
      I1 => txsim_counter_10_FROM,
      O => txsim_counter_n0000(10)
    );
  txsim_counter_10_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => txsim_counter(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => txsim_counter_10_FROM
    );
  txsim_counter_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => txsim_counter(11),
      ADR3 => VCC,
      O => txsim_counter_10_GROM
    );
  txsim_counter_10_COUTUSED : X_BUF
    port map (
      I => txsim_counter_10_CYMUXG,
      O => txsim_counter_Madd_n0000_inst_cy_114
    );
  txsim_counter_Madd_n0000_inst_cy_114_561 : X_MUX2
    port map (
      IA => txsim_counter_10_LOGIC_ZERO,
      IB => txsim_counter_Madd_n0000_inst_cy_113,
      SEL => txsim_counter_10_GROM,
      O => txsim_counter_10_CYMUXG
    );
  txsim_counter_Madd_n0000_inst_sum_114 : X_XOR2
    port map (
      I0 => txsim_counter_Madd_n0000_inst_cy_113,
      I1 => txsim_counter_10_GROM,
      O => txsim_counter_n0000(11)
    );
  txsim_counter_10_CYINIT_562 : X_BUF
    port map (
      I => txsim_counter_Madd_n0000_inst_cy_112,
      O => txsim_counter_10_CYINIT
    );
  txsim_counter_12_LOGIC_ZERO_563 : X_ZERO
    port map (
      O => txsim_counter_12_LOGIC_ZERO
    );
  txsim_counter_Madd_n0000_inst_cy_115_564 : X_MUX2
    port map (
      IA => txsim_counter_12_LOGIC_ZERO,
      IB => txsim_counter_12_CYINIT,
      SEL => txsim_counter_12_FROM,
      O => txsim_counter_Madd_n0000_inst_cy_115
    );
  txsim_counter_Madd_n0000_inst_sum_115 : X_XOR2
    port map (
      I0 => txsim_counter_12_CYINIT,
      I1 => txsim_counter_12_FROM,
      O => txsim_counter_n0000(12)
    );
  txsim_counter_12_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => txsim_counter(12),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => txsim_counter_12_FROM
    );
  txsim_counter_12_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => txsim_counter(13),
      ADR3 => VCC,
      O => txsim_counter_12_GROM
    );
  txsim_counter_12_COUTUSED : X_BUF
    port map (
      I => txsim_counter_12_CYMUXG,
      O => txsim_counter_Madd_n0000_inst_cy_116
    );
  txsim_counter_Madd_n0000_inst_cy_116_565 : X_MUX2
    port map (
      IA => txsim_counter_12_LOGIC_ZERO,
      IB => txsim_counter_Madd_n0000_inst_cy_115,
      SEL => txsim_counter_12_GROM,
      O => txsim_counter_12_CYMUXG
    );
  txsim_counter_Madd_n0000_inst_sum_116 : X_XOR2
    port map (
      I0 => txsim_counter_Madd_n0000_inst_cy_115,
      I1 => txsim_counter_12_GROM,
      O => txsim_counter_n0000(13)
    );
  txsim_counter_12_CYINIT_566 : X_BUF
    port map (
      I => txsim_counter_Madd_n0000_inst_cy_114,
      O => txsim_counter_12_CYINIT
    );
  txsim_counter_14_LOGIC_ZERO_567 : X_ZERO
    port map (
      O => txsim_counter_14_LOGIC_ZERO
    );
  txsim_counter_Madd_n0000_inst_cy_117_568 : X_MUX2
    port map (
      IA => txsim_counter_14_LOGIC_ZERO,
      IB => txsim_counter_14_CYINIT,
      SEL => txsim_counter_14_FROM,
      O => txsim_counter_Madd_n0000_inst_cy_117
    );
  txsim_counter_Madd_n0000_inst_sum_117 : X_XOR2
    port map (
      I0 => txsim_counter_14_CYINIT,
      I1 => txsim_counter_14_FROM,
      O => txsim_counter_n0000(14)
    );
  txsim_counter_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => txsim_counter(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => txsim_counter_14_FROM
    );
  txsim_counter_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => txsim_counter(15),
      ADR3 => VCC,
      O => txsim_counter_14_GROM
    );
  txsim_counter_14_COUTUSED : X_BUF
    port map (
      I => txsim_counter_14_CYMUXG,
      O => txsim_counter_Madd_n0000_inst_cy_118
    );
  txsim_counter_Madd_n0000_inst_cy_118_569 : X_MUX2
    port map (
      IA => txsim_counter_14_LOGIC_ZERO,
      IB => txsim_counter_Madd_n0000_inst_cy_117,
      SEL => txsim_counter_14_GROM,
      O => txsim_counter_14_CYMUXG
    );
  txsim_counter_Madd_n0000_inst_sum_118 : X_XOR2
    port map (
      I0 => txsim_counter_Madd_n0000_inst_cy_117,
      I1 => txsim_counter_14_GROM,
      O => txsim_counter_n0000(15)
    );
  txsim_counter_14_CYINIT_570 : X_BUF
    port map (
      I => txsim_counter_Madd_n0000_inst_cy_116,
      O => txsim_counter_14_CYINIT
    );
  txsim_counter_16_LOGIC_ZERO_571 : X_ZERO
    port map (
      O => txsim_counter_16_LOGIC_ZERO
    );
  txsim_counter_Madd_n0000_inst_cy_119_572 : X_MUX2
    port map (
      IA => txsim_counter_16_LOGIC_ZERO,
      IB => txsim_counter_16_CYINIT,
      SEL => txsim_counter_16_FROM,
      O => txsim_counter_Madd_n0000_inst_cy_119
    );
  txsim_counter_Madd_n0000_inst_sum_119 : X_XOR2
    port map (
      I0 => txsim_counter_16_CYINIT,
      I1 => txsim_counter_16_FROM,
      O => txsim_counter_n0000(16)
    );
  txsim_counter_16_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => txsim_counter(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => txsim_counter_16_FROM
    );
  txsim_counter_17_rt_573 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => txsim_counter(17),
      ADR3 => VCC,
      O => txsim_counter_17_rt
    );
  txsim_counter_Madd_n0000_inst_sum_120 : X_XOR2
    port map (
      I0 => txsim_counter_Madd_n0000_inst_cy_119,
      I1 => txsim_counter_17_rt,
      O => txsim_counter_n0000(17)
    );
  txsim_counter_16_CYINIT_574 : X_BUF
    port map (
      I => txsim_counter_Madd_n0000_inst_cy_118,
      O => txsim_counter_16_CYINIT
    );
  memtest2_Mcompar_n0028_inst_cy_145_LOGIC_ONE_575 : X_ONE
    port map (
      O => memtest2_Mcompar_n0028_inst_cy_145_LOGIC_ONE
    );
  memtest2_Mcompar_n0028_inst_cy_145_LOGIC_ZERO_576 : X_ZERO
    port map (
      O => memtest2_Mcompar_n0028_inst_cy_145_LOGIC_ZERO
    );
  memtest2_Mcompar_n0028_inst_cy_144_577 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0028_inst_cy_145_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0028_inst_cy_145_LOGIC_ONE,
      SEL => memtest2_Mcompar_n0028_inst_lut1_0,
      O => memtest2_Mcompar_n0028_inst_cy_144
    );
  memtest2_Mcompar_n0028_inst_lut1_01 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memtest2_cnt(0),
      ADR3 => VCC,
      O => memtest2_Mcompar_n0028_inst_lut1_0
    );
  memtest2_Mcompar_n0028_inst_lut1_11 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memtest2_cnt(0),
      ADR3 => VCC,
      O => memtest2_Mcompar_n0028_inst_lut1_1
    );
  memtest2_Mcompar_n0028_inst_cy_145_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0028_inst_cy_145_CYMUXG,
      O => memtest2_Mcompar_n0028_inst_cy_145
    );
  memtest2_Mcompar_n0028_inst_cy_145_578 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0028_inst_cy_145_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0028_inst_cy_144,
      SEL => memtest2_Mcompar_n0028_inst_lut1_1,
      O => memtest2_Mcompar_n0028_inst_cy_145_CYMUXG
    );
  memtest2_Mcompar_n0028_inst_cy_147_LOGIC_ONE_579 : X_ONE
    port map (
      O => memtest2_Mcompar_n0028_inst_cy_147_LOGIC_ONE
    );
  memtest2_Mcompar_n0028_inst_cy_146_580 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0028_inst_cy_147_LOGIC_ONE,
      IB => memtest2_Mcompar_n0028_inst_cy_147_CYINIT,
      SEL => memtest2_Mcompar_n0028_inst_lut2_121,
      O => memtest2_Mcompar_n0028_inst_cy_146
    );
  memtest2_Mcompar_n0028_inst_lut2_1211 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => memtest2_cnt(1),
      ADR1 => VCC,
      ADR2 => memtest2_cnt(2),
      ADR3 => VCC,
      O => memtest2_Mcompar_n0028_inst_lut2_121
    );
  memtest2_Mcompar_n0028_inst_lut2_1221 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => memtest2_cnt(1),
      ADR1 => memtest2_cnt(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_Mcompar_n0028_inst_lut2_122
    );
  memtest2_Mcompar_n0028_inst_cy_147_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0028_inst_cy_147_CYMUXG,
      O => memtest2_Mcompar_n0028_inst_cy_147
    );
  memtest2_Mcompar_n0028_inst_cy_147_581 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0028_inst_cy_147_LOGIC_ONE,
      IB => memtest2_Mcompar_n0028_inst_cy_146,
      SEL => memtest2_Mcompar_n0028_inst_lut2_122,
      O => memtest2_Mcompar_n0028_inst_cy_147_CYMUXG
    );
  memtest2_Mcompar_n0028_inst_cy_147_CYINIT_582 : X_BUF
    port map (
      I => memtest2_Mcompar_n0028_inst_cy_145,
      O => memtest2_Mcompar_n0028_inst_cy_147_CYINIT
    );
  memtest2_Mcompar_n0028_inst_lut4_16_LOGIC_ZERO_583 : X_ZERO
    port map (
      O => memtest2_Mcompar_n0028_inst_lut4_16_LOGIC_ZERO
    );
  memtest2_Mcompar_n0028_inst_cy_148_584 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0028_inst_lut4_16_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0028_inst_lut4_16_CYINIT,
      SEL => memtest2_Mcompar_n0028_inst_lut4_16_FROM,
      O => memtest2_Mcompar_n0028_inst_cy_148
    );
  memtest2_Mcompar_n0028_inst_lut4_161 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(4),
      ADR1 => memtest2_cnt(6),
      ADR2 => memtest2_cnt(5),
      ADR3 => memtest2_cnt(3),
      O => memtest2_Mcompar_n0028_inst_lut4_16_FROM
    );
  memtest2_Mcompar_n0028_inst_lut4_171 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(9),
      ADR1 => memtest2_cnt(7),
      ADR2 => memtest2_cnt(8),
      ADR3 => memtest2_cnt(10),
      O => memtest2_Mcompar_n0028_inst_lut4_17
    );
  memtest2_Mcompar_n0028_inst_lut4_16_COUTUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0028_inst_lut4_16_CYMUXG,
      O => memtest2_Mcompar_n0028_inst_cy_149
    );
  memtest2_Mcompar_n0028_inst_lut4_16_XUSED : X_BUF
    port map (
      I => memtest2_Mcompar_n0028_inst_lut4_16_FROM,
      O => memtest2_Mcompar_n0028_inst_lut4_16
    );
  memtest2_Mcompar_n0028_inst_cy_149_585 : X_MUX2
    port map (
      IA => memtest2_Mcompar_n0028_inst_lut4_16_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0028_inst_cy_148,
      SEL => memtest2_Mcompar_n0028_inst_lut4_17,
      O => memtest2_Mcompar_n0028_inst_lut4_16_CYMUXG
    );
  memtest2_Mcompar_n0028_inst_lut4_16_CYINIT_586 : X_BUF
    port map (
      I => memtest2_Mcompar_n0028_inst_cy_147,
      O => memtest2_Mcompar_n0028_inst_lut4_16_CYINIT
    );
  memtest2_n0028_LOGIC_ZERO_587 : X_ZERO
    port map (
      O => memtest2_n0028_LOGIC_ZERO
    );
  memtest2_Mcompar_n0028_inst_cy_150_588 : X_MUX2
    port map (
      IA => memtest2_n0028_LOGIC_ZERO,
      IB => memtest2_n0028_CYINIT,
      SEL => memtest2_Mcompar_n0028_inst_lut4_18,
      O => memtest2_Mcompar_n0028_inst_cy_150
    );
  memtest2_Mcompar_n0028_inst_lut4_181 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(12),
      ADR1 => memtest2_cnt(13),
      ADR2 => memtest2_cnt(11),
      ADR3 => memtest2_cnt(14),
      O => memtest2_Mcompar_n0028_inst_lut4_18
    );
  memtest2_Mcompar_n0028_inst_lut2_1231 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(16),
      ADR2 => memtest2_cnt(15),
      ADR3 => VCC,
      O => memtest2_Mcompar_n0028_inst_lut2_123
    );
  memtest2_n0028_COUTUSED : X_BUF
    port map (
      I => memtest2_n0028_CYMUXG,
      O => memtest2_n0028
    );
  memtest2_Mcompar_n0028_inst_cy_151 : X_MUX2
    port map (
      IA => memtest2_n0028_LOGIC_ZERO,
      IB => memtest2_Mcompar_n0028_inst_cy_150,
      SEL => memtest2_Mcompar_n0028_inst_lut2_123,
      O => memtest2_n0028_CYMUXG
    );
  memtest2_n0028_CYINIT_589 : X_BUF
    port map (
      I => memtest2_Mcompar_n0028_inst_cy_149,
      O => memtest2_n0028_CYINIT
    );
  d1_0_LOGIC_ZERO_590 : X_ZERO
    port map (
      O => d1_0_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_38_591 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_37,
      IB => d1_0_LOGIC_ZERO,
      SEL => memtest_datacnt_Madd_n0000_inst_lut2_38,
      O => memtest_datacnt_Madd_n0000_inst_cy_38
    );
  memtest_datacnt_Madd_n0000_inst_lut2_381 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_37,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(0),
      O => memtest_datacnt_Madd_n0000_inst_lut2_38
    );
  d1_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_26,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(1),
      O => d1_0_GROM
    );
  d1_0_COUTUSED : X_BUF
    port map (
      I => d1_0_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_39
    );
  memtest_datacnt_Madd_n0000_inst_cy_39_592 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_26,
      IB => memtest_datacnt_Madd_n0000_inst_cy_38,
      SEL => d1_0_GROM,
      O => d1_0_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_38,
      I1 => d1_0_GROM,
      O => memtest_datacnt_n0000(1)
    );
  d1_2_LOGIC_ZERO_593 : X_ZERO
    port map (
      O => d1_2_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_40_594 : X_MUX2
    port map (
      IA => d1_2_LOGIC_ZERO,
      IB => d1_2_CYINIT,
      SEL => d1_2_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_40
    );
  memtest_datacnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => d1_2_CYINIT,
      I1 => d1_2_FROM,
      O => memtest_datacnt_n0000(2)
    );
  d1_2_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(2),
      ADR3 => VCC,
      O => d1_2_FROM
    );
  d1_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(3),
      O => d1_2_GROM
    );
  d1_2_COUTUSED : X_BUF
    port map (
      I => d1_2_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_41
    );
  memtest_datacnt_Madd_n0000_inst_cy_41_595 : X_MUX2
    port map (
      IA => d1_2_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_40,
      SEL => d1_2_GROM,
      O => d1_2_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_40,
      I1 => d1_2_GROM,
      O => memtest_datacnt_n0000(3)
    );
  d1_2_CYINIT_596 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_39,
      O => d1_2_CYINIT
    );
  d1_4_LOGIC_ZERO_597 : X_ZERO
    port map (
      O => d1_4_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_42_598 : X_MUX2
    port map (
      IA => d1_4_LOGIC_ZERO,
      IB => d1_4_CYINIT,
      SEL => d1_4_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_42
    );
  memtest_datacnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => d1_4_CYINIT,
      I1 => d1_4_FROM,
      O => memtest_datacnt_n0000(4)
    );
  d1_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => d1_4_FROM
    );
  d1_4_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => d1_4_GROM
    );
  d1_4_COUTUSED : X_BUF
    port map (
      I => d1_4_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_43
    );
  memtest_datacnt_Madd_n0000_inst_cy_43_599 : X_MUX2
    port map (
      IA => d1_4_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_42,
      SEL => d1_4_GROM,
      O => d1_4_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_42,
      I1 => d1_4_GROM,
      O => memtest_datacnt_n0000(5)
    );
  d1_4_CYINIT_600 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_41,
      O => d1_4_CYINIT
    );
  d1_6_LOGIC_ZERO_601 : X_ZERO
    port map (
      O => d1_6_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_44_602 : X_MUX2
    port map (
      IA => d1_6_LOGIC_ZERO,
      IB => d1_6_CYINIT,
      SEL => d1_6_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_44
    );
  memtest_datacnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => d1_6_CYINIT,
      I1 => d1_6_FROM,
      O => memtest_datacnt_n0000(6)
    );
  d1_6_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(6),
      ADR3 => VCC,
      O => d1_6_FROM
    );
  d1_6_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(7),
      ADR3 => VCC,
      O => d1_6_GROM
    );
  d1_6_COUTUSED : X_BUF
    port map (
      I => d1_6_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_45
    );
  memtest_datacnt_Madd_n0000_inst_cy_45_603 : X_MUX2
    port map (
      IA => d1_6_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_44,
      SEL => d1_6_GROM,
      O => d1_6_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_44,
      I1 => d1_6_GROM,
      O => memtest_datacnt_n0000(7)
    );
  d1_6_CYINIT_604 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_43,
      O => d1_6_CYINIT
    );
  memcontroller_addr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_6_OD,
      CE => MA_6_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_6_OFF_RST,
      O => memcontroller_ADDREXT(6)
    );
  MA_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_6_OFF_RST
    );
  d1_8_LOGIC_ZERO_605 : X_ZERO
    port map (
      O => d1_8_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_46_606 : X_MUX2
    port map (
      IA => d1_8_LOGIC_ZERO,
      IB => d1_8_CYINIT,
      SEL => d1_8_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_46
    );
  memtest_datacnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => d1_8_CYINIT,
      I1 => d1_8_FROM,
      O => memtest_datacnt_n0000(8)
    );
  d1_8_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(8),
      O => d1_8_FROM
    );
  d1_8_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(9),
      O => d1_8_GROM
    );
  d1_8_COUTUSED : X_BUF
    port map (
      I => d1_8_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_47
    );
  memtest_datacnt_Madd_n0000_inst_cy_47_607 : X_MUX2
    port map (
      IA => d1_8_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_46,
      SEL => d1_8_GROM,
      O => d1_8_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_46,
      I1 => d1_8_GROM,
      O => memtest_datacnt_n0000(9)
    );
  d1_8_CYINIT_608 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_45,
      O => d1_8_CYINIT
    );
  d1_10_LOGIC_ZERO_609 : X_ZERO
    port map (
      O => d1_10_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_48_610 : X_MUX2
    port map (
      IA => d1_10_LOGIC_ZERO,
      IB => d1_10_CYINIT,
      SEL => d1_10_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_48
    );
  memtest_datacnt_Madd_n0000_inst_sum_48 : X_XOR2
    port map (
      I0 => d1_10_CYINIT,
      I1 => d1_10_FROM,
      O => memtest_datacnt_n0000(10)
    );
  d1_10_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(10),
      O => d1_10_FROM
    );
  d1_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(11),
      ADR3 => VCC,
      O => d1_10_GROM
    );
  d1_10_COUTUSED : X_BUF
    port map (
      I => d1_10_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_49
    );
  memtest_datacnt_Madd_n0000_inst_cy_49_611 : X_MUX2
    port map (
      IA => d1_10_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_48,
      SEL => d1_10_GROM,
      O => d1_10_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_49 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_48,
      I1 => d1_10_GROM,
      O => memtest_datacnt_n0000(11)
    );
  d1_10_CYINIT_612 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_47,
      O => d1_10_CYINIT
    );
  d1_12_LOGIC_ZERO_613 : X_ZERO
    port map (
      O => d1_12_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_50_614 : X_MUX2
    port map (
      IA => d1_12_LOGIC_ZERO,
      IB => d1_12_CYINIT,
      SEL => d1_12_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_50
    );
  memtest_datacnt_Madd_n0000_inst_sum_50 : X_XOR2
    port map (
      I0 => d1_12_CYINIT,
      I1 => d1_12_FROM,
      O => memtest_datacnt_n0000(12)
    );
  d1_12_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(12),
      ADR3 => VCC,
      O => d1_12_FROM
    );
  d1_12_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(13),
      ADR3 => VCC,
      O => d1_12_GROM
    );
  d1_12_COUTUSED : X_BUF
    port map (
      I => d1_12_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_51
    );
  memtest_datacnt_Madd_n0000_inst_cy_51_615 : X_MUX2
    port map (
      IA => d1_12_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_50,
      SEL => d1_12_GROM,
      O => d1_12_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_51 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_50,
      I1 => d1_12_GROM,
      O => memtest_datacnt_n0000(13)
    );
  d1_12_CYINIT_616 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_49,
      O => d1_12_CYINIT
    );
  d1_14_LOGIC_ZERO_617 : X_ZERO
    port map (
      O => d1_14_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_52_618 : X_MUX2
    port map (
      IA => d1_14_LOGIC_ZERO,
      IB => d1_14_CYINIT,
      SEL => d1_14_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_52
    );
  memtest_datacnt_Madd_n0000_inst_sum_52 : X_XOR2
    port map (
      I0 => d1_14_CYINIT,
      I1 => d1_14_FROM,
      O => memtest_datacnt_n0000(14)
    );
  d1_14_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(14),
      O => d1_14_FROM
    );
  d1_14_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(15),
      ADR2 => VCC,
      ADR3 => VCC,
      O => d1_14_GROM
    );
  d1_14_COUTUSED : X_BUF
    port map (
      I => d1_14_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_53
    );
  memtest_datacnt_Madd_n0000_inst_cy_53_619 : X_MUX2
    port map (
      IA => d1_14_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_52,
      SEL => d1_14_GROM,
      O => d1_14_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_53 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_52,
      I1 => d1_14_GROM,
      O => memtest_datacnt_n0000(15)
    );
  d1_14_CYINIT_620 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_51,
      O => d1_14_CYINIT
    );
  d1_16_LOGIC_ZERO_621 : X_ZERO
    port map (
      O => d1_16_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_54_622 : X_MUX2
    port map (
      IA => d1_16_LOGIC_ZERO,
      IB => d1_16_CYINIT,
      SEL => d1_16_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_54
    );
  memtest_datacnt_Madd_n0000_inst_sum_54 : X_XOR2
    port map (
      I0 => d1_16_CYINIT,
      I1 => d1_16_FROM,
      O => memtest_datacnt_n0000(16)
    );
  d1_16_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(16),
      O => d1_16_FROM
    );
  d1_16_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(17),
      O => d1_16_GROM
    );
  d1_16_COUTUSED : X_BUF
    port map (
      I => d1_16_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_55
    );
  memtest_datacnt_Madd_n0000_inst_cy_55_623 : X_MUX2
    port map (
      IA => d1_16_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_54,
      SEL => d1_16_GROM,
      O => d1_16_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_55 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_54,
      I1 => d1_16_GROM,
      O => memtest_datacnt_n0000(17)
    );
  d1_16_CYINIT_624 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_53,
      O => d1_16_CYINIT
    );
  d1_18_LOGIC_ZERO_625 : X_ZERO
    port map (
      O => d1_18_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_56_626 : X_MUX2
    port map (
      IA => d1_18_LOGIC_ZERO,
      IB => d1_18_CYINIT,
      SEL => d1_18_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_56
    );
  memtest_datacnt_Madd_n0000_inst_sum_56 : X_XOR2
    port map (
      I0 => d1_18_CYINIT,
      I1 => d1_18_FROM,
      O => memtest_datacnt_n0000(18)
    );
  d1_18_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(18),
      ADR3 => VCC,
      O => d1_18_FROM
    );
  d1_18_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(19),
      ADR2 => VCC,
      ADR3 => VCC,
      O => d1_18_GROM
    );
  d1_18_COUTUSED : X_BUF
    port map (
      I => d1_18_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_57
    );
  memtest_datacnt_Madd_n0000_inst_cy_57_627 : X_MUX2
    port map (
      IA => d1_18_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_56,
      SEL => d1_18_GROM,
      O => d1_18_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_57 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_56,
      I1 => d1_18_GROM,
      O => memtest_datacnt_n0000(19)
    );
  d1_18_CYINIT_628 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_55,
      O => d1_18_CYINIT
    );
  d1_20_LOGIC_ZERO_629 : X_ZERO
    port map (
      O => d1_20_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_58_630 : X_MUX2
    port map (
      IA => d1_20_LOGIC_ZERO,
      IB => d1_20_CYINIT,
      SEL => d1_20_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_58
    );
  memtest_datacnt_Madd_n0000_inst_sum_58 : X_XOR2
    port map (
      I0 => d1_20_CYINIT,
      I1 => d1_20_FROM,
      O => memtest_datacnt_n0000(20)
    );
  d1_20_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(20),
      ADR3 => VCC,
      O => d1_20_FROM
    );
  d1_20_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(21),
      O => d1_20_GROM
    );
  d1_20_COUTUSED : X_BUF
    port map (
      I => d1_20_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_59
    );
  memtest_datacnt_Madd_n0000_inst_cy_59_631 : X_MUX2
    port map (
      IA => d1_20_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_58,
      SEL => d1_20_GROM,
      O => d1_20_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_59 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_58,
      I1 => d1_20_GROM,
      O => memtest_datacnt_n0000(21)
    );
  d1_20_CYINIT_632 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_57,
      O => d1_20_CYINIT
    );
  d1_22_LOGIC_ZERO_633 : X_ZERO
    port map (
      O => d1_22_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_60_634 : X_MUX2
    port map (
      IA => d1_22_LOGIC_ZERO,
      IB => d1_22_CYINIT,
      SEL => d1_22_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_60
    );
  memtest_datacnt_Madd_n0000_inst_sum_60 : X_XOR2
    port map (
      I0 => d1_22_CYINIT,
      I1 => d1_22_FROM,
      O => memtest_datacnt_n0000(22)
    );
  d1_22_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(22),
      O => d1_22_FROM
    );
  d1_22_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(23),
      ADR3 => VCC,
      O => d1_22_GROM
    );
  d1_22_COUTUSED : X_BUF
    port map (
      I => d1_22_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_61
    );
  memtest_datacnt_Madd_n0000_inst_cy_61_635 : X_MUX2
    port map (
      IA => d1_22_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_60,
      SEL => d1_22_GROM,
      O => d1_22_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_61 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_60,
      I1 => d1_22_GROM,
      O => memtest_datacnt_n0000(23)
    );
  d1_22_CYINIT_636 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_59,
      O => d1_22_CYINIT
    );
  d1_24_LOGIC_ZERO_637 : X_ZERO
    port map (
      O => d1_24_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_62_638 : X_MUX2
    port map (
      IA => d1_24_LOGIC_ZERO,
      IB => d1_24_CYINIT,
      SEL => d1_24_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_62
    );
  memtest_datacnt_Madd_n0000_inst_sum_62 : X_XOR2
    port map (
      I0 => d1_24_CYINIT,
      I1 => d1_24_FROM,
      O => memtest_datacnt_n0000(24)
    );
  d1_24_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(24),
      ADR3 => VCC,
      O => d1_24_FROM
    );
  d1_24_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(25),
      ADR3 => VCC,
      O => d1_24_GROM
    );
  d1_24_COUTUSED : X_BUF
    port map (
      I => d1_24_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_63
    );
  memtest_datacnt_Madd_n0000_inst_cy_63_639 : X_MUX2
    port map (
      IA => d1_24_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_62,
      SEL => d1_24_GROM,
      O => d1_24_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_63 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_62,
      I1 => d1_24_GROM,
      O => memtest_datacnt_n0000(25)
    );
  d1_24_CYINIT_640 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_61,
      O => d1_24_CYINIT
    );
  d1_26_LOGIC_ZERO_641 : X_ZERO
    port map (
      O => d1_26_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_64_642 : X_MUX2
    port map (
      IA => d1_26_LOGIC_ZERO,
      IB => d1_26_CYINIT,
      SEL => d1_26_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_64
    );
  memtest_datacnt_Madd_n0000_inst_sum_64 : X_XOR2
    port map (
      I0 => d1_26_CYINIT,
      I1 => d1_26_FROM,
      O => memtest_datacnt_n0000(26)
    );
  d1_26_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(26),
      O => d1_26_FROM
    );
  d1_26_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(27),
      ADR3 => VCC,
      O => d1_26_GROM
    );
  d1_26_COUTUSED : X_BUF
    port map (
      I => d1_26_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_65
    );
  memtest_datacnt_Madd_n0000_inst_cy_65_643 : X_MUX2
    port map (
      IA => d1_26_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_64,
      SEL => d1_26_GROM,
      O => d1_26_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_65 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_64,
      I1 => d1_26_GROM,
      O => memtest_datacnt_n0000(27)
    );
  d1_26_CYINIT_644 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_63,
      O => d1_26_CYINIT
    );
  d1_28_LOGIC_ZERO_645 : X_ZERO
    port map (
      O => d1_28_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_66_646 : X_MUX2
    port map (
      IA => d1_28_LOGIC_ZERO,
      IB => d1_28_CYINIT,
      SEL => d1_28_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_66
    );
  memtest_datacnt_Madd_n0000_inst_sum_66 : X_XOR2
    port map (
      I0 => d1_28_CYINIT,
      I1 => d1_28_FROM,
      O => memtest_datacnt_n0000(28)
    );
  d1_28_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(28),
      O => d1_28_FROM
    );
  d1_28_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(29),
      O => d1_28_GROM
    );
  d1_28_COUTUSED : X_BUF
    port map (
      I => d1_28_CYMUXG,
      O => memtest_datacnt_Madd_n0000_inst_cy_67
    );
  memtest_datacnt_Madd_n0000_inst_cy_67_647 : X_MUX2
    port map (
      IA => d1_28_LOGIC_ZERO,
      IB => memtest_datacnt_Madd_n0000_inst_cy_66,
      SEL => d1_28_GROM,
      O => d1_28_CYMUXG
    );
  memtest_datacnt_Madd_n0000_inst_sum_67 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_66,
      I1 => d1_28_GROM,
      O => memtest_datacnt_n0000(29)
    );
  d1_28_CYINIT_648 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_65,
      O => d1_28_CYINIT
    );
  d1_30_LOGIC_ZERO_649 : X_ZERO
    port map (
      O => d1_30_LOGIC_ZERO
    );
  memtest_datacnt_Madd_n0000_inst_cy_68_650 : X_MUX2
    port map (
      IA => d1_30_LOGIC_ZERO,
      IB => d1_30_CYINIT,
      SEL => d1_30_FROM,
      O => memtest_datacnt_Madd_n0000_inst_cy_68
    );
  memtest_datacnt_Madd_n0000_inst_sum_68 : X_XOR2
    port map (
      I0 => d1_30_CYINIT,
      I1 => d1_30_FROM,
      O => memtest_datacnt_n0000(30)
    );
  d1_30_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(30),
      O => d1_30_FROM
    );
  d1_31_rt_651 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(31),
      ADR3 => VCC,
      O => d1_31_rt
    );
  memtest_datacnt_Madd_n0000_inst_sum_69 : X_XOR2
    port map (
      I0 => memtest_datacnt_Madd_n0000_inst_cy_68,
      I1 => d1_31_rt,
      O => memtest_datacnt_n0000(31)
    );
  d1_30_CYINIT_652 : X_BUF
    port map (
      I => memtest_datacnt_Madd_n0000_inst_cy_67,
      O => d1_30_CYINIT
    );
  addr1_0_LOGIC_ZERO_653 : X_ZERO
    port map (
      O => addr1_0_LOGIC_ZERO
    );
  memtest_addrcnt_Madd_n0000_inst_cy_70_654 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_22,
      IB => addr1_0_LOGIC_ZERO,
      SEL => memtest_addrcnt_Madd_n0000_inst_lut2_70,
      O => memtest_addrcnt_Madd_n0000_inst_cy_70
    );
  memtest_addrcnt_Madd_n0000_inst_lut2_701 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_22,
      ADR1 => addr1(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest_addrcnt_Madd_n0000_inst_lut2_70
    );
  addr1_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_8,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr1(1),
      O => addr1_0_GROM
    );
  addr1_0_COUTUSED : X_BUF
    port map (
      I => addr1_0_CYMUXG,
      O => memtest_addrcnt_Madd_n0000_inst_cy_71
    );
  memtest_addrcnt_Madd_n0000_inst_cy_71_655 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_8,
      IB => memtest_addrcnt_Madd_n0000_inst_cy_70,
      SEL => addr1_0_GROM,
      O => addr1_0_CYMUXG
    );
  memtest_addrcnt_Madd_n0000_inst_sum_71 : X_XOR2
    port map (
      I0 => memtest_addrcnt_Madd_n0000_inst_cy_70,
      I1 => addr1_0_GROM,
      O => memtest_addrcnt_n0000(1)
    );
  addr1_2_LOGIC_ZERO_656 : X_ZERO
    port map (
      O => addr1_2_LOGIC_ZERO
    );
  memtest_addrcnt_Madd_n0000_inst_cy_72_657 : X_MUX2
    port map (
      IA => addr1_2_LOGIC_ZERO,
      IB => addr1_2_CYINIT,
      SEL => addr1_2_FROM,
      O => memtest_addrcnt_Madd_n0000_inst_cy_72
    );
  memtest_addrcnt_Madd_n0000_inst_sum_72 : X_XOR2
    port map (
      I0 => addr1_2_CYINIT,
      I1 => addr1_2_FROM,
      O => memtest_addrcnt_n0000(2)
    );
  addr1_2_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => addr1(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr1_2_FROM
    );
  addr1_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr1(3),
      ADR3 => VCC,
      O => addr1_2_GROM
    );
  addr1_2_COUTUSED : X_BUF
    port map (
      I => addr1_2_CYMUXG,
      O => memtest_addrcnt_Madd_n0000_inst_cy_73
    );
  memtest_addrcnt_Madd_n0000_inst_cy_73_658 : X_MUX2
    port map (
      IA => addr1_2_LOGIC_ZERO,
      IB => memtest_addrcnt_Madd_n0000_inst_cy_72,
      SEL => addr1_2_GROM,
      O => addr1_2_CYMUXG
    );
  memtest_addrcnt_Madd_n0000_inst_sum_73 : X_XOR2
    port map (
      I0 => memtest_addrcnt_Madd_n0000_inst_cy_72,
      I1 => addr1_2_GROM,
      O => memtest_addrcnt_n0000(3)
    );
  addr1_2_CYINIT_659 : X_BUF
    port map (
      I => memtest_addrcnt_Madd_n0000_inst_cy_71,
      O => addr1_2_CYINIT
    );
  addr1_4_LOGIC_ZERO_660 : X_ZERO
    port map (
      O => addr1_4_LOGIC_ZERO
    );
  memtest_addrcnt_Madd_n0000_inst_cy_74_661 : X_MUX2
    port map (
      IA => addr1_4_LOGIC_ZERO,
      IB => addr1_4_CYINIT,
      SEL => addr1_4_FROM,
      O => memtest_addrcnt_Madd_n0000_inst_cy_74
    );
  memtest_addrcnt_Madd_n0000_inst_sum_74 : X_XOR2
    port map (
      I0 => addr1_4_CYINIT,
      I1 => addr1_4_FROM,
      O => memtest_addrcnt_n0000(4)
    );
  addr1_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr1(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr1_4_FROM
    );
  addr1_4_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => addr1(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr1_4_GROM
    );
  addr1_4_COUTUSED : X_BUF
    port map (
      I => addr1_4_CYMUXG,
      O => memtest_addrcnt_Madd_n0000_inst_cy_75
    );
  memtest_addrcnt_Madd_n0000_inst_cy_75_662 : X_MUX2
    port map (
      IA => addr1_4_LOGIC_ZERO,
      IB => memtest_addrcnt_Madd_n0000_inst_cy_74,
      SEL => addr1_4_GROM,
      O => addr1_4_CYMUXG
    );
  memtest_addrcnt_Madd_n0000_inst_sum_75 : X_XOR2
    port map (
      I0 => memtest_addrcnt_Madd_n0000_inst_cy_74,
      I1 => addr1_4_GROM,
      O => memtest_addrcnt_n0000(5)
    );
  addr1_4_CYINIT_663 : X_BUF
    port map (
      I => memtest_addrcnt_Madd_n0000_inst_cy_73,
      O => addr1_4_CYINIT
    );
  addr1_6_LOGIC_ZERO_664 : X_ZERO
    port map (
      O => addr1_6_LOGIC_ZERO
    );
  memtest_addrcnt_Madd_n0000_inst_cy_76_665 : X_MUX2
    port map (
      IA => addr1_6_LOGIC_ZERO,
      IB => addr1_6_CYINIT,
      SEL => addr1_6_FROM,
      O => memtest_addrcnt_Madd_n0000_inst_cy_76
    );
  memtest_addrcnt_Madd_n0000_inst_sum_76 : X_XOR2
    port map (
      I0 => addr1_6_CYINIT,
      I1 => addr1_6_FROM,
      O => memtest_addrcnt_n0000(6)
    );
  addr1_6_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr1(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr1_6_FROM
    );
  addr1_6_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr1(7),
      O => addr1_6_GROM
    );
  addr1_6_COUTUSED : X_BUF
    port map (
      I => addr1_6_CYMUXG,
      O => memtest_addrcnt_Madd_n0000_inst_cy_77
    );
  memtest_addrcnt_Madd_n0000_inst_cy_77_666 : X_MUX2
    port map (
      IA => addr1_6_LOGIC_ZERO,
      IB => memtest_addrcnt_Madd_n0000_inst_cy_76,
      SEL => addr1_6_GROM,
      O => addr1_6_CYMUXG
    );
  memtest_addrcnt_Madd_n0000_inst_sum_77 : X_XOR2
    port map (
      I0 => memtest_addrcnt_Madd_n0000_inst_cy_76,
      I1 => addr1_6_GROM,
      O => memtest_addrcnt_n0000(7)
    );
  addr1_6_CYINIT_667 : X_BUF
    port map (
      I => memtest_addrcnt_Madd_n0000_inst_cy_75,
      O => addr1_6_CYINIT
    );
  addr1_8_LOGIC_ZERO_668 : X_ZERO
    port map (
      O => addr1_8_LOGIC_ZERO
    );
  memtest_addrcnt_Madd_n0000_inst_cy_78_669 : X_MUX2
    port map (
      IA => addr1_8_LOGIC_ZERO,
      IB => addr1_8_CYINIT,
      SEL => addr1_8_FROM,
      O => memtest_addrcnt_Madd_n0000_inst_cy_78
    );
  memtest_addrcnt_Madd_n0000_inst_sum_78 : X_XOR2
    port map (
      I0 => addr1_8_CYINIT,
      I1 => addr1_8_FROM,
      O => memtest_addrcnt_n0000(8)
    );
  addr1_8_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => addr1(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr1_8_FROM
    );
  addr1_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr1(9),
      ADR3 => VCC,
      O => addr1_8_GROM
    );
  addr1_8_COUTUSED : X_BUF
    port map (
      I => addr1_8_CYMUXG,
      O => memtest_addrcnt_Madd_n0000_inst_cy_79
    );
  memtest_addrcnt_Madd_n0000_inst_cy_79_670 : X_MUX2
    port map (
      IA => addr1_8_LOGIC_ZERO,
      IB => memtest_addrcnt_Madd_n0000_inst_cy_78,
      SEL => addr1_8_GROM,
      O => addr1_8_CYMUXG
    );
  memtest_addrcnt_Madd_n0000_inst_sum_79 : X_XOR2
    port map (
      I0 => memtest_addrcnt_Madd_n0000_inst_cy_78,
      I1 => addr1_8_GROM,
      O => memtest_addrcnt_n0000(9)
    );
  addr1_8_CYINIT_671 : X_BUF
    port map (
      I => memtest_addrcnt_Madd_n0000_inst_cy_77,
      O => addr1_8_CYINIT
    );
  addr1_10_LOGIC_ZERO_672 : X_ZERO
    port map (
      O => addr1_10_LOGIC_ZERO
    );
  memtest_addrcnt_Madd_n0000_inst_cy_80_673 : X_MUX2
    port map (
      IA => addr1_10_LOGIC_ZERO,
      IB => addr1_10_CYINIT,
      SEL => addr1_10_FROM,
      O => memtest_addrcnt_Madd_n0000_inst_cy_80
    );
  memtest_addrcnt_Madd_n0000_inst_sum_80 : X_XOR2
    port map (
      I0 => addr1_10_CYINIT,
      I1 => addr1_10_FROM,
      O => memtest_addrcnt_n0000(10)
    );
  addr1_10_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => addr1(10),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr1_10_FROM
    );
  addr1_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr1(11),
      O => addr1_10_GROM
    );
  addr1_10_COUTUSED : X_BUF
    port map (
      I => addr1_10_CYMUXG,
      O => memtest_addrcnt_Madd_n0000_inst_cy_81
    );
  memtest_addrcnt_Madd_n0000_inst_cy_81_674 : X_MUX2
    port map (
      IA => addr1_10_LOGIC_ZERO,
      IB => memtest_addrcnt_Madd_n0000_inst_cy_80,
      SEL => addr1_10_GROM,
      O => addr1_10_CYMUXG
    );
  memtest_addrcnt_Madd_n0000_inst_sum_81 : X_XOR2
    port map (
      I0 => memtest_addrcnt_Madd_n0000_inst_cy_80,
      I1 => addr1_10_GROM,
      O => memtest_addrcnt_n0000(11)
    );
  addr1_10_CYINIT_675 : X_BUF
    port map (
      I => memtest_addrcnt_Madd_n0000_inst_cy_79,
      O => addr1_10_CYINIT
    );
  addr1_12_LOGIC_ZERO_676 : X_ZERO
    port map (
      O => addr1_12_LOGIC_ZERO
    );
  memtest_addrcnt_Madd_n0000_inst_cy_82_677 : X_MUX2
    port map (
      IA => addr1_12_LOGIC_ZERO,
      IB => addr1_12_CYINIT,
      SEL => addr1_12_FROM,
      O => memtest_addrcnt_Madd_n0000_inst_cy_82
    );
  memtest_addrcnt_Madd_n0000_inst_sum_82 : X_XOR2
    port map (
      I0 => addr1_12_CYINIT,
      I1 => addr1_12_FROM,
      O => memtest_addrcnt_n0000(12)
    );
  addr1_12_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => addr1(12),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr1_12_FROM
    );
  addr1_12_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr1(13),
      O => addr1_12_GROM
    );
  addr1_12_COUTUSED : X_BUF
    port map (
      I => addr1_12_CYMUXG,
      O => memtest_addrcnt_Madd_n0000_inst_cy_83
    );
  memtest_addrcnt_Madd_n0000_inst_cy_83_678 : X_MUX2
    port map (
      IA => addr1_12_LOGIC_ZERO,
      IB => memtest_addrcnt_Madd_n0000_inst_cy_82,
      SEL => addr1_12_GROM,
      O => addr1_12_CYMUXG
    );
  memtest_addrcnt_Madd_n0000_inst_sum_83 : X_XOR2
    port map (
      I0 => memtest_addrcnt_Madd_n0000_inst_cy_82,
      I1 => addr1_12_GROM,
      O => memtest_addrcnt_n0000(13)
    );
  addr1_12_CYINIT_679 : X_BUF
    port map (
      I => memtest_addrcnt_Madd_n0000_inst_cy_81,
      O => addr1_12_CYINIT
    );
  memcontroller_addr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_7_OD,
      CE => MA_7_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_7_OFF_RST,
      O => memcontroller_ADDREXT(7)
    );
  MA_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_7_OFF_RST
    );
  addr1_14_LOGIC_ZERO_680 : X_ZERO
    port map (
      O => addr1_14_LOGIC_ZERO
    );
  memtest_addrcnt_Madd_n0000_inst_cy_84_681 : X_MUX2
    port map (
      IA => addr1_14_LOGIC_ZERO,
      IB => addr1_14_CYINIT,
      SEL => addr1_14_FROM,
      O => memtest_addrcnt_Madd_n0000_inst_cy_84
    );
  memtest_addrcnt_Madd_n0000_inst_sum_84 : X_XOR2
    port map (
      I0 => addr1_14_CYINIT,
      I1 => addr1_14_FROM,
      O => memtest_addrcnt_n0000(14)
    );
  addr1_14_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => addr1(14),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr1_14_FROM
    );
  addr1_15_rt_682 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr1(15),
      ADR3 => VCC,
      O => addr1_15_rt
    );
  memtest_addrcnt_Madd_n0000_inst_sum_85 : X_XOR2
    port map (
      I0 => memtest_addrcnt_Madd_n0000_inst_cy_84,
      I1 => addr1_15_rt,
      O => memtest_addrcnt_n0000(15)
    );
  addr1_14_CYINIT_683 : X_BUF
    port map (
      I => memtest_addrcnt_Madd_n0000_inst_cy_83,
      O => addr1_14_CYINIT
    );
  memcontroller_Ker256691 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => memcontroller_clknum(0),
      O => addr2_13_FROM
    );
  memtest2_n00511_1_684 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memtest2_cs(0),
      ADR3 => memcontroller_Ker256691_O,
      O => addr2_13_GROM
    );
  addr2_13_XUSED : X_BUF
    port map (
      I => addr2_13_FROM,
      O => memcontroller_Ker256691_O
    );
  addr2_13_YUSED : X_BUF
    port map (
      I => addr2_13_GROM,
      O => memtest2_n00511_1
    );
  memtest2_datain_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_11_FFY_RST
    );
  memtest2_datain_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(10),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_11_FFY_RST,
      O => memtest2_datain(10)
    );
  memtest2_n00511 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cs(0),
      ADR2 => memcontroller_Ker256691_O,
      ADR3 => VCC,
      O => memtest2_datain_11_GROM
    );
  memtest2_datain_11_YUSED : X_BUF
    port map (
      I => memtest2_datain_11_GROM,
      O => memtest2_n00511_O
    );
  memtest2_datain_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_30_FFY_RST
    );
  memtest2_Mshreg_data4_10_59_685 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_10_net107,
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_30_FFY_RST,
      O => memtest2_Mshreg_data4_10_59
    );
  memtest2_n00511_4_686 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => memtest2_cs(0),
      ADR1 => VCC,
      ADR2 => memcontroller_Ker256691_O,
      ADR3 => VCC,
      O => memtest2_datain_30_FROM
    );
  memtest2_Mshreg_data4_10_srl_53 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_14,
      A1 => GLOBAL_LOGIC1_32,
      A2 => GLOBAL_LOGIC0_11,
      A3 => GLOBAL_LOGIC0_14,
      D => memtest2_ldata(10),
      CE => memtest2_n00511_4,
      CLK => clk,
      Q => memtest2_Mshreg_data4_10_net107
    );
  memtest2_datain_30_XUSED : X_BUF
    port map (
      I => memtest2_datain_30_FROM,
      O => memtest2_n00511_4
    );
  maccontrol_Mmux_n0023_Result_0_92_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_CHOICE1443,
      ADR1 => maccontrol_CHOICE1439,
      ADR2 => maccontrol_N30162,
      ADR3 => maccontrol_CHOICE1446,
      O => maccontrol_dout_0_FROM
    );
  maccontrol_Mmux_n0023_Result_0_92 : X_LUT4
    generic map(
      INIT => X"AAA8"
    )
    port map (
      ADR0 => maccontrol_N30238,
      ADR1 => maccontrol_CHOICE1426,
      ADR2 => maccontrol_CHOICE1433,
      ADR3 => maccontrol_Mmux_n0023_Result_0_92_SW0_O,
      O => maccontrol_Mmux_n0023_Result_0_92_O
    );
  maccontrol_dout_0_XUSED : X_BUF
    port map (
      I => maccontrol_dout_0_FROM,
      O => maccontrol_Mmux_n0023_Result_0_92_SW0_O
    );
  maccontrol_dout_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_14_FFY_RST
    );
  maccontrol_dout_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_1_58_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_14_FFY_RST,
      O => maccontrol_dout(1)
    );
  maccontrol_Mmux_n0023_Result_14_58 : X_LUT4
    generic map(
      INIT => X"D5C0"
    )
    port map (
      ADR0 => maccontrol_CHOICE1055,
      ADR1 => maccontrol_Mmux_n0023_Result_14_58_SW0_O,
      ADR2 => maccontrol_N30238,
      ADR3 => maccontrol_dout(13),
      O => maccontrol_Mmux_n0023_Result_14_58_O
    );
  maccontrol_Mmux_n0023_Result_1_58 : X_LUT4
    generic map(
      INIT => X"DC50"
    )
    port map (
      ADR0 => maccontrol_CHOICE1055,
      ADR1 => maccontrol_Mmux_n0023_Result_1_58_SW0_O,
      ADR2 => maccontrol_dout(0),
      ADR3 => maccontrol_N30238,
      O => maccontrol_Mmux_n0023_Result_1_58_O
    );
  maccontrol_dout_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_2_FFY_RST
    );
  maccontrol_dout_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_2_58_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_2_FFY_RST,
      O => maccontrol_dout(2)
    );
  maccontrol_Mmux_n0023_Result_2_58_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_CHOICE1471,
      ADR1 => maccontrol_CHOICE1474,
      ADR2 => maccontrol_Mmux_n0023_Result_2_26_SW0_O,
      ADR3 => maccontrol_Mmux_n0023_Result_2_26_2,
      O => maccontrol_dout_2_FROM
    );
  maccontrol_Mmux_n0023_Result_2_58 : X_LUT4
    generic map(
      INIT => X"F444"
    )
    port map (
      ADR0 => maccontrol_n00541_1,
      ADR1 => maccontrol_dout(1),
      ADR2 => maccontrol_N30238,
      ADR3 => maccontrol_Mmux_n0023_Result_2_58_SW0_O,
      O => maccontrol_Mmux_n0023_Result_2_58_O
    );
  maccontrol_dout_2_XUSED : X_BUF
    port map (
      I => maccontrol_dout_2_FROM,
      O => maccontrol_Mmux_n0023_Result_2_58_SW0_O
    );
  maccontrol_Ker302361 : X_LUT4
    generic map(
      INIT => X"0040"
    )
    port map (
      ADR0 => maccontrol_addr(5),
      ADR1 => maccontrol_N30218,
      ADR2 => maccontrol_sclkdeltall,
      ADR3 => maccontrol_bitcnt_90,
      O => maccontrol_dout_3_FROM
    );
  maccontrol_Mmux_n0023_Result_3_76 : X_LUT4
    generic map(
      INIT => X"DC50"
    )
    port map (
      ADR0 => maccontrol_n00541_1,
      ADR1 => maccontrol_N46555,
      ADR2 => maccontrol_dout(2),
      ADR3 => maccontrol_N30238,
      O => maccontrol_Mmux_n0023_Result_3_76_O
    );
  maccontrol_dout_3_XUSED : X_BUF
    port map (
      I => maccontrol_dout_3_FROM,
      O => maccontrol_N30238
    );
  maccontrol_dout_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_4_FFY_RST
    );
  maccontrol_dout_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_4_68_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_4_FFY_RST,
      O => maccontrol_dout(4)
    );
  maccontrol_Mmux_n0023_Result_4_32 : X_LUT4
    generic map(
      INIT => X"DCCC"
    )
    port map (
      ADR0 => maccontrol_addr_1_1,
      ADR1 => maccontrol_N46518,
      ADR2 => maccontrol_addr_0_1,
      ADR3 => maccontrol_CHOICE1269,
      O => maccontrol_dout_4_FROM
    );
  maccontrol_Mmux_n0023_Result_4_68 : X_LUT4
    generic map(
      INIT => X"FAF8"
    )
    port map (
      ADR0 => maccontrol_N30238,
      ADR1 => maccontrol_CHOICE1266,
      ADR2 => maccontrol_CHOICE1281,
      ADR3 => maccontrol_Mmux_n0023_Result_4_32_O,
      O => maccontrol_Mmux_n0023_Result_4_68_O
    );
  maccontrol_dout_4_XUSED : X_BUF
    port map (
      I => maccontrol_dout_4_FROM,
      O => maccontrol_Mmux_n0023_Result_4_32_O
    );
  maccontrol_Mmux_n0023_Result_5_58_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_CHOICE1507,
      ADR1 => maccontrol_CHOICE1510,
      ADR2 => maccontrol_Mmux_n0023_Result_5_26_SW0_O,
      ADR3 => maccontrol_Mmux_n0023_Result_5_26_2,
      O => maccontrol_dout_5_FROM
    );
  maccontrol_Mmux_n0023_Result_5_58 : X_LUT4
    generic map(
      INIT => X"AE0C"
    )
    port map (
      ADR0 => maccontrol_N30238,
      ADR1 => maccontrol_dout(4),
      ADR2 => maccontrol_n00541_1,
      ADR3 => maccontrol_Mmux_n0023_Result_5_58_SW0_O,
      O => maccontrol_Mmux_n0023_Result_5_58_O
    );
  maccontrol_dout_5_XUSED : X_BUF
    port map (
      I => maccontrol_dout_5_FROM,
      O => maccontrol_Mmux_n0023_Result_5_58_SW0_O
    );
  maccontrol_Mmux_n0023_Result_8_58 : X_LUT4
    generic map(
      INIT => X"CE0A"
    )
    port map (
      ADR0 => maccontrol_dout(7),
      ADR1 => maccontrol_N30238,
      ADR2 => maccontrol_n00541_1,
      ADR3 => maccontrol_Mmux_n0023_Result_8_58_SW0_O,
      O => maccontrol_Mmux_n0023_Result_8_58_O
    );
  maccontrol_Mmux_n0023_Result_6_58 : X_LUT4
    generic map(
      INIT => X"CE0A"
    )
    port map (
      ADR0 => maccontrol_dout(5),
      ADR1 => maccontrol_Mmux_n0023_Result_6_58_SW0_O,
      ADR2 => maccontrol_n00541_1,
      ADR3 => maccontrol_N30238,
      O => maccontrol_Mmux_n0023_Result_6_58_O
    );
  maccontrol_dout_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_7_FFY_RST
    );
  maccontrol_dout_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_7_76_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_7_FFY_RST,
      O => maccontrol_dout(7)
    );
  maccontrol_Mmux_n0023_Result_7_76_SW0 : X_LUT4
    generic map(
      INIT => X"FEFA"
    )
    port map (
      ADR0 => maccontrol_CHOICE1364,
      ADR1 => maccontrol_n00691_1,
      ADR2 => maccontrol_CHOICE1376,
      ADR3 => maccontrol_phyaddr(7),
      O => maccontrol_dout_7_FROM
    );
  maccontrol_Mmux_n0023_Result_7_76 : X_LUT4
    generic map(
      INIT => X"F222"
    )
    port map (
      ADR0 => maccontrol_dout(6),
      ADR1 => maccontrol_n00541_1,
      ADR2 => maccontrol_N30238,
      ADR3 => maccontrol_Mmux_n0023_Result_7_76_SW0_O,
      O => maccontrol_Mmux_n0023_Result_7_76_O
    );
  maccontrol_dout_7_XUSED : X_BUF
    port map (
      I => maccontrol_dout_7_FROM,
      O => maccontrol_Mmux_n0023_Result_7_76_SW0_O
    );
  memtest2_n01161 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => memtest2_cs(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_Ker256691_O,
      O => d2_0_GROM
    );
  d2_0_YUSED : X_BUF
    port map (
      I => d2_0_GROM,
      O => memtest2_n0116
    );
  maccontrol_dout_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_9_FFY_RST
    );
  maccontrol_dout_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_9_68_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_9_FFY_RST,
      O => maccontrol_dout(9)
    );
  maccontrol_Mmux_n0023_Result_9_32 : X_LUT4
    generic map(
      INIT => X"BAAA"
    )
    port map (
      ADR0 => maccontrol_N46526,
      ADR1 => maccontrol_addr_1_1,
      ADR2 => maccontrol_addr_0_1,
      ADR3 => maccontrol_CHOICE1288,
      O => maccontrol_dout_9_FROM
    );
  maccontrol_Mmux_n0023_Result_9_68 : X_LUT4
    generic map(
      INIT => X"EEEA"
    )
    port map (
      ADR0 => maccontrol_CHOICE1300,
      ADR1 => maccontrol_N30238,
      ADR2 => maccontrol_CHOICE1285,
      ADR3 => maccontrol_Mmux_n0023_Result_9_32_O,
      O => maccontrol_Mmux_n0023_Result_9_68_O
    );
  maccontrol_dout_9_XUSED : X_BUF
    port map (
      I => maccontrol_dout_9_FROM,
      O => maccontrol_Mmux_n0023_Result_9_32_O
    );
  memtest2_n01161_1_687 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_Ker256691_O,
      ADR3 => memtest2_cs(0),
      O => d2_3_GROM
    );
  d2_3_YUSED : X_BUF
    port map (
      I => d2_3_GROM,
      O => memtest2_n01161_1
    );
  memtest2_Mshreg_data4_13_56_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_13_56_FFY_RST
    );
  memtest2_Mshreg_data4_20_49_688 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_20_net87,
      CE => memtest2_n00511_3,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_13_56_FFY_RST,
      O => memtest2_Mshreg_data4_20_49
    );
  memtest2_n00511_3_689 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cs(0),
      ADR2 => VCC,
      ADR3 => memcontroller_Ker256691_O,
      O => memtest2_Mshreg_data4_13_56_FROM
    );
  memtest2_Mshreg_data4_20_srl_43 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_27,
      A1 => GLOBAL_LOGIC1_11,
      A2 => GLOBAL_LOGIC0_45,
      A3 => GLOBAL_LOGIC0_45,
      D => memtest2_ldata(20),
      CE => memtest2_n00511_3,
      CLK => clk,
      Q => memtest2_Mshreg_data4_20_net87
    );
  memtest2_Mshreg_data4_13_56_XUSED : X_BUF
    port map (
      I => memtest2_Mshreg_data4_13_56_FROM,
      O => memtest2_n00511_3
    );
  memtest2_Mshreg_data4_21_48_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_21_48_FFY_RST
    );
  memtest2_Mshreg_data4_24_45_690 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_24_net79,
      CE => memtest2_n00511_2,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_21_48_FFY_RST,
      O => memtest2_Mshreg_data4_24_45
    );
  memtest2_n00511_2_691 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_Ker256691_O,
      ADR3 => memtest2_cs(0),
      O => memtest2_Mshreg_data4_21_48_FROM
    );
  memtest2_Mshreg_data4_24_srl_39 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_25,
      A1 => GLOBAL_LOGIC1_29,
      A2 => GLOBAL_LOGIC0_25,
      A3 => GLOBAL_LOGIC0_25,
      D => memtest2_ldata(24),
      CE => memtest2_n00511_2,
      CLK => clk,
      Q => memtest2_Mshreg_data4_24_net79
    );
  memtest2_Mshreg_data4_21_48_XUSED : X_BUF
    port map (
      I => memtest2_Mshreg_data4_21_48_FROM,
      O => memtest2_n00511_2
    );
  maccontrol_Mmux_n0023_Result_13_18 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(29),
      ADR1 => maccontrol_phydo(13),
      ADR2 => maccontrol_N30192,
      ADR3 => maccontrol_N30212,
      O => maccontrol_Mmux_n0023_Result_13_18_O_FROM
    );
  maccontrol_Mmux_n0023_Result_13_32_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n0067,
      ADR1 => maccontrol_N30292,
      ADR2 => maccontrol_phystat(13),
      ADR3 => maccontrol_Mmux_n0023_Result_13_18_O,
      O => maccontrol_Mmux_n0023_Result_13_18_O_GROM
    );
  maccontrol_Mmux_n0023_Result_13_18_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_13_18_O_FROM,
      O => maccontrol_Mmux_n0023_Result_13_18_O
    );
  maccontrol_Mmux_n0023_Result_13_18_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_13_18_O_GROM,
      O => maccontrol_N46514
    );
  maccontrol_dout_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_10_FFY_RST
    );
  maccontrol_dout_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_10_58_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_10_FFY_RST,
      O => maccontrol_dout(10)
    );
  maccontrol_Mmux_n0023_Result_10_58_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_Mmux_n0023_Result_10_26_SW0_O,
      ADR1 => maccontrol_CHOICE1543,
      ADR2 => maccontrol_CHOICE1546,
      ADR3 => maccontrol_Mmux_n0023_Result_10_26_2,
      O => maccontrol_dout_10_FROM
    );
  maccontrol_Mmux_n0023_Result_10_58 : X_LUT4
    generic map(
      INIT => X"BA30"
    )
    port map (
      ADR0 => maccontrol_N30238,
      ADR1 => maccontrol_CHOICE1055,
      ADR2 => maccontrol_dout(9),
      ADR3 => maccontrol_Mmux_n0023_Result_10_58_SW0_O,
      O => maccontrol_Mmux_n0023_Result_10_58_O
    );
  maccontrol_dout_10_XUSED : X_BUF
    port map (
      I => maccontrol_dout_10_FROM,
      O => maccontrol_Mmux_n0023_Result_10_58_SW0_O
    );
  memcontroller_addr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_8_OD,
      CE => MA_8_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_8_OFF_RST,
      O => memcontroller_ADDREXT(8)
    );
  MA_8_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_8_OFF_RST
    );
  maccontrol_Ker303141_2_692 : X_LUT4
    generic map(
      INIT => X"0010"
    )
    port map (
      ADR0 => maccontrol_N42043,
      ADR1 => maccontrol_bitcnt_89,
      ADR2 => maccontrol_bitcnt_88,
      ADR3 => maccontrol_N46368,
      O => maccontrol_PHY_status_phyaddrws_FROM
    );
  maccontrol_PHY_status_n00151 : X_LUT4
    generic map(
      INIT => X"0E0A"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd1,
      ADR1 => maccontrol_n0069,
      ADR2 => maccontrol_PHY_status_n00151_1,
      ADR3 => maccontrol_Ker303141_2,
      O => maccontrol_PHY_status_phyaddrws_GROM
    );
  maccontrol_PHY_status_phyaddrws_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_phyaddrws_FROM,
      O => maccontrol_Ker303141_2
    );
  maccontrol_PHY_status_phyaddrws_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_phyaddrws_GROM,
      O => maccontrol_PHY_status_n00151_O
    );
  maccontrol_PHY_status_phyaddrws_BYMUX : X_INV
    port map (
      I => maccontrol_PHY_status_cs_FFd1,
      O => maccontrol_PHY_status_phyaddrws_BYMUXNOT
    );
  maccontrol_dout_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_11_FFY_RST
    );
  maccontrol_dout_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_11_76_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_11_FFY_RST,
      O => maccontrol_dout(11)
    );
  maccontrol_Mmux_n0023_Result_11_76_SW0 : X_LUT4
    generic map(
      INIT => X"FEFA"
    )
    port map (
      ADR0 => maccontrol_CHOICE1385,
      ADR1 => maccontrol_phyaddr(11),
      ADR2 => maccontrol_CHOICE1397,
      ADR3 => maccontrol_n0069,
      O => maccontrol_dout_11_FROM
    );
  maccontrol_Mmux_n0023_Result_11_76 : X_LUT4
    generic map(
      INIT => X"DC50"
    )
    port map (
      ADR0 => maccontrol_CHOICE1055,
      ADR1 => maccontrol_N30238,
      ADR2 => maccontrol_dout(10),
      ADR3 => maccontrol_Mmux_n0023_Result_11_76_SW0_O,
      O => maccontrol_Mmux_n0023_Result_11_76_O
    );
  maccontrol_dout_11_XUSED : X_BUF
    port map (
      I => maccontrol_dout_11_FROM,
      O => maccontrol_Mmux_n0023_Result_11_76_SW0_O
    );
  maccontrol_Mmux_n0023_Result_12_32 : X_LUT4
    generic map(
      INIT => X"DCCC"
    )
    port map (
      ADR0 => maccontrol_addr_1_1,
      ADR1 => maccontrol_N46522,
      ADR2 => maccontrol_CHOICE1307,
      ADR3 => maccontrol_addr_0_1,
      O => maccontrol_dout_12_FROM
    );
  maccontrol_Mmux_n0023_Result_12_68 : X_LUT4
    generic map(
      INIT => X"FAEA"
    )
    port map (
      ADR0 => maccontrol_CHOICE1319,
      ADR1 => maccontrol_CHOICE1304,
      ADR2 => maccontrol_N30238,
      ADR3 => maccontrol_Mmux_n0023_Result_12_32_O,
      O => maccontrol_Mmux_n0023_Result_12_68_O
    );
  maccontrol_dout_12_XUSED : X_BUF
    port map (
      I => maccontrol_dout_12_FROM,
      O => maccontrol_Mmux_n0023_Result_12_32_O
    );
  maccontrol_Mmux_n0023_Result_20_22_SW0 : X_LUT4
    generic map(
      INIT => X"FAF0"
    )
    port map (
      ADR0 => maccontrol_n00691_1,
      ADR1 => VCC,
      ADR2 => maccontrol_CHOICE1120,
      ADR3 => maccontrol_phyaddr(20),
      O => maccontrol_dout_20_FROM
    );
  maccontrol_Mmux_n0023_Result_20_22 : X_LUT4
    generic map(
      INIT => X"F444"
    )
    port map (
      ADR0 => maccontrol_CHOICE1055,
      ADR1 => maccontrol_dout(19),
      ADR2 => maccontrol_N30238,
      ADR3 => maccontrol_Mmux_n0023_Result_20_22_SW0_O,
      O => maccontrol_Mmux_n0023_Result_20_22_O
    );
  maccontrol_dout_20_XUSED : X_BUF
    port map (
      I => maccontrol_dout_20_FROM,
      O => maccontrol_Mmux_n0023_Result_20_22_SW0_O
    );
  maccontrol_Mmux_n0023_Result_21_12 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n00671_1,
      ADR1 => maccontrol_N30212,
      ADR2 => maccontrol_phystat(21),
      ADR3 => maccontrol_CHOICE1245,
      O => maccontrol_dout_21_FROM
    );
  maccontrol_Mmux_n0023_Result_21_36 : X_LUT4
    generic map(
      INIT => X"EEEA"
    )
    port map (
      ADR0 => maccontrol_CHOICE1251,
      ADR1 => maccontrol_N30238,
      ADR2 => maccontrol_N30162,
      ADR3 => maccontrol_Mmux_n0023_Result_21_12_O,
      O => maccontrol_Mmux_n0023_Result_21_36_O
    );
  maccontrol_dout_21_XUSED : X_BUF
    port map (
      I => maccontrol_dout_21_FROM,
      O => maccontrol_Mmux_n0023_Result_21_12_O
    );
  maccontrol_Mmux_n0023_Result_13_32 : X_LUT4
    generic map(
      INIT => X"F0F8"
    )
    port map (
      ADR0 => maccontrol_CHOICE1326,
      ADR1 => maccontrol_addr_0_1,
      ADR2 => maccontrol_N46514,
      ADR3 => maccontrol_addr_1_1,
      O => maccontrol_dout_13_FROM
    );
  maccontrol_Mmux_n0023_Result_13_68 : X_LUT4
    generic map(
      INIT => X"FAEA"
    )
    port map (
      ADR0 => maccontrol_CHOICE1338,
      ADR1 => maccontrol_CHOICE1323,
      ADR2 => maccontrol_N30238,
      ADR3 => maccontrol_Mmux_n0023_Result_13_32_O,
      O => maccontrol_Mmux_n0023_Result_13_68_O
    );
  maccontrol_dout_13_XUSED : X_BUF
    port map (
      I => maccontrol_dout_13_FROM,
      O => maccontrol_Mmux_n0023_Result_13_32_O
    );
  maccontrol_Mmux_n0023_Result_30_22_SW0 : X_LUT4
    generic map(
      INIT => X"FCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_CHOICE1165,
      ADR2 => maccontrol_phyaddr(30),
      ADR3 => maccontrol_n00691_1,
      O => maccontrol_dout_30_FROM
    );
  maccontrol_Mmux_n0023_Result_30_22 : X_LUT4
    generic map(
      INIT => X"BA30"
    )
    port map (
      ADR0 => maccontrol_N30238,
      ADR1 => maccontrol_n00541_1,
      ADR2 => maccontrol_dout(29),
      ADR3 => maccontrol_Mmux_n0023_Result_30_22_SW0_O,
      O => maccontrol_Mmux_n0023_Result_30_22_O
    );
  maccontrol_dout_30_XUSED : X_BUF
    port map (
      I => maccontrol_dout_30_FROM,
      O => maccontrol_Mmux_n0023_Result_30_22_SW0_O
    );
  maccontrol_Mmux_n0023_Result_22_22_SW0 : X_LUT4
    generic map(
      INIT => X"FAAA"
    )
    port map (
      ADR0 => maccontrol_CHOICE1129,
      ADR1 => VCC,
      ADR2 => maccontrol_phyaddr(22),
      ADR3 => maccontrol_n00691_1,
      O => maccontrol_dout_22_FROM
    );
  maccontrol_Mmux_n0023_Result_22_22 : X_LUT4
    generic map(
      INIT => X"AE0C"
    )
    port map (
      ADR0 => maccontrol_N30238,
      ADR1 => maccontrol_dout(21),
      ADR2 => maccontrol_CHOICE1055,
      ADR3 => maccontrol_Mmux_n0023_Result_22_22_SW0_O,
      O => maccontrol_Mmux_n0023_Result_22_22_O
    );
  maccontrol_dout_22_XUSED : X_BUF
    port map (
      I => maccontrol_dout_22_FROM,
      O => maccontrol_Mmux_n0023_Result_22_22_SW0_O
    );
  maccontrol_Mmux_n0023_Result_23_25_SW0 : X_LUT4
    generic map(
      INIT => X"0105"
    )
    port map (
      ADR0 => maccontrol_CHOICE1204,
      ADR1 => maccontrol_n00671_1,
      ADR2 => maccontrol_n0068,
      ADR3 => maccontrol_phystat(23),
      O => maccontrol_dout_23_FROM
    );
  maccontrol_Mmux_n0023_Result_23_25 : X_LUT4
    generic map(
      INIT => X"5072"
    )
    port map (
      ADR0 => maccontrol_CHOICE1055,
      ADR1 => maccontrol_addr(5),
      ADR2 => maccontrol_dout(22),
      ADR3 => maccontrol_Mmux_n0023_Result_23_25_SW0_O,
      O => maccontrol_Mmux_n0023_Result_23_25_O
    );
  maccontrol_dout_23_XUSED : X_BUF
    port map (
      I => maccontrol_dout_23_FROM,
      O => maccontrol_Mmux_n0023_Result_23_25_SW0_O
    );
  maccontrol_Mmux_n0023_Result_31_25_SW0 : X_LUT4
    generic map(
      INIT => X"0103"
    )
    port map (
      ADR0 => maccontrol_phystat(31),
      ADR1 => maccontrol_CHOICE1184,
      ADR2 => maccontrol_n0068,
      ADR3 => maccontrol_n00671_1,
      O => maccontrol_dout_31_FROM
    );
  maccontrol_Mmux_n0023_Result_31_25 : X_LUT4
    generic map(
      INIT => X"0C5C"
    )
    port map (
      ADR0 => maccontrol_addr(5),
      ADR1 => maccontrol_dout(30),
      ADR2 => maccontrol_n00541_1,
      ADR3 => maccontrol_Mmux_n0023_Result_31_25_SW0_O,
      O => maccontrol_Mmux_n0023_Result_31_25_O
    );
  maccontrol_dout_31_XUSED : X_BUF
    port map (
      I => maccontrol_dout_31_FROM,
      O => maccontrol_Mmux_n0023_Result_31_25_SW0_O
    );
  maccontrol_Mmux_n0023_Result_15_76_SW0 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => maccontrol_phyaddr(15),
      ADR1 => maccontrol_n00691_1,
      ADR2 => maccontrol_CHOICE1406,
      ADR3 => maccontrol_CHOICE1418,
      O => maccontrol_dout_15_FROM
    );
  maccontrol_Mmux_n0023_Result_15_76 : X_LUT4
    generic map(
      INIT => X"8F88"
    )
    port map (
      ADR0 => maccontrol_N30238,
      ADR1 => maccontrol_Mmux_n0023_Result_15_76_SW0_O,
      ADR2 => maccontrol_CHOICE1055,
      ADR3 => maccontrol_dout(14),
      O => maccontrol_Mmux_n0023_Result_15_76_O
    );
  maccontrol_dout_15_XUSED : X_BUF
    port map (
      I => maccontrol_dout_15_FROM,
      O => maccontrol_Mmux_n0023_Result_15_76_SW0_O
    );
  maccontrol_Mmux_n0023_Result_24_12 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_CHOICE1256,
      ADR1 => maccontrol_N30212,
      ADR2 => maccontrol_n00671_1,
      ADR3 => maccontrol_phystat(24),
      O => maccontrol_dout_24_FROM
    );
  maccontrol_Mmux_n0023_Result_24_36 : X_LUT4
    generic map(
      INIT => X"EEEC"
    )
    port map (
      ADR0 => maccontrol_N30238,
      ADR1 => maccontrol_CHOICE1262,
      ADR2 => maccontrol_N30162,
      ADR3 => maccontrol_Mmux_n0023_Result_24_12_O,
      O => maccontrol_Mmux_n0023_Result_24_36_O
    );
  maccontrol_dout_24_XUSED : X_BUF
    port map (
      I => maccontrol_dout_24_FROM,
      O => maccontrol_Mmux_n0023_Result_24_12_O
    );
  maccontrol_Mmux_n0023_Result_16_12 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n00671_1,
      ADR1 => maccontrol_N30212,
      ADR2 => maccontrol_phystat(16),
      ADR3 => maccontrol_CHOICE1223,
      O => maccontrol_dout_16_FROM
    );
  maccontrol_Mmux_n0023_Result_16_36 : X_LUT4
    generic map(
      INIT => X"FCF8"
    )
    port map (
      ADR0 => maccontrol_N30162,
      ADR1 => maccontrol_N30238,
      ADR2 => maccontrol_CHOICE1229,
      ADR3 => maccontrol_Mmux_n0023_Result_16_12_O,
      O => maccontrol_Mmux_n0023_Result_16_36_O
    );
  maccontrol_dout_16_XUSED : X_BUF
    port map (
      I => maccontrol_dout_16_FROM,
      O => maccontrol_Mmux_n0023_Result_16_12_O
    );
  maccontrol_Mmux_n0023_Result_17_12 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_n00671_1,
      ADR1 => maccontrol_phystat(17),
      ADR2 => maccontrol_N30212,
      ADR3 => maccontrol_CHOICE1234,
      O => maccontrol_dout_17_FROM
    );
  maccontrol_Mmux_n0023_Result_17_36 : X_LUT4
    generic map(
      INIT => X"FAEA"
    )
    port map (
      ADR0 => maccontrol_CHOICE1240,
      ADR1 => maccontrol_N30162,
      ADR2 => maccontrol_N30238,
      ADR3 => maccontrol_Mmux_n0023_Result_17_12_O,
      O => maccontrol_Mmux_n0023_Result_17_36_O
    );
  maccontrol_dout_17_XUSED : X_BUF
    port map (
      I => maccontrol_dout_17_FROM,
      O => maccontrol_Mmux_n0023_Result_17_12_O
    );
  maccontrol_Mmux_n0023_Result_25_22_SW0 : X_LUT4
    generic map(
      INIT => X"FF88"
    )
    port map (
      ADR0 => maccontrol_phyaddr(25),
      ADR1 => maccontrol_n00691_1,
      ADR2 => VCC,
      ADR3 => maccontrol_CHOICE1138,
      O => maccontrol_dout_25_FROM
    );
  maccontrol_Mmux_n0023_Result_25_22 : X_LUT4
    generic map(
      INIT => X"CE0A"
    )
    port map (
      ADR0 => maccontrol_dout(24),
      ADR1 => maccontrol_N30238,
      ADR2 => maccontrol_CHOICE1055,
      ADR3 => maccontrol_Mmux_n0023_Result_25_22_SW0_O,
      O => maccontrol_Mmux_n0023_Result_25_22_O
    );
  maccontrol_dout_25_XUSED : X_BUF
    port map (
      I => maccontrol_dout_25_FROM,
      O => maccontrol_Mmux_n0023_Result_25_22_SW0_O
    );
  maccontrol_Mmux_n0023_Result_18_22_SW0 : X_LUT4
    generic map(
      INIT => X"FF88"
    )
    port map (
      ADR0 => maccontrol_phyaddr(18),
      ADR1 => maccontrol_n00691_1,
      ADR2 => VCC,
      ADR3 => maccontrol_CHOICE1111,
      O => maccontrol_dout_18_FROM
    );
  maccontrol_Mmux_n0023_Result_18_22 : X_LUT4
    generic map(
      INIT => X"F444"
    )
    port map (
      ADR0 => maccontrol_CHOICE1055,
      ADR1 => maccontrol_dout(17),
      ADR2 => maccontrol_N30238,
      ADR3 => maccontrol_Mmux_n0023_Result_18_22_SW0_O,
      O => maccontrol_Mmux_n0023_Result_18_22_O
    );
  maccontrol_dout_18_XUSED : X_BUF
    port map (
      I => maccontrol_dout_18_FROM,
      O => maccontrol_Mmux_n0023_Result_18_22_SW0_O
    );
  maccontrol_Mmux_n0023_Result_26_22_SW0 : X_LUT4
    generic map(
      INIT => X"FCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_CHOICE1147,
      ADR2 => maccontrol_n00691_1,
      ADR3 => maccontrol_phyaddr(26),
      O => maccontrol_dout_26_FROM
    );
  maccontrol_Mmux_n0023_Result_26_22 : X_LUT4
    generic map(
      INIT => X"F222"
    )
    port map (
      ADR0 => maccontrol_dout(25),
      ADR1 => maccontrol_n00541_1,
      ADR2 => maccontrol_N30238,
      ADR3 => maccontrol_Mmux_n0023_Result_26_22_SW0_O,
      O => maccontrol_Mmux_n0023_Result_26_22_O
    );
  maccontrol_dout_26_XUSED : X_BUF
    port map (
      I => maccontrol_dout_26_FROM,
      O => maccontrol_Mmux_n0023_Result_26_22_SW0_O
    );
  maccontrol_Mmux_n0023_Result_27_25_SW0 : X_LUT4
    generic map(
      INIT => X"0013"
    )
    port map (
      ADR0 => maccontrol_phystat(27),
      ADR1 => maccontrol_n0068,
      ADR2 => maccontrol_n00671_1,
      ADR3 => maccontrol_CHOICE1214,
      O => maccontrol_dout_27_FROM
    );
  maccontrol_Mmux_n0023_Result_27_25 : X_LUT4
    generic map(
      INIT => X"0C5C"
    )
    port map (
      ADR0 => maccontrol_addr(5),
      ADR1 => maccontrol_dout(26),
      ADR2 => maccontrol_n00541_1,
      ADR3 => maccontrol_Mmux_n0023_Result_27_25_SW0_O,
      O => maccontrol_Mmux_n0023_Result_27_25_O
    );
  maccontrol_dout_27_XUSED : X_BUF
    port map (
      I => maccontrol_dout_27_FROM,
      O => maccontrol_Mmux_n0023_Result_27_25_SW0_O
    );
  maccontrol_Mmux_n0023_Result_19_25_SW0 : X_LUT4
    generic map(
      INIT => X"0111"
    )
    port map (
      ADR0 => maccontrol_n0068,
      ADR1 => maccontrol_CHOICE1194,
      ADR2 => maccontrol_n00671_1,
      ADR3 => maccontrol_phystat(19),
      O => maccontrol_dout_19_FROM
    );
  maccontrol_Mmux_n0023_Result_19_25 : X_LUT4
    generic map(
      INIT => X"444E"
    )
    port map (
      ADR0 => maccontrol_CHOICE1055,
      ADR1 => maccontrol_dout(18),
      ADR2 => maccontrol_addr(5),
      ADR3 => maccontrol_Mmux_n0023_Result_19_25_SW0_O,
      O => maccontrol_Mmux_n0023_Result_19_25_O
    );
  maccontrol_dout_19_XUSED : X_BUF
    port map (
      I => maccontrol_dout_19_FROM,
      O => maccontrol_Mmux_n0023_Result_19_25_SW0_O
    );
  memcontroller_addr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_9_OD,
      CE => MA_9_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_9_OFF_RST,
      O => memcontroller_ADDREXT(9)
    );
  MA_9_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_9_OFF_RST
    );
  maccontrol_Mmux_n0023_Result_28_22_SW0 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => maccontrol_phyaddr(28),
      ADR1 => VCC,
      ADR2 => maccontrol_n00691_1,
      ADR3 => maccontrol_CHOICE1156,
      O => maccontrol_dout_28_FROM
    );
  maccontrol_Mmux_n0023_Result_28_22 : X_LUT4
    generic map(
      INIT => X"CE0A"
    )
    port map (
      ADR0 => maccontrol_dout(27),
      ADR1 => maccontrol_N30238,
      ADR2 => maccontrol_n00541_1,
      ADR3 => maccontrol_Mmux_n0023_Result_28_22_SW0_O,
      O => maccontrol_Mmux_n0023_Result_28_22_O
    );
  maccontrol_dout_28_XUSED : X_BUF
    port map (
      I => maccontrol_dout_28_FROM,
      O => maccontrol_Mmux_n0023_Result_28_22_SW0_O
    );
  maccontrol_Mmux_n0023_Result_29_22_SW0 : X_LUT4
    generic map(
      INIT => X"FF88"
    )
    port map (
      ADR0 => maccontrol_phyaddr(29),
      ADR1 => maccontrol_n00691_1,
      ADR2 => VCC,
      ADR3 => maccontrol_CHOICE1174,
      O => maccontrol_dout_29_FROM
    );
  maccontrol_Mmux_n0023_Result_29_22 : X_LUT4
    generic map(
      INIT => X"DC50"
    )
    port map (
      ADR0 => maccontrol_n00541_1,
      ADR1 => maccontrol_N30238,
      ADR2 => maccontrol_dout(28),
      ADR3 => maccontrol_Mmux_n0023_Result_29_22_SW0_O,
      O => maccontrol_Mmux_n0023_Result_29_22_O
    );
  maccontrol_dout_29_XUSED : X_BUF
    port map (
      I => maccontrol_dout_29_FROM,
      O => maccontrol_Mmux_n0023_Result_29_22_SW0_O
    );
  maccontrol_Mmux_n0023_Result_6_26_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_n0070,
      ADR1 => maccontrol_phydi(6),
      ADR2 => maccontrol_phydo(6),
      ADR3 => maccontrol_n0071,
      O => maccontrol_Mmux_n0023_Result_6_26_SW0_O_FROM
    );
  maccontrol_Mmux_n0023_Result_6_58_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_Mmux_n0023_Result_6_26_2,
      ADR1 => maccontrol_CHOICE1492,
      ADR2 => maccontrol_CHOICE1489,
      ADR3 => maccontrol_Mmux_n0023_Result_6_26_SW0_O,
      O => maccontrol_Mmux_n0023_Result_6_26_SW0_O_GROM
    );
  maccontrol_Mmux_n0023_Result_6_26_SW0_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_6_26_SW0_O_FROM,
      O => maccontrol_Mmux_n0023_Result_6_26_SW0_O
    );
  maccontrol_Mmux_n0023_Result_6_26_SW0_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_6_26_SW0_O_GROM,
      O => maccontrol_Mmux_n0023_Result_6_58_SW0_O
    );
  maccontrol_n00671 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => maccontrol_N30292,
      ADR1 => maccontrol_addr(4),
      ADR2 => maccontrol_addr(2),
      ADR3 => maccontrol_addr(3),
      O => maccontrol_n0067_FROM
    );
  maccontrol_Mmux_n0023_Result_2_9 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(18),
      ADR1 => maccontrol_phystat(2),
      ADR2 => maccontrol_n0084,
      ADR3 => maccontrol_n0067,
      O => maccontrol_n0067_GROM
    );
  maccontrol_n0067_XUSED : X_BUF
    port map (
      I => maccontrol_n0067_FROM,
      O => maccontrol_n0067
    );
  maccontrol_n0067_YUSED : X_BUF
    port map (
      I => maccontrol_n0067_GROM,
      O => maccontrol_CHOICE1474
    );
  maccontrol_n00691_1_693 : X_LUT4
    generic map(
      INIT => X"0200"
    )
    port map (
      ADR0 => maccontrol_addr(3),
      ADR1 => maccontrol_addr(2),
      ADR2 => maccontrol_addr(4),
      ADR3 => maccontrol_N30305,
      O => maccontrol_n00691_1_FROM
    );
  maccontrol_Mmux_n0023_Result_4_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_phyaddr(4),
      ADR1 => maccontrol_n0085,
      ADR2 => maccontrol_lmacaddr(36),
      ADR3 => maccontrol_n00691_1,
      O => maccontrol_n00691_1_GROM
    );
  maccontrol_n00691_1_XUSED : X_BUF
    port map (
      I => maccontrol_n00691_1_FROM,
      O => maccontrol_n00691_1
    );
  maccontrol_n00691_1_YUSED : X_BUF
    port map (
      I => maccontrol_n00691_1_GROM,
      O => maccontrol_CHOICE1266
    );
  maccontrol_n00831 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_addr(3),
      ADR1 => maccontrol_N30285,
      ADR2 => maccontrol_addr(4),
      ADR3 => maccontrol_addr(2),
      O => maccontrol_n0083_FROM
    );
  maccontrol_Mmux_n0023_Result_5_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n0085,
      ADR1 => maccontrol_lmacaddr(5),
      ADR2 => maccontrol_lmacaddr(37),
      ADR3 => maccontrol_n0083,
      O => maccontrol_n0083_GROM
    );
  maccontrol_n0083_XUSED : X_BUF
    port map (
      I => maccontrol_n0083_FROM,
      O => maccontrol_n0083
    );
  maccontrol_n0083_YUSED : X_BUF
    port map (
      I => maccontrol_n0083_GROM,
      O => maccontrol_CHOICE1507
    );
  memcontroller_qn_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(0),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_0_IFF_RST,
      O => memcontroller_qn(0)
    );
  MD_0_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_0_IFF_RST
    );
  maccontrol_Ker301901 : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_addr(3),
      ADR2 => maccontrol_addr(2),
      ADR3 => maccontrol_addr(4),
      O => maccontrol_N30192_FROM
    );
  maccontrol_Mmux_n0023_Result_4_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_phydi(4),
      ADR1 => maccontrol_N30212,
      ADR2 => maccontrol_lmacaddr(4),
      ADR3 => maccontrol_N30192,
      O => maccontrol_N30192_GROM
    );
  maccontrol_N30192_XUSED : X_BUF
    port map (
      I => maccontrol_N30192_FROM,
      O => maccontrol_N30192
    );
  maccontrol_N30192_YUSED : X_BUF
    port map (
      I => maccontrol_N30192_GROM,
      O => maccontrol_CHOICE1269
    );
  maccontrol_n00671_1_694 : X_LUT4
    generic map(
      INIT => X"0004"
    )
    port map (
      ADR0 => maccontrol_addr(3),
      ADR1 => maccontrol_N30292,
      ADR2 => maccontrol_addr(2),
      ADR3 => maccontrol_addr(4),
      O => maccontrol_n00671_1_FROM
    );
  maccontrol_Mmux_n0023_Result_6_9 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n0084,
      ADR1 => maccontrol_phystat(6),
      ADR2 => maccontrol_lmacaddr(22),
      ADR3 => maccontrol_n00671_1,
      O => maccontrol_n00671_1_GROM
    );
  maccontrol_n00671_1_XUSED : X_BUF
    port map (
      I => maccontrol_n00671_1_FROM,
      O => maccontrol_n00671_1
    );
  maccontrol_n00671_1_YUSED : X_BUF
    port map (
      I => maccontrol_n00671_1_GROM,
      O => maccontrol_CHOICE1492
    );
  memtest2_Ker2265830 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => memtest2_cnt(1),
      ADR1 => memtest2_cnt(15),
      ADR2 => memtest2_cnt(2),
      ADR3 => memtest2_cnt(14),
      O => memtest2_Ker2265830_O_FROM
    );
  memtest2_Ker2265849 : X_LUT4
    generic map(
      INIT => X"0400"
    )
    port map (
      ADR0 => memtest2_cnt(0),
      ADR1 => memtest2_Ker2265849_2,
      ADR2 => memtest2_cnt(16),
      ADR3 => memtest2_Ker2265830_O,
      O => memtest2_Ker2265830_O_GROM
    );
  memtest2_Ker2265830_O_XUSED : X_BUF
    port map (
      I => memtest2_Ker2265830_O_FROM,
      O => memtest2_Ker2265830_O
    );
  memtest2_Ker2265830_O_YUSED : X_BUF
    port map (
      I => memtest2_Ker2265830_O_GROM,
      O => memtest2_N22660
    );
  maccontrol_Mmux_n0023_Result_9_18 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_N30192,
      ADR1 => maccontrol_lmacaddr(25),
      ADR2 => maccontrol_phydo(9),
      ADR3 => maccontrol_N30212,
      O => maccontrol_Mmux_n0023_Result_9_18_O_FROM
    );
  maccontrol_Mmux_n0023_Result_9_32_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_phystat(9),
      ADR1 => maccontrol_n00671_1,
      ADR2 => maccontrol_N30292,
      ADR3 => maccontrol_Mmux_n0023_Result_9_18_O,
      O => maccontrol_Mmux_n0023_Result_9_18_O_GROM
    );
  maccontrol_Mmux_n0023_Result_9_18_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_9_18_O_FROM,
      O => maccontrol_Mmux_n0023_Result_9_18_O
    );
  maccontrol_Mmux_n0023_Result_9_18_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_9_18_O_GROM,
      O => maccontrol_N46526
    );
  maccontrol_Mmux_n0023_Result_14_26_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_phydi(14),
      ADR1 => maccontrol_phydo(14),
      ADR2 => maccontrol_n0070,
      ADR3 => maccontrol_n0071,
      O => maccontrol_Mmux_n0023_Result_14_26_SW0_O_FROM
    );
  maccontrol_Mmux_n0023_Result_14_58_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_Mmux_n0023_Result_14_26_2,
      ADR1 => maccontrol_CHOICE1561,
      ADR2 => maccontrol_CHOICE1564,
      ADR3 => maccontrol_Mmux_n0023_Result_14_26_SW0_O,
      O => maccontrol_Mmux_n0023_Result_14_26_SW0_O_GROM
    );
  maccontrol_Mmux_n0023_Result_14_26_SW0_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_14_26_SW0_O_FROM,
      O => maccontrol_Mmux_n0023_Result_14_26_SW0_O
    );
  maccontrol_Mmux_n0023_Result_14_26_SW0_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_14_26_SW0_O_GROM,
      O => maccontrol_Mmux_n0023_Result_14_58_SW0_O
    );
  maccontrol_Mmux_n0023_Result_8_26_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_phydo(8),
      ADR1 => maccontrol_phydi(8),
      ADR2 => maccontrol_n0071,
      ADR3 => maccontrol_n0070,
      O => maccontrol_Mmux_n0023_Result_8_26_SW0_O_FROM
    );
  maccontrol_Mmux_n0023_Result_8_58_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_Mmux_n0023_Result_8_26_2,
      ADR1 => maccontrol_CHOICE1528,
      ADR2 => maccontrol_CHOICE1525,
      ADR3 => maccontrol_Mmux_n0023_Result_8_26_SW0_O,
      O => maccontrol_Mmux_n0023_Result_8_26_SW0_O_GROM
    );
  maccontrol_Mmux_n0023_Result_8_26_SW0_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_8_26_SW0_O_FROM,
      O => maccontrol_Mmux_n0023_Result_8_26_SW0_O
    );
  maccontrol_Mmux_n0023_Result_8_26_SW0_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_8_26_SW0_O_GROM,
      O => maccontrol_Mmux_n0023_Result_8_58_SW0_O
    );
  maccontrol_n00841 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_N30292,
      ADR1 => maccontrol_addr(2),
      ADR2 => maccontrol_addr(3),
      ADR3 => maccontrol_addr(4),
      O => maccontrol_n0084_FROM
    );
  maccontrol_Mmux_n0023_Result_14_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_phystat(14),
      ADR1 => maccontrol_n0067,
      ADR2 => maccontrol_lmacaddr(30),
      ADR3 => maccontrol_n0084,
      O => maccontrol_n0084_GROM
    );
  maccontrol_n0084_XUSED : X_BUF
    port map (
      I => maccontrol_n0084_FROM,
      O => maccontrol_n0084
    );
  maccontrol_n0084_YUSED : X_BUF
    port map (
      I => maccontrol_n0084_GROM,
      O => maccontrol_CHOICE1564
    );
  maccontrol_n00701_1_695 : X_LUT4
    generic map(
      INIT => X"0400"
    )
    port map (
      ADR0 => maccontrol_addr(2),
      ADR1 => maccontrol_addr(3),
      ADR2 => maccontrol_addr(4),
      ADR3 => maccontrol_N30285,
      O => maccontrol_n00701_1_FROM
    );
  maccontrol_Mmux_n0023_Result_31_7 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_phyaddr(31),
      ADR1 => maccontrol_n0069,
      ADR2 => maccontrol_phydi(31),
      ADR3 => maccontrol_n00701_1,
      O => maccontrol_n00701_1_GROM
    );
  maccontrol_n00701_1_XUSED : X_BUF
    port map (
      I => maccontrol_n00701_1_FROM,
      O => maccontrol_n00701_1
    );
  maccontrol_n00701_1_YUSED : X_BUF
    port map (
      I => maccontrol_n00701_1_GROM,
      O => maccontrol_CHOICE1184
    );
  maccontrol_Mmux_n0023_Result_1_26_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_phydi(1),
      ADR1 => maccontrol_phydo(1),
      ADR2 => maccontrol_n0070,
      ADR3 => maccontrol_n0071,
      O => maccontrol_Mmux_n0023_Result_1_26_SW0_O_FROM
    );
  maccontrol_Mmux_n0023_Result_1_58_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_CHOICE1453,
      ADR1 => maccontrol_Mmux_n0023_Result_1_26_2,
      ADR2 => maccontrol_CHOICE1456,
      ADR3 => maccontrol_Mmux_n0023_Result_1_26_SW0_O,
      O => maccontrol_Mmux_n0023_Result_1_26_SW0_O_GROM
    );
  maccontrol_Mmux_n0023_Result_1_26_SW0_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_1_26_SW0_O_FROM,
      O => maccontrol_Mmux_n0023_Result_1_26_SW0_O
    );
  maccontrol_Mmux_n0023_Result_1_26_SW0_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_1_26_SW0_O_GROM,
      O => maccontrol_Mmux_n0023_Result_1_58_SW0_O
    );
  maccontrol_Mmux_n0023_Result_0_11 : X_LUT4
    generic map(
      INIT => X"0200"
    )
    port map (
      ADR0 => maccontrol_lrxucast,
      ADR1 => maccontrol_addr(1),
      ADR2 => maccontrol_addr_0_1,
      ADR3 => maccontrol_N30192,
      O => maccontrol_Mmux_n0023_Result_0_11_O_FROM
    );
  maccontrol_Mmux_n0023_Result_0_19 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => maccontrol_phydo(0),
      ADR1 => maccontrol_CHOICE1429,
      ADR2 => maccontrol_n0071,
      ADR3 => maccontrol_Mmux_n0023_Result_0_11_O,
      O => maccontrol_Mmux_n0023_Result_0_11_O_GROM
    );
  maccontrol_Mmux_n0023_Result_0_11_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_0_11_O_FROM,
      O => maccontrol_Mmux_n0023_Result_0_11_O
    );
  maccontrol_Mmux_n0023_Result_0_11_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_0_11_O_GROM,
      O => maccontrol_CHOICE1433
    );
  maccontrol_Mmux_n0023_Result_3_40_SW0_SW0 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => maccontrol_addr(0),
      ADR1 => VCC,
      ADR2 => maccontrol_lmacaddr(19),
      ADR3 => maccontrol_lmacaddr(35),
      O => maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O_FROM
    );
  maccontrol_Mmux_n0023_Result_3_40_SW0 : X_LUT4
    generic map(
      INIT => X"F808"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(3),
      ADR1 => maccontrol_addr(0),
      ADR2 => maccontrol_addr(1),
      ADR3 => maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O,
      O => maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O_GROM
    );
  maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O_FROM,
      O => maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O
    );
  maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_3_40_SW0_SW0_O_GROM,
      O => maccontrol_N46462
    );
  maccontrol_Ker303091 : X_LUT4
    generic map(
      INIT => X"0005"
    )
    port map (
      ADR0 => maccontrol_bitcnt_88,
      ADR1 => VCC,
      ADR2 => maccontrol_bitcnt_89,
      ADR3 => maccontrol_bitcnt_90,
      O => maccontrol_N30311_FROM
    );
  maccontrol_n001223_SW0 : X_LUT4
    generic map(
      INIT => X"FFDD"
    )
    port map (
      ADR0 => maccontrol_sclkdelta,
      ADR1 => maccontrol_addr(7),
      ADR2 => VCC,
      ADR3 => maccontrol_N30311,
      O => maccontrol_N30311_GROM
    );
  maccontrol_N30311_XUSED : X_BUF
    port map (
      I => maccontrol_N30311_FROM,
      O => maccontrol_N30311
    );
  maccontrol_N30311_YUSED : X_BUF
    port map (
      I => maccontrol_N30311_GROM,
      O => maccontrol_N46628
    );
  maccontrol_Mmux_n0023_Result_4_18 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_N30192,
      ADR1 => maccontrol_lmacaddr(20),
      ADR2 => maccontrol_phydo(4),
      ADR3 => maccontrol_N30212,
      O => maccontrol_Mmux_n0023_Result_4_18_O_FROM
    );
  maccontrol_Mmux_n0023_Result_4_32_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_phystat(4),
      ADR1 => maccontrol_n00671_1,
      ADR2 => maccontrol_N30292,
      ADR3 => maccontrol_Mmux_n0023_Result_4_18_O,
      O => maccontrol_Mmux_n0023_Result_4_18_O_GROM
    );
  maccontrol_Mmux_n0023_Result_4_18_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_4_18_O_FROM,
      O => maccontrol_Mmux_n0023_Result_4_18_O
    );
  maccontrol_Mmux_n0023_Result_4_18_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_4_18_O_GROM,
      O => maccontrol_N46518
    );
  maccontrol_Mmux_n0023_Result_3_6 : X_LUT4
    generic map(
      INIT => X"A800"
    )
    port map (
      ADR0 => maccontrol_addr_1_1,
      ADR1 => maccontrol_phystat(3),
      ADR2 => maccontrol_addr_0_1,
      ADR3 => maccontrol_N30199,
      O => maccontrol_Mmux_n0023_Result_3_6_O_FROM
    );
  maccontrol_Mmux_n0023_Result_3_76_SW0 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => maccontrol_n00691_1,
      ADR1 => maccontrol_phyaddr(3),
      ADR2 => maccontrol_CHOICE1355,
      ADR3 => maccontrol_Mmux_n0023_Result_3_6_O,
      O => maccontrol_Mmux_n0023_Result_3_6_O_GROM
    );
  maccontrol_Mmux_n0023_Result_3_6_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_3_6_O_FROM,
      O => maccontrol_Mmux_n0023_Result_3_6_O
    );
  maccontrol_Mmux_n0023_Result_3_6_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_3_6_O_GROM,
      O => maccontrol_N46555
    );
  maccontrol_Ker301971 : X_LUT4
    generic map(
      INIT => X"0011"
    )
    port map (
      ADR0 => maccontrol_addr(3),
      ADR1 => maccontrol_addr(2),
      ADR2 => VCC,
      ADR3 => maccontrol_addr(4),
      O => maccontrol_N30199_FROM
    );
  maccontrol_Ker301601 : X_LUT4
    generic map(
      INIT => X"A500"
    )
    port map (
      ADR0 => maccontrol_addr(1),
      ADR1 => VCC,
      ADR2 => maccontrol_addr(0),
      ADR3 => maccontrol_N30199,
      O => maccontrol_N30199_GROM
    );
  maccontrol_N30199_XUSED : X_BUF
    port map (
      I => maccontrol_N30199_FROM,
      O => maccontrol_N30199
    );
  maccontrol_N30199_YUSED : X_BUF
    port map (
      I => maccontrol_N30199_GROM,
      O => maccontrol_N30162
    );
  maccontrol_Ker30216_SW0 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_bitcnt_85,
      ADR2 => VCC,
      ADR3 => maccontrol_bitcnt_87,
      O => maccontrol_N42043_FROM
    );
  maccontrol_Ker30216 : X_LUT4
    generic map(
      INIT => X"0004"
    )
    port map (
      ADR0 => maccontrol_bitcnt_89,
      ADR1 => maccontrol_bitcnt_88,
      ADR2 => maccontrol_bitcnt_86,
      ADR3 => maccontrol_N42043,
      O => maccontrol_N42043_GROM
    );
  maccontrol_N42043_XUSED : X_BUF
    port map (
      I => maccontrol_N42043_FROM,
      O => maccontrol_N42043
    );
  maccontrol_N42043_YUSED : X_BUF
    port map (
      I => maccontrol_N42043_GROM,
      O => maccontrol_N30218
    );
  memcontroller_qn_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(1),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_1_IFF_RST,
      O => memcontroller_qn(1)
    );
  MD_1_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_1_IFF_RST
    );
  maccontrol_n00397 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_103,
      ADR1 => maccontrol_phyrstcnt_102,
      ADR2 => maccontrol_phyrstcnt_101,
      ADR3 => maccontrol_phyrstcnt_91,
      O => maccontrol_n00397_O_FROM
    );
  maccontrol_n003910 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_99,
      ADR1 => maccontrol_phyrstcnt_98,
      ADR2 => maccontrol_phyrstcnt_100,
      ADR3 => maccontrol_n00397_O,
      O => maccontrol_n00397_O_GROM
    );
  maccontrol_n00397_O_XUSED : X_BUF
    port map (
      I => maccontrol_n00397_O_FROM,
      O => maccontrol_n00397_O
    );
  maccontrol_n00397_O_YUSED : X_BUF
    port map (
      I => maccontrol_n00397_O_GROM,
      O => maccontrol_CHOICE1582
    );
  maccontrol_Ker301791 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => maccontrol_newcmd,
      ADR1 => RESET_IBUF,
      ADR2 => clkslen,
      ADR3 => maccontrol_addr(7),
      O => maccontrol_N30181_FROM
    );
  maccontrol_n00341 : X_LUT4
    generic map(
      INIT => X"0200"
    )
    port map (
      ADR0 => maccontrol_N30192,
      ADR1 => maccontrol_addr_0_1,
      ADR2 => maccontrol_addr_1_1,
      ADR3 => maccontrol_N30181,
      O => maccontrol_N30181_GROM
    );
  maccontrol_N30181_XUSED : X_BUF
    port map (
      I => maccontrol_N30181_FROM,
      O => maccontrol_N30181
    );
  maccontrol_N30181_YUSED : X_BUF
    port map (
      I => maccontrol_N30181_GROM,
      O => maccontrol_n0034
    );
  maccontrol_n003923 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_92,
      ADR1 => maccontrol_phyrstcnt_109,
      ADR2 => maccontrol_phyrstcnt_110,
      ADR3 => maccontrol_phyrstcnt_108,
      O => maccontrol_n003923_O_FROM
    );
  maccontrol_n003924 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_CHOICE1585,
      ADR2 => VCC,
      ADR3 => maccontrol_n003923_O,
      O => maccontrol_n003923_O_GROM
    );
  maccontrol_n003923_O_XUSED : X_BUF
    port map (
      I => maccontrol_n003923_O_FROM,
      O => maccontrol_n003923_O
    );
  maccontrol_n003923_O_YUSED : X_BUF
    port map (
      I => maccontrol_n003923_O_GROM,
      O => maccontrol_CHOICE1589
    );
  maccontrol_Ker302901 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => maccontrol_addr(0),
      ADR3 => maccontrol_addr(1),
      O => maccontrol_N30292_FROM
    );
  maccontrol_n00711 : X_LUT4
    generic map(
      INIT => X"0200"
    )
    port map (
      ADR0 => maccontrol_addr(3),
      ADR1 => maccontrol_addr(2),
      ADR2 => maccontrol_addr(4),
      ADR3 => maccontrol_N30292,
      O => maccontrol_N30292_GROM
    );
  maccontrol_N30292_XUSED : X_BUF
    port map (
      I => maccontrol_N30292_FROM,
      O => maccontrol_N30292
    );
  maccontrol_N30292_YUSED : X_BUF
    port map (
      I => maccontrol_N30292_GROM,
      O => maccontrol_n0071
    );
  maccontrol_Mmux_n0023_Result_12_18 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_N30192,
      ADR1 => maccontrol_N30212,
      ADR2 => maccontrol_lmacaddr(28),
      ADR3 => maccontrol_phydo(12),
      O => maccontrol_Mmux_n0023_Result_12_18_O_FROM
    );
  maccontrol_Mmux_n0023_Result_12_32_SW0 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_N30292,
      ADR1 => maccontrol_n0067,
      ADR2 => maccontrol_phystat(12),
      ADR3 => maccontrol_Mmux_n0023_Result_12_18_O,
      O => maccontrol_Mmux_n0023_Result_12_18_O_GROM
    );
  maccontrol_Mmux_n0023_Result_12_18_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_12_18_O_FROM,
      O => maccontrol_Mmux_n0023_Result_12_18_O
    );
  maccontrol_Mmux_n0023_Result_12_18_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_12_18_O_GROM,
      O => maccontrol_N46522
    );
  memcontroller_dnout_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_0_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_0_OFF_RST,
      O => memcontroller_dnout(0)
    );
  MD_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_0_OFF_RST
    );
  maccontrol_Ker302971 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_addr(1),
      ADR2 => maccontrol_addr(0),
      ADR3 => VCC,
      O => maccontrol_N30299_FROM
    );
  maccontrol_n00851 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_addr(3),
      ADR1 => maccontrol_addr(4),
      ADR2 => maccontrol_addr(2),
      ADR3 => maccontrol_N30299,
      O => maccontrol_N30299_GROM
    );
  maccontrol_N30299_XUSED : X_BUF
    port map (
      I => maccontrol_N30299_FROM,
      O => maccontrol_N30299
    );
  maccontrol_N30299_YUSED : X_BUF
    port map (
      I => maccontrol_N30299_GROM,
      O => maccontrol_n0085
    );
  maccontrol_n00511 : X_LUT4
    generic map(
      INIT => X"BFBF"
    )
    port map (
      ADR0 => maccontrol_addr(7),
      ADR1 => maccontrol_newcmd,
      ADR2 => maccontrol_n0069,
      ADR3 => VCC,
      O => maccontrol_phyaddr_31_FROM
    );
  maccontrol_PHY_status_n00171 : X_LUT4
    generic map(
      INIT => X"4050"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => maccontrol_PHY_status_cs_FFd1,
      ADR2 => clkslen,
      ADR3 => maccontrol_PHY_status_n00181_O,
      O => maccontrol_phyaddr_31_GROM
    );
  maccontrol_phyaddr_31_XUSED : X_BUF
    port map (
      I => maccontrol_phyaddr_31_FROM,
      O => maccontrol_PHY_status_n00181_O
    );
  maccontrol_phyaddr_31_YUSED : X_BUF
    port map (
      I => maccontrol_phyaddr_31_GROM,
      O => maccontrol_PHY_status_n00171_O
    );
  memtest_Mshreg_dataw4_4_srl_27 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_39,
      A1 => GLOBAL_LOGIC0_29,
      A2 => GLOBAL_LOGIC0_29,
      A3 => GLOBAL_LOGIC0_29,
      D => memtest_dataw1(4),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_4_net55
    );
  memtest_Mshreg_dataw4_5_srl_26 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_20,
      A1 => GLOBAL_LOGIC0_6,
      A2 => GLOBAL_LOGIC0_6,
      A3 => GLOBAL_LOGIC0_10,
      D => memtest_dataw1(5),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_5_net53
    );
  memtest2_Mshreg_data4_11_srl_52 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_34,
      A1 => GLOBAL_LOGIC1_36,
      A2 => GLOBAL_LOGIC0_34,
      A3 => GLOBAL_LOGIC0_34,
      D => memtest2_ldata(11),
      CE => memtest2_n00511_4,
      CLK => clk,
      Q => memtest2_Mshreg_data4_11_net105
    );
  memtest_Mshreg_dataw4_6_srl_25 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_39,
      A1 => GLOBAL_LOGIC0_29,
      A2 => GLOBAL_LOGIC0_29,
      A3 => GLOBAL_LOGIC0_29,
      D => memtest_dataw1(6),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_6_net51
    );
  memtest2_Mshreg_data4_12_srl_51 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_21,
      A1 => GLOBAL_LOGIC1_28,
      A2 => GLOBAL_LOGIC0_15,
      A3 => GLOBAL_LOGIC0_37,
      D => memtest2_ldata(12),
      CE => memtest2_n00511_3,
      CLK => clk,
      Q => memtest2_Mshreg_data4_12_net103
    );
  memtest_Mshreg_dataw4_7_srl_24 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_42,
      A1 => GLOBAL_LOGIC0_3,
      A2 => GLOBAL_LOGIC0_6,
      A3 => GLOBAL_LOGIC0_6,
      D => memtest_dataw1(7),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_7_net49
    );
  memcontroller_ts_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_0_TFF_RST,
      O => memcontroller_ts(0)
    );
  MD_0_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_0_TFF_RST
    );
  memtest_Mshreg_dataw4_8_srl_23 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_39,
      A1 => GLOBAL_LOGIC0_29,
      A2 => GLOBAL_LOGIC0_29,
      A3 => GLOBAL_LOGIC0_29,
      D => memtest_dataw1(8),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_8_net47
    );
  maccontrol_PHY_status_MII_Interface_n001120 : X_LUT4
    generic map(
      INIT => X"1110"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_mdccnt(1),
      ADR1 => maccontrol_PHY_status_MII_Interface_mdccnt(0),
      ADR2 => maccontrol_PHY_status_MII_Interface_cs_FFd3,
      ADR3 => maccontrol_PHY_status_MII_Interface_cs_FFd4,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd3_FROM
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd3_In_696 : X_LUT4
    generic map(
      INIT => X"50DC"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_n0004,
      ADR1 => maccontrol_PHY_status_MII_Interface_cs_FFd4,
      ADR2 => maccontrol_PHY_status_MII_Interface_cs_FFd3,
      ADR3 => maccontrol_PHY_status_MII_Interface_N41734,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd3_In
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd3_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_cs_FFd3_FROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE925
    );
  memtest2_Mshreg_data4_14_srl_49 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_44,
      A1 => GLOBAL_LOGIC1_11,
      A2 => GLOBAL_LOGIC0_46,
      A3 => GLOBAL_LOGIC0_39,
      D => memtest2_ldata(14),
      CE => memtest2_n00511_3,
      CLK => clk,
      Q => memtest2_Mshreg_data4_14_net99
    );
  memtest2_Mshreg_data4_22_srl_41 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_25,
      A1 => GLOBAL_LOGIC1_17,
      A2 => GLOBAL_LOGIC0_25,
      A3 => GLOBAL_LOGIC0_27,
      D => memtest2_ldata(22),
      CE => memtest2_n00511_2,
      CLK => clk,
      Q => memtest2_Mshreg_data4_22_net83
    );
  memtest2_Mshreg_data4_30_srl_33 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_31,
      A1 => GLOBAL_LOGIC1_17,
      A2 => GLOBAL_LOGIC0_31,
      A3 => GLOBAL_LOGIC0_31,
      D => memtest2_ldata(30),
      CE => memtest2_n00511_1,
      CLK => clk,
      Q => memtest2_Mshreg_data4_30_net67
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"F0E0"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd3,
      ADR1 => maccontrol_PHY_status_cs_FFd8,
      ADR2 => maccontrol_PHY_status_MII_Interface_cs_FFd6,
      ADR3 => maccontrol_PHY_status_cs_FFd6,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd5_In
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"EFCC"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_mdccnt(5),
      ADR1 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      ADR2 => MDC_OBUF,
      ADR3 => maccontrol_PHY_status_MII_Interface_cs_FFd4,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd4_In
    );
  memtest_Mshreg_dataw4_9_srl_22 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_38,
      A1 => GLOBAL_LOGIC0_30,
      A2 => GLOBAL_LOGIC0_30,
      A3 => GLOBAL_LOGIC0_30,
      D => memtest_dataw1(9),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_9_net45
    );
  memtest2_Mshreg_data4_15_srl_48 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_39,
      A1 => GLOBAL_LOGIC1_10,
      A2 => GLOBAL_LOGIC0_46,
      A3 => GLOBAL_LOGIC0_44,
      D => memtest2_ldata(15),
      CE => memtest2_n00511_3,
      CLK => clk,
      Q => memtest2_Mshreg_data4_15_net97
    );
  memtest2_Mshreg_data4_23_srl_40 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_25,
      A1 => GLOBAL_LOGIC1_14,
      A2 => GLOBAL_LOGIC0_22,
      A3 => GLOBAL_LOGIC0_25,
      D => memtest2_ldata(23),
      CE => memtest2_n00511_2,
      CLK => clk,
      Q => memtest2_Mshreg_data4_23_net81
    );
  memtest2_Mshreg_data4_31_srl_32 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_40,
      A1 => GLOBAL_LOGIC1_32,
      A2 => GLOBAL_LOGIC0_35,
      A3 => GLOBAL_LOGIC0_35,
      D => memtest2_ldata(31),
      CE => memtest2_n00511_1,
      CLK => clk,
      Q => memtest2_Mshreg_data4_31_net65
    );
  memtest2_Mshreg_data4_16_srl_47 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_45,
      A1 => GLOBAL_LOGIC1_11,
      A2 => GLOBAL_LOGIC0_45,
      A3 => GLOBAL_LOGIC0_27,
      D => memtest2_ldata(16),
      CE => memtest2_n00511_3,
      CLK => clk,
      Q => memtest2_Mshreg_data4_16_net95
    );
  memtest2_Mshreg_data4_17_srl_46 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_25,
      A1 => GLOBAL_LOGIC1_28,
      A2 => GLOBAL_LOGIC0_21,
      A3 => GLOBAL_LOGIC0_25,
      D => memtest2_ldata(17),
      CE => memtest2_n00511_3,
      CLK => clk,
      Q => memtest2_Mshreg_data4_17_net93
    );
  memtest2_Mshreg_data4_25_srl_38 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_45,
      A1 => GLOBAL_LOGIC1_13,
      A2 => GLOBAL_LOGIC0_45,
      A3 => GLOBAL_LOGIC0_45,
      D => memtest2_ldata(25),
      CE => memtest2_n00511_2,
      CLK => clk,
      Q => memtest2_Mshreg_data4_25_net77
    );
  memtest2_Mshreg_data4_18_srl_45 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_31,
      A1 => GLOBAL_LOGIC1_19,
      A2 => GLOBAL_LOGIC0_48,
      A3 => GLOBAL_LOGIC0_31,
      D => memtest2_ldata(18),
      CE => memtest2_n00511_3,
      CLK => clk,
      Q => memtest2_Mshreg_data4_18_net91
    );
  memtest2_Mshreg_data4_26_srl_37 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_45,
      A1 => GLOBAL_LOGIC1_28,
      A2 => GLOBAL_LOGIC0_45,
      A3 => GLOBAL_LOGIC0_45,
      D => memtest2_ldata(26),
      CE => memtest2_n00511_2,
      CLK => clk,
      Q => memtest2_Mshreg_data4_26_net75
    );
  memtest2_Mshreg_data4_19_srl_44 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_31,
      A1 => GLOBAL_LOGIC1_9,
      A2 => GLOBAL_LOGIC0_51,
      A3 => GLOBAL_LOGIC0_31,
      D => memtest2_ldata(19),
      CE => memtest2_n00511_3,
      CLK => clk,
      Q => memtest2_Mshreg_data4_19_net89
    );
  memtest2_Mshreg_data4_27_srl_36 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_41,
      A1 => GLOBAL_LOGIC1_31,
      A2 => GLOBAL_LOGIC0_40,
      A3 => GLOBAL_LOGIC0_40,
      D => memtest2_ldata(27),
      CE => memtest2_n00511_2,
      CLK => clk,
      Q => memtest2_Mshreg_data4_27_net73
    );
  memcontroller_Mmux_dn_inst_mux_f5_181 : X_LUT4
    generic map(
      INIT => X"0E02"
    )
    port map (
      ADR0 => d1(1),
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d2(1),
      O => memcontroller_dn(1)
    );
  memcontroller_Mmux_dn_inst_mux_f5_171 : X_LUT4
    generic map(
      INIT => X"0E02"
    )
    port map (
      ADR0 => d1(0),
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d2(0),
      O => memcontroller_dn(0)
    );
  memcontroller_dnl1_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_1_CEMUXNOT
    );
  memtest2_Mshreg_data4_28_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_28_41_FFY_RST
    );
  memtest2_Mshreg_data4_28_41_697 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_28_net71,
      CE => memtest2_n00511_2,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_28_41_FFY_RST,
      O => memtest2_Mshreg_data4_28_41
    );
  memtest2_Mshreg_data4_28_srl_35 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_21,
      A1 => GLOBAL_LOGIC1_14,
      A2 => GLOBAL_LOGIC0_21,
      A3 => GLOBAL_LOGIC0_21,
      D => memtest2_ldata(28),
      CE => memtest2_n00511_2,
      CLK => clk,
      Q => memtest2_Mshreg_data4_28_net71
    );
  memcontroller_Mmux_dn_inst_mux_f5_201 : X_LUT4
    generic map(
      INIT => X"0B08"
    )
    port map (
      ADR0 => d2(3),
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d1(3),
      O => memcontroller_dn(3)
    );
  memcontroller_Mmux_dn_inst_mux_f5_191 : X_LUT4
    generic map(
      INIT => X"0B08"
    )
    port map (
      ADR0 => d2(2),
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d1(2),
      O => memcontroller_dn(2)
    );
  memcontroller_dnl1_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_3_CEMUXNOT
    );
  memcontroller_dnl1_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_5_FFY_RST
    );
  memcontroller_dnl1_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(4),
      CE => memcontroller_dnl1_5_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_5_FFY_RST,
      O => memcontroller_dnl1(4)
    );
  memcontroller_Mmux_dn_inst_mux_f5_221 : X_LUT4
    generic map(
      INIT => X"4450"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => d2(5),
      ADR2 => d1(5),
      ADR3 => memcontroller_clknum_0_2,
      O => memcontroller_dn(5)
    );
  memcontroller_Mmux_dn_inst_mux_f5_211 : X_LUT4
    generic map(
      INIT => X"5404"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => d1(4),
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => d2(4),
      O => memcontroller_dn(4)
    );
  memcontroller_dnl1_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_5_CEMUXNOT
    );
  memcontroller_dnl1_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_7_FFY_RST
    );
  memcontroller_dnl1_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(6),
      CE => memcontroller_dnl1_7_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_7_FFY_RST,
      O => memcontroller_dnl1(6)
    );
  memcontroller_Mmux_dn_inst_mux_f5_241 : X_LUT4
    generic map(
      INIT => X"3120"
    )
    port map (
      ADR0 => memcontroller_clknum_0_2,
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => d2(7),
      ADR3 => d1(7),
      O => memcontroller_dn(7)
    );
  memcontroller_Mmux_dn_inst_mux_f5_231 : X_LUT4
    generic map(
      INIT => X"00E4"
    )
    port map (
      ADR0 => memcontroller_clknum_0_2,
      ADR1 => d1(6),
      ADR2 => d2(6),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_dn(6)
    );
  memcontroller_dnl1_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_7_CEMUXNOT
    );
  txsim_Mshreg_TX_EN_70 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TX_EN_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => TX_EN_OFF_RST,
      O => txsim_TX_EN_OBUF
    );
  TX_EN_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TX_EN_OFF_RST
    );
  memcontroller_dnl1_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_9_FFY_RST
    );
  memcontroller_dnl1_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(8),
      CE => memcontroller_dnl1_9_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_9_FFY_RST,
      O => memcontroller_dnl1(8)
    );
  memcontroller_Mmux_dn_inst_mux_f5_261 : X_LUT4
    generic map(
      INIT => X"2320"
    )
    port map (
      ADR0 => d2(9),
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => d1(9),
      O => memcontroller_dn(9)
    );
  memcontroller_Mmux_dn_inst_mux_f5_251 : X_LUT4
    generic map(
      INIT => X"3202"
    )
    port map (
      ADR0 => d1(8),
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => d2(8),
      O => memcontroller_dn(8)
    );
  memcontroller_dnl1_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_9_CEMUXNOT
    );
  memcontroller_clknum_1_2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_1_2_FFY_RST
    );
  memcontroller_clknum_1_1_698 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_1_2_GROM,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memcontroller_clknum_1_2_FFY_RST,
      O => memcontroller_clknum_1_1
    );
  memcontroller_clknum_Mmux_n0001_Result_1_1 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_clknum_1_2_GROM
    );
  memcontroller_clknum_1_2_YUSED : X_BUF
    port map (
      I => memcontroller_clknum_1_2_GROM,
      O => memcontroller_clknum_n0001(1)
    );
  memcontroller_dnout_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_1_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_1_OFF_RST,
      O => memcontroller_dnout(1)
    );
  MD_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_1_OFF_RST
    );
  memtest2_Mshreg_data4_29_40_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_29_40_FFY_RST
    );
  memtest2_Mshreg_data4_29_40_699 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_29_net69,
      CE => memtest2_n00511_2,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_29_40_FFY_RST,
      O => memtest2_Mshreg_data4_29_40
    );
  memtest2_Mshreg_data4_29_srl_34 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_45,
      A1 => GLOBAL_LOGIC1_28,
      A2 => GLOBAL_LOGIC0_41,
      A3 => GLOBAL_LOGIC0_41,
      D => memtest2_ldata(29),
      CE => memtest2_n00511_2,
      CLK => clk,
      Q => memtest2_Mshreg_data4_29_net69
    );
  maccontrol_Mshreg_scslll_srl_66 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_0,
      A1 => GLOBAL_LOGIC0_63,
      A2 => GLOBAL_LOGIC0_62,
      A3 => GLOBAL_LOGIC0_62,
      D => SCS_IBUF,
      CE => maccontrol_N30273,
      CLK => clk,
      Q => maccontrol_Mshreg_scslll_net281
    );
  maccontrol_PHY_status_MII_Interface_n0004_2_700 : X_LUT4
    generic map(
      INIT => X"FEFE"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(0),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(1),
      ADR3 => VCC,
      O => maccontrol_PHY_status_MII_Interface_statecnt_0_FROM
    );
  maccontrol_PHY_status_MII_Interface_n0014_0_1 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => VCC,
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(0),
      ADR3 => VCC,
      O => maccontrol_PHY_status_MII_Interface_n0014(0)
    );
  maccontrol_PHY_status_MII_Interface_statecnt_0_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_statecnt_0_FROM,
      O => maccontrol_PHY_status_MII_Interface_n0004_2
    );
  maccontrol_PHY_status_MII_Interface_n0014_3_1 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_n0079,
      ADR1 => maccontrol_PHY_status_MII_Interface_n0078(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => maccontrol_PHY_status_MII_Interface_n0014(3)
    );
  maccontrol_PHY_status_MII_Interface_n0014_2_1 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_n0078(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_n0079,
      O => maccontrol_PHY_status_MII_Interface_n0014(2)
    );
  maccontrol_PHY_status_MII_Interface_n0014_5_1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_MII_Interface_n0078(5),
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_n0079,
      O => maccontrol_PHY_status_MII_Interface_n0014(5)
    );
  maccontrol_PHY_status_MII_Interface_n0014_4_1 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_n0078(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_n0079,
      O => maccontrol_PHY_status_MII_Interface_n0014(4)
    );
  memcontroller_Mmux_dn_inst_mux_f5_281 : X_LUT4
    generic map(
      INIT => X"5404"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => d1(11),
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => d2(11),
      O => memcontroller_dn(11)
    );
  memcontroller_Mmux_dn_inst_mux_f5_271 : X_LUT4
    generic map(
      INIT => X"5044"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => d1(10),
      ADR2 => d2(10),
      ADR3 => memcontroller_clknum_0_2,
      O => memcontroller_dn(10)
    );
  memcontroller_dnl1_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_11_CEMUXNOT
    );
  memcontroller_dnl1_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_21_FFY_RST
    );
  memcontroller_dnl1_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(20),
      CE => memcontroller_dnl1_21_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_21_FFY_RST,
      O => memcontroller_dnl1(20)
    );
  memcontroller_Mmux_dn_inst_mux_f5_381 : X_LUT4
    generic map(
      INIT => X"3120"
    )
    port map (
      ADR0 => memcontroller_clknum_0_2,
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => d2(21),
      ADR3 => d1(21),
      O => memcontroller_dn(21)
    );
  memcontroller_Mmux_dn_inst_mux_f5_371 : X_LUT4
    generic map(
      INIT => X"3202"
    )
    port map (
      ADR0 => d1(20),
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => d2(20),
      O => memcontroller_dn(20)
    );
  memcontroller_dnl1_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_21_CEMUXNOT
    );
  memcontroller_dnl1_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_13_FFY_RST
    );
  memcontroller_dnl1_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(12),
      CE => memcontroller_dnl1_13_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_13_FFY_RST,
      O => memcontroller_dnl1(12)
    );
  memcontroller_Mmux_dn_inst_mux_f5_301 : X_LUT4
    generic map(
      INIT => X"00E4"
    )
    port map (
      ADR0 => memcontroller_clknum_0_2,
      ADR1 => d1(13),
      ADR2 => d2(13),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_dn(13)
    );
  memcontroller_Mmux_dn_inst_mux_f5_291 : X_LUT4
    generic map(
      INIT => X"00D8"
    )
    port map (
      ADR0 => memcontroller_clknum_0_2,
      ADR1 => d2(12),
      ADR2 => d1(12),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_dn(12)
    );
  memcontroller_dnl1_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_13_CEMUXNOT
    );
  memcontroller_ts_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_1_TFF_RST,
      O => memcontroller_ts(1)
    );
  MD_1_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_1_TFF_RST
    );
  memcontroller_dnl1_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_31_FFY_RST
    );
  memcontroller_dnl1_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(30),
      CE => memcontroller_dnl1_31_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_31_FFY_RST,
      O => memcontroller_dnl1(30)
    );
  memcontroller_Mmux_dn_inst_mux_f5_481 : X_LUT4
    generic map(
      INIT => X"2230"
    )
    port map (
      ADR0 => d2(31),
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => d1(31),
      ADR3 => memcontroller_clknum_0_2,
      O => memcontroller_dn(31)
    );
  memcontroller_Mmux_dn_inst_mux_f5_471 : X_LUT4
    generic map(
      INIT => X"00B8"
    )
    port map (
      ADR0 => d2(30),
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => d1(30),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_dn(30)
    );
  memcontroller_dnl1_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_31_CEMUXNOT
    );
  memcontroller_dnl1_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_23_FFY_RST
    );
  memcontroller_dnl1_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(22),
      CE => memcontroller_dnl1_23_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_23_FFY_RST,
      O => memcontroller_dnl1(22)
    );
  memcontroller_Mmux_dn_inst_mux_f5_401 : X_LUT4
    generic map(
      INIT => X"3120"
    )
    port map (
      ADR0 => memcontroller_clknum_0_2,
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => d2(23),
      ADR3 => d1(23),
      O => memcontroller_dn(23)
    );
  memcontroller_Mmux_dn_inst_mux_f5_391 : X_LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => d1(22),
      ADR3 => d2(22),
      O => memcontroller_dn(22)
    );
  memcontroller_dnl1_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_23_CEMUXNOT
    );
  memcontroller_dnl1_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_15_FFY_RST
    );
  memcontroller_dnl1_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(14),
      CE => memcontroller_dnl1_15_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_15_FFY_RST,
      O => memcontroller_dnl1(14)
    );
  memcontroller_Mmux_dn_inst_mux_f5_321 : X_LUT4
    generic map(
      INIT => X"0E04"
    )
    port map (
      ADR0 => memcontroller_clknum_0_2,
      ADR1 => d1(15),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d2(15),
      O => memcontroller_dn(15)
    );
  memcontroller_Mmux_dn_inst_mux_f5_311 : X_LUT4
    generic map(
      INIT => X"0D08"
    )
    port map (
      ADR0 => memcontroller_clknum_0_2,
      ADR1 => d2(14),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d1(14),
      O => memcontroller_dn(14)
    );
  memcontroller_dnl1_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_15_CEMUXNOT
    );
  memcontroller_dnl1_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_25_FFY_RST
    );
  memcontroller_dnl1_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(24),
      CE => memcontroller_dnl1_25_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_25_FFY_RST,
      O => memcontroller_dnl1(24)
    );
  memcontroller_Mmux_dn_inst_mux_f5_421 : X_LUT4
    generic map(
      INIT => X"3202"
    )
    port map (
      ADR0 => d1(25),
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => d2(25),
      O => memcontroller_dn(25)
    );
  memcontroller_Mmux_dn_inst_mux_f5_411 : X_LUT4
    generic map(
      INIT => X"4540"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => d2(24),
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => d1(24),
      O => memcontroller_dn(24)
    );
  memcontroller_dnl1_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_25_CEMUXNOT
    );
  memcontroller_dnl1_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_17_FFY_RST
    );
  memcontroller_dnl1_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(16),
      CE => memcontroller_dnl1_17_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_17_FFY_RST,
      O => memcontroller_dnl1(16)
    );
  memcontroller_Mmux_dn_inst_mux_f5_341 : X_LUT4
    generic map(
      INIT => X"5140"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => d2(17),
      ADR3 => d1(17),
      O => memcontroller_dn(17)
    );
  memcontroller_Mmux_dn_inst_mux_f5_331 : X_LUT4
    generic map(
      INIT => X"00B8"
    )
    port map (
      ADR0 => d2(16),
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => d1(16),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_dn(16)
    );
  memcontroller_dnl1_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_17_CEMUXNOT
    );
  memcontroller_dnl1_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_27_FFY_RST
    );
  memcontroller_dnl1_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(26),
      CE => memcontroller_dnl1_27_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_27_FFY_RST,
      O => memcontroller_dnl1(26)
    );
  memcontroller_Mmux_dn_inst_mux_f5_441 : X_LUT4
    generic map(
      INIT => X"0E02"
    )
    port map (
      ADR0 => d1(27),
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d2(27),
      O => memcontroller_dn(27)
    );
  memcontroller_Mmux_dn_inst_mux_f5_431 : X_LUT4
    generic map(
      INIT => X"0E02"
    )
    port map (
      ADR0 => d1(26),
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d2(26),
      O => memcontroller_dn(26)
    );
  memcontroller_dnl1_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_27_CEMUXNOT
    );
  memcontroller_dnl1_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_19_FFY_RST
    );
  memcontroller_dnl1_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(18),
      CE => memcontroller_dnl1_19_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_19_FFY_RST,
      O => memcontroller_dnl1(18)
    );
  memcontroller_Mmux_dn_inst_mux_f5_361 : X_LUT4
    generic map(
      INIT => X"2320"
    )
    port map (
      ADR0 => d2(19),
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => d1(19),
      O => memcontroller_dn(19)
    );
  memcontroller_Mmux_dn_inst_mux_f5_351 : X_LUT4
    generic map(
      INIT => X"00CA"
    )
    port map (
      ADR0 => d1(18),
      ADR1 => d2(18),
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_dn(18)
    );
  memcontroller_dnl1_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_19_CEMUXNOT
    );
  memcontroller_dnl1_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_29_FFY_RST
    );
  memcontroller_dnl1_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(28),
      CE => memcontroller_dnl1_29_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_29_FFY_RST,
      O => memcontroller_dnl1(28)
    );
  memcontroller_Mmux_dn_inst_mux_f5_461 : X_LUT4
    generic map(
      INIT => X"0C0A"
    )
    port map (
      ADR0 => d1(29),
      ADR1 => d2(29),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => memcontroller_clknum_0_2,
      O => memcontroller_dn(29)
    );
  memcontroller_Mmux_dn_inst_mux_f5_451 : X_LUT4
    generic map(
      INIT => X"2230"
    )
    port map (
      ADR0 => d2(28),
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => d1(28),
      ADR3 => memcontroller_clknum_0_2,
      O => memcontroller_dn(28)
    );
  memcontroller_dnl1_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_29_CEMUXNOT
    );
  memtest2_datalfsr_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_n0214,
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(0)
    );
  memtest2_n02141 : X_LUT4
    generic map(
      INIT => X"9669"
    )
    port map (
      ADR0 => memtest2_datalfsr(31),
      ADR1 => memtest2_datalfsr(0),
      ADR2 => memtest2_datalfsr(1),
      ADR3 => memtest2_datalfsr(21),
      O => memtest2_n0214
    );
  clken_clkcnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => clken_clkcnt_n0000(2),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => clken_n0002,
      O => clken_clkcnt(2)
    );
  clken_n00021 : X_LUT4
    generic map(
      INIT => X"8080"
    )
    port map (
      ADR0 => clken_clkcnt(1),
      ADR1 => clken_clkcnt(2),
      ADR2 => clken_clkcnt(0),
      ADR3 => VCC,
      O => clken_clkcnt_2_FROM
    );
  clken_clkcnt_Madd_n0000_Mxor_Result_2_Result1 : X_LUT4
    generic map(
      INIT => X"3FC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => clken_clkcnt(0),
      ADR2 => clken_clkcnt(1),
      ADR3 => clken_clkcnt(2),
      O => clken_clkcnt_n0000(2)
    );
  clken_clkcnt_2_XUSED : X_BUF
    port map (
      I => clken_clkcnt_2_FROM,
      O => clken_n0002
    );
  maccontrol_PHY_status_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"AAFA"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd3,
      ADR1 => VCC,
      ADR2 => maccontrol_PHY_status_cs_FFd2,
      ADR3 => maccontrol_PHY_status_done,
      O => maccontrol_PHY_status_cs_FFd2_In
    );
  maccontrol_PHY_status_cs_FFd1_In1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_done,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_cs_FFd2,
      O => maccontrol_PHY_status_cs_FFd1_In
    );
  maccontrol_PHY_status_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_done,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_cs_FFd5,
      O => maccontrol_PHY_status_cs_FFd4_In
    );
  maccontrol_PHY_status_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => maccontrol_PHY_status_phyaddrws,
      ADR1 => VCC,
      ADR2 => maccontrol_PHY_status_cs_FFd4,
      ADR3 => VCC,
      O => maccontrol_PHY_status_cs_FFd3_In
    );
  maccontrol_PHY_status_cs_FFd6_In1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_done,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_cs_FFd7,
      O => maccontrol_PHY_status_cs_FFd6_In
    );
  maccontrol_PHY_status_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"CFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_cs_FFd6,
      ADR2 => maccontrol_PHY_status_done,
      ADR3 => maccontrol_PHY_status_cs_FFd5,
      O => maccontrol_PHY_status_cs_FFd5_In
    );
  maccontrol_PHY_status_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"AAEE"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd1,
      ADR1 => maccontrol_PHY_status_cs_FFd4,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_phyaddrws,
      O => maccontrol_PHY_status_cs_FFd8_In
    );
  maccontrol_PHY_status_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"DCDC"
    )
    port map (
      ADR0 => maccontrol_PHY_status_done,
      ADR1 => maccontrol_PHY_status_cs_FFd8,
      ADR2 => maccontrol_PHY_status_cs_FFd7,
      ADR3 => VCC,
      O => maccontrol_PHY_status_cs_FFd7_In
    );
  memtest2_Mshreg_data4_0_srl_63 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_14,
      A1 => GLOBAL_LOGIC1_36,
      A2 => GLOBAL_LOGIC0_14,
      A3 => GLOBAL_LOGIC0_14,
      D => memtest2_ldata(0),
      CE => memtest2_n00511_4,
      CLK => clk,
      Q => memtest2_Mshreg_data4_0_net127
    );
  memtest2_Mshreg_data4_1_srl_62 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_41,
      A1 => GLOBAL_LOGIC1_28,
      A2 => GLOBAL_LOGIC0_21,
      A3 => GLOBAL_LOGIC0_21,
      D => memtest2_ldata(1),
      CE => memtest2_n00511_3,
      CLK => clk,
      Q => memtest2_Mshreg_data4_1_net125
    );
  maccontrol_Mshreg_sinlll_srl_65 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_5,
      A1 => GLOBAL_LOGIC0_55,
      A2 => GLOBAL_LOGIC0_53,
      A3 => GLOBAL_LOGIC0_55,
      D => SIN_IBUF,
      CE => maccontrol_N30273,
      CLK => clk,
      Q => maccontrol_Mshreg_sinlll_net279
    );
  memtest_Mshreg_dataw4_10_srl_21 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_39,
      A1 => GLOBAL_LOGIC0_29,
      A2 => GLOBAL_LOGIC0_29,
      A3 => GLOBAL_LOGIC0_29,
      D => memtest_dataw1(10),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_10_net43
    );
  memtest2_Mshreg_data4_2_srl_61 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_47,
      A1 => GLOBAL_LOGIC1_46,
      A2 => GLOBAL_LOGIC0_20,
      A3 => GLOBAL_LOGIC0_44,
      D => memtest2_ldata(2),
      CE => memtest2_n00511_1,
      CLK => clk,
      Q => memtest2_Mshreg_data4_2_net123
    );
  memtest_Mshreg_dataw4_11_srl_20 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_39,
      A1 => GLOBAL_LOGIC0_29,
      A2 => GLOBAL_LOGIC0_18,
      A3 => GLOBAL_LOGIC0_29,
      D => memtest_dataw1(11),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_11_net41
    );
  memcontroller_qn_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(2),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_2_IFF_RST,
      O => memcontroller_qn(2)
    );
  MD_2_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_2_IFF_RST
    );
  memtest2_Mshreg_data4_3_srl_60 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_46,
      A1 => GLOBAL_LOGIC1_11,
      A2 => GLOBAL_LOGIC0_50,
      A3 => GLOBAL_LOGIC0_46,
      D => memtest2_ldata(3),
      CE => memtest2_n00511_1,
      CLK => clk,
      Q => memtest2_Mshreg_data4_3_net121
    );
  memtest_Mshreg_dataw4_12_srl_19 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_34,
      A1 => GLOBAL_LOGIC0_36,
      A2 => GLOBAL_LOGIC0_36,
      A3 => GLOBAL_LOGIC0_36,
      D => memtest_dataw1(12),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_12_net39
    );
  memtest_Mshreg_dataw4_20_srl_11 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_41,
      A1 => GLOBAL_LOGIC0_16,
      A2 => GLOBAL_LOGIC0_16,
      A3 => GLOBAL_LOGIC0_23,
      D => memtest_dataw1(20),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_20_net23
    );
  memtest2_Mshreg_data4_4_srl_59 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_19,
      A1 => GLOBAL_LOGIC1_15,
      A2 => GLOBAL_LOGIC0_47,
      A3 => GLOBAL_LOGIC0_33,
      D => memtest2_ldata(4),
      CE => memtest2_n00511_1,
      CLK => clk,
      Q => memtest2_Mshreg_data4_4_net119
    );
  memtest_Mshreg_dataw4_13_srl_18 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_23,
      A1 => GLOBAL_LOGIC0_2,
      A2 => GLOBAL_LOGIC0_2,
      A3 => GLOBAL_LOGIC0_2,
      D => memtest_dataw1(13),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_13_net37
    );
  memtest_Mshreg_dataw4_21_srl_10 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_26,
      A1 => GLOBAL_LOGIC0_2,
      A2 => GLOBAL_LOGIC0_2,
      A3 => GLOBAL_LOGIC0_2,
      D => memtest_dataw1(21),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_21_net21
    );
  memtest2_Mshreg_data4_5_srl_58 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_39,
      A1 => GLOBAL_LOGIC1_33,
      A2 => GLOBAL_LOGIC0_39,
      A3 => GLOBAL_LOGIC0_19,
      D => memtest2_ldata(5),
      CE => memtest2_n00511_1,
      CLK => clk,
      Q => memtest2_Mshreg_data4_5_net117
    );
  testrx_n00081 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => testrx_cs_FFd2,
      ADR3 => testrx_cs_FFd3,
      O => testrx_cs_FFd2_FROM
    );
  testrx_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"F020"
    )
    port map (
      ADR0 => testrx_cs_FFd2,
      ADR1 => testrx_n0004,
      ADR2 => testrx_rx_dvl,
      ADR3 => testrx_cs_FFd3,
      O => testrx_cs_FFd2_In
    );
  testrx_cs_FFd2_XUSED : X_BUF
    port map (
      I => testrx_cs_FFd2_FROM,
      O => testrx_n0008
    );
  memtest_Mshreg_dataw4_14_srl_17 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_21,
      A1 => GLOBAL_LOGIC0_9,
      A2 => GLOBAL_LOGIC0_5,
      A3 => GLOBAL_LOGIC0_9,
      D => memtest_dataw1(14),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_14_net35
    );
  memtest_Mshreg_dataw4_22_srl_9 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_41,
      A1 => GLOBAL_LOGIC0_16,
      A2 => GLOBAL_LOGIC0_16,
      A3 => GLOBAL_LOGIC0_16,
      D => memtest_dataw1(22),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_22_net19
    );
  testrx_cs_FFd1_In_SW0 : X_LUT4
    generic map(
      INIT => X"BBBB"
    )
    port map (
      ADR0 => testrx_nextfl,
      ADR1 => testrx_cs_FFd1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => testrx_cs_FFd3_FROM
    );
  testrx_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"B3A0"
    )
    port map (
      ADR0 => testrx_nextfl,
      ADR1 => testrx_rx_dvl,
      ADR2 => testrx_cs_FFd1,
      ADR3 => testrx_cs_FFd3,
      O => testrx_cs_FFd3_In
    );
  testrx_cs_FFd3_XUSED : X_BUF
    port map (
      I => testrx_cs_FFd3_FROM,
      O => testrx_N41780
    );
  memtest2_Mshreg_data4_6_srl_57 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_33,
      A1 => GLOBAL_LOGIC1_12,
      A2 => GLOBAL_LOGIC0_19,
      A3 => GLOBAL_LOGIC0_19,
      D => memtest2_ldata(6),
      CE => memtest2_n00511_1,
      CLK => clk,
      Q => memtest2_Mshreg_data4_6_net115
    );
  memtest_Mshreg_dataw4_15_srl_16 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_44,
      A1 => GLOBAL_LOGIC0_42,
      A2 => GLOBAL_LOGIC0_2,
      A3 => GLOBAL_LOGIC0_2,
      D => memtest_dataw1(15),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_15_net33
    );
  memtest_Mshreg_dataw4_23_srl_8 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_26,
      A1 => GLOBAL_LOGIC0_0,
      A2 => GLOBAL_LOGIC0_0,
      A3 => GLOBAL_LOGIC0_1,
      D => memtest_dataw1(23),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_23_net17
    );
  memtest2_Mshreg_data4_7_srl_56 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_19,
      A1 => GLOBAL_LOGIC1_33,
      A2 => GLOBAL_LOGIC0_13,
      A3 => GLOBAL_LOGIC0_19,
      D => memtest2_ldata(7),
      CE => memtest2_n00511_1,
      CLK => clk,
      Q => memtest2_Mshreg_data4_7_net113
    );
  txsim_Mshreg_TX_EN_net129_LOGIC_ONE_701 : X_ONE
    port map (
      O => txsim_Mshreg_TX_EN_net129_LOGIC_ONE
    );
  txsim_Mshreg_TX_EN_srl_64 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_7,
      A1 => GLOBAL_LOGIC0_56,
      A2 => GLOBAL_LOGIC0_56,
      A3 => GLOBAL_LOGIC0_56,
      D => txsim_llltx,
      CE => txsim_Mshreg_TX_EN_net129_LOGIC_ONE,
      CLK => clk,
      Q => txsim_Mshreg_TX_EN_net129_GSHIFT
    );
  txsim_Mshreg_TX_EN_net129_YUSED : X_BUF
    port map (
      I => txsim_Mshreg_TX_EN_net129_GSHIFT,
      O => txsim_Mshreg_TX_EN_net129
    );
  memtest2_n002184_SW0_2_702 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cnt(9),
      ADR2 => memtest2_cnt(16),
      ADR3 => memtest2_cnt(0),
      O => memtest2_n002184_SW0_2_GROM
    );
  memtest2_n002184_SW0_2_YUSED : X_BUF
    port map (
      I => memtest2_n002184_SW0_2_GROM,
      O => memtest2_n002184_SW0_2
    );
  memcontroller_addr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_12_OD,
      CE => MA_12_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_12_OFF_RST,
      O => memcontroller_ADDREXT(12)
    );
  MA_12_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_12_OFF_RST
    );
  maccontrol_din_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_13_FFY_RST
    );
  maccontrol_din_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(11),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_13_FFY_RST,
      O => maccontrol_din(12)
    );
  maccontrol_n00221 : X_LUT4
    generic map(
      INIT => X"00C8"
    )
    port map (
      ADR0 => maccontrol_sclkdelta,
      ADR1 => clkslen,
      ADR2 => maccontrol_Mshreg_scslll_84,
      ADR3 => RESET_IBUF,
      O => maccontrol_n0022_FROM
    );
  maccontrol_PHY_status_n0019_703 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => clkslen,
      ADR1 => maccontrol_PHY_status_cs_FFd3,
      ADR2 => maccontrol_PHY_status_N23520,
      ADR3 => maccontrol_PHY_status_N42089,
      O => maccontrol_n0022_GROM
    );
  maccontrol_n0022_XUSED : X_BUF
    port map (
      I => maccontrol_n0022_FROM,
      O => maccontrol_n0022
    );
  maccontrol_n0022_YUSED : X_BUF
    port map (
      I => maccontrol_n0022_GROM,
      O => maccontrol_PHY_status_n0019
    );
  memcontroller_addr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_13_OD,
      CE => MA_13_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_13_OFF_RST,
      O => memcontroller_ADDREXT(13)
    );
  MA_13_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_13_OFF_RST
    );
  memtest2_addrlfsr_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(11),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(12)
    );
  memcontroller_oel_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_oel_CEMUXNOT
    );
  memcontroller_oel_BYMUX : X_INV
    port map (
      I => memcontroller_oe,
      O => memcontroller_oel_BYMUXNOT
    );
  maccontrol_Ker303141_1_704 : X_LUT4
    generic map(
      INIT => X"0010"
    )
    port map (
      ADR0 => maccontrol_N46368,
      ADR1 => maccontrol_N42043,
      ADR2 => maccontrol_bitcnt_88,
      ADR3 => maccontrol_bitcnt_89,
      O => maccontrol_Ker303141_1_FROM
    );
  maccontrol_phyrstcnt_inst_lut3_1231 : X_LUT4
    generic map(
      INIT => X"8F0F"
    )
    port map (
      ADR0 => maccontrol_N30199,
      ADR1 => maccontrol_N46337,
      ADR2 => maccontrol_phyrstcnt_91,
      ADR3 => maccontrol_Ker303141_1,
      O => maccontrol_Ker303141_1_GROM
    );
  maccontrol_Ker303141_1_XUSED : X_BUF
    port map (
      I => maccontrol_Ker303141_1_FROM,
      O => maccontrol_Ker303141_1
    );
  maccontrol_Ker303141_1_YUSED : X_BUF
    port map (
      I => maccontrol_Ker303141_1_GROM,
      O => maccontrol_phyrstcnt_inst_lut3_1231_O
    );
  memtest2_deq_0_rt_705 : X_XOR2
    port map (
      I0 => memtest2_deql_0_CYINIT,
      I1 => memtest2_deql_0_FROM,
      O => memtest2_deq_0_rt
    );
  memtest2_deql_0_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_deql_0_FROM
    );
  memtest2_deql_0_CYINIT_706 : X_BUF
    port map (
      I => memtest2_deq(0),
      O => memtest2_deql_0_CYINIT
    );
  txsim_SF2275667_SW0 : X_LUT4
    generic map(
      INIT => X"FFF3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => txsim_counter(2),
      ADR2 => txsim_counter(4),
      ADR3 => txsim_counter(9),
      O => txsim_N46398_GROM
    );
  txsim_N46398_YUSED : X_BUF
    port map (
      I => txsim_N46398_GROM,
      O => txsim_N46398
    );
  memtest2_deq_2_rt_707 : X_XOR2
    port map (
      I0 => memtest2_deql_2_CYINIT,
      I1 => memtest2_deql_2_FROM,
      O => memtest2_deq_2_rt
    );
  memtest2_deql_2_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memtest2_deql_2_FROM
    );
  memtest2_deql_2_CYINIT_708 : X_BUF
    port map (
      I => memtest2_deq(2),
      O => memtest2_deql_2_CYINIT
    );
  maccontrol_PHY_status_cs_Out51 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_cs_FFd6,
      ADR2 => maccontrol_PHY_status_cs_FFd8,
      ADR3 => maccontrol_PHY_status_cs_FFd3,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd6_FROM
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd6_In1 : X_LUT4
    generic map(
      INIT => X"F0FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_MII_Interface_cs_FFd6,
      ADR2 => maccontrol_PHY_status_done,
      ADR3 => maccontrol_PHY_status_start,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd6_In
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd6_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_cs_FFd6_FROM,
      O => maccontrol_PHY_status_start
    );
  maccontrol_Mmux_n0023_Result_11_40_SW0 : X_LUT4
    generic map(
      INIT => X"EA40"
    )
    port map (
      ADR0 => maccontrol_addr(1),
      ADR1 => maccontrol_lmacaddr(11),
      ADR2 => maccontrol_addr(0),
      ADR3 => maccontrol_N46685,
      O => maccontrol_Mmux_n0023_Result_11_40_SW0_O_FROM
    );
  maccontrol_Mmux_n0023_Result_11_40 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_N30192,
      ADR1 => maccontrol_N30212,
      ADR2 => maccontrol_CHOICE1389,
      ADR3 => maccontrol_Mmux_n0023_Result_11_40_SW0_O,
      O => maccontrol_Mmux_n0023_Result_11_40_SW0_O_GROM
    );
  maccontrol_Mmux_n0023_Result_11_40_SW0_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_11_40_SW0_O_FROM,
      O => maccontrol_Mmux_n0023_Result_11_40_SW0_O
    );
  maccontrol_Mmux_n0023_Result_11_40_SW0_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_11_40_SW0_O_GROM,
      O => maccontrol_CHOICE1397
    );
  memtest_Mshreg_dataw4_16_srl_15 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_26,
      A1 => GLOBAL_LOGIC0_17,
      A2 => GLOBAL_LOGIC0_17,
      A3 => GLOBAL_LOGIC0_17,
      D => memtest_dataw1(16),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_16_net31
    );
  memcontroller_qn_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(3),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_3_IFF_RST,
      O => memcontroller_qn(3)
    );
  MD_3_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_3_IFF_RST
    );
  memtest_Mshreg_dataw4_24_srl_7 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_22,
      A1 => GLOBAL_LOGIC0_8,
      A2 => GLOBAL_LOGIC0_4,
      A3 => GLOBAL_LOGIC0_43,
      D => memtest_dataw1(24),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_24_net15
    );
  memtest2_Mshreg_data4_8_srl_55 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_46,
      A1 => GLOBAL_LOGIC1_27,
      A2 => GLOBAL_LOGIC0_46,
      A3 => GLOBAL_LOGIC0_46,
      D => memtest2_ldata(8),
      CE => memtest2_n00511_1,
      CLK => clk,
      Q => memtest2_Mshreg_data4_8_net111
    );
  memtest_Mshreg_dataw4_17_srl_14 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_26,
      A1 => GLOBAL_LOGIC0_1,
      A2 => GLOBAL_LOGIC0_1,
      A3 => GLOBAL_LOGIC0_1,
      D => memtest_dataw1(17),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_17_net29
    );
  memcontroller_dnout_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_2_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_2_OFF_RST,
      O => memcontroller_dnout(2)
    );
  MD_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_2_OFF_RST
    );
  memtest_Mshreg_dataw4_25_srl_6 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_24,
      A1 => GLOBAL_LOGIC0_1,
      A2 => GLOBAL_LOGIC0_1,
      A3 => GLOBAL_LOGIC0_1,
      D => memtest_dataw1(25),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_25_net13
    );
  memtest2_Mshreg_data4_9_srl_54 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_14,
      A1 => GLOBAL_LOGIC1_35,
      A2 => GLOBAL_LOGIC0_34,
      A3 => GLOBAL_LOGIC0_34,
      D => memtest2_ldata(9),
      CE => memtest2_n00511_1,
      CLK => clk,
      Q => memtest2_Mshreg_data4_9_net109
    );
  memtest_Mshreg_dataw4_26_srl_5 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_25,
      A1 => GLOBAL_LOGIC0_0,
      A2 => GLOBAL_LOGIC0_0,
      A3 => GLOBAL_LOGIC0_0,
      D => memtest_dataw1(26),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_26_net11
    );
  memtest_Mshreg_dataw4_18_srl_13 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_23,
      A1 => GLOBAL_LOGIC0_2,
      A2 => GLOBAL_LOGIC0_2,
      A3 => GLOBAL_LOGIC0_2,
      D => memtest_dataw1(18),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_18_net27
    );
  memtest_Mshreg_dataw4_27_srl_4 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_45,
      A1 => GLOBAL_LOGIC0_0,
      A2 => GLOBAL_LOGIC0_0,
      A3 => GLOBAL_LOGIC0_0,
      D => memtest_dataw1(27),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_27_net9
    );
  memtest_Mshreg_dataw4_19_srl_12 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_24,
      A1 => GLOBAL_LOGIC0_2,
      A2 => GLOBAL_LOGIC0_2,
      A3 => GLOBAL_LOGIC0_2,
      D => memtest_dataw1(19),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_19_net25
    );
  maccontrol_lsclkdelta1 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_sclkl,
      ADR2 => maccontrol_sclkll,
      ADR3 => VCC,
      O => maccontrol_lsclkdelta
    );
  memcontroller_n01161 : X_LUT4
    generic map(
      INIT => X"FF30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mwe2,
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_oe_FROM
    );
  memcontroller_wen1 : X_LUT4
    generic map(
      INIT => X"00BB"
    )
    port map (
      ADR0 => mwe2,
      ADR1 => memcontroller_clknum_0_2,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_wen
    );
  memcontroller_oe_XUSED : X_BUF
    port map (
      I => memcontroller_oe_FROM,
      O => memcontroller_n0116
    );
  memcontroller_ts_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_2_TFF_RST,
      O => memcontroller_ts(2)
    );
  MD_2_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_2_TFF_RST
    );
  memtest_Mshreg_dataw4_30_srl_1 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_40,
      A1 => GLOBAL_LOGIC0_23,
      A2 => GLOBAL_LOGIC0_23,
      A3 => GLOBAL_LOGIC0_28,
      D => memtest_dataw1(30),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_30_net3
    );
  memtest2_n01501 : X_LUT4
    generic map(
      INIT => X"9669"
    )
    port map (
      ADR0 => memtest2_addrlfsr(3),
      ADR1 => memtest2_addrlfsr(15),
      ADR2 => memtest2_addrlfsr(12),
      ADR3 => memtest2_addrlfsr(14),
      O => memtest2_n0150
    );
  memtest_Mshreg_dataw4_31_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_31_6_FFY_RST
    );
  memtest_Mshreg_dataw4_31_6_709 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_31_net1,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_31_6_FFY_RST,
      O => memtest_Mshreg_dataw4_31_6
    );
  memtest_Mshreg_dataw4_31_srl_0 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_25,
      A1 => GLOBAL_LOGIC0,
      A2 => GLOBAL_LOGIC0,
      A3 => GLOBAL_LOGIC0,
      D => memtest_dataw1(31),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_31_net1
    );
  memtest_Mshreg_dataw4_28_srl_3 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_43,
      A1 => GLOBAL_LOGIC0_16,
      A2 => GLOBAL_LOGIC0_12,
      A3 => GLOBAL_LOGIC0_12,
      D => memtest_dataw1(28),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_28_net7
    );
  memtest_Mshreg_dataw4_29_srl_2 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_26,
      A1 => GLOBAL_LOGIC0_0,
      A2 => GLOBAL_LOGIC0_0,
      A3 => GLOBAL_LOGIC0_0,
      D => memtest_dataw1(29),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_29_net5
    );
  memtest_Mshreg_dataw4_0_srl_31 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_38,
      A1 => GLOBAL_LOGIC0_30,
      A2 => GLOBAL_LOGIC0_24,
      A3 => GLOBAL_LOGIC0_24,
      D => memtest_dataw1(0),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_0_net63
    );
  memtest_Mshreg_dataw4_1_srl_30 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_38,
      A1 => GLOBAL_LOGIC0_30,
      A2 => GLOBAL_LOGIC0_30,
      A3 => GLOBAL_LOGIC0_30,
      D => memtest_dataw1(1),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_1_net61
    );
  memtest_Mshreg_dataw4_2_srl_29 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_37,
      A1 => GLOBAL_LOGIC0_32,
      A2 => GLOBAL_LOGIC0_32,
      A3 => GLOBAL_LOGIC0_32,
      D => memtest_dataw1(2),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_2_net59
    );
  memtest_Mshreg_dataw4_3_srl_28 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_20,
      A1 => GLOBAL_LOGIC0_7,
      A2 => GLOBAL_LOGIC0_10,
      A3 => GLOBAL_LOGIC0_10,
      D => memtest_dataw1(3),
      CE => clken4,
      CLK => clk,
      Q => memtest_Mshreg_dataw4_3_net57
    );
  memtest2_datain_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_13_FFY_RST
    );
  memtest2_datain_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(12),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_13_FFY_RST,
      O => memtest2_datain(12)
    );
  memtest2_datain_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_21_FFY_RST
    );
  memtest2_datain_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(20),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_21_FFY_RST,
      O => memtest2_datain(20)
    );
  memtest2_datain_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_15_FFY_RST
    );
  memtest2_datain_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(14),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_15_FFY_RST,
      O => memtest2_datain(14)
    );
  memtest2_datain_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_23_FFY_RST
    );
  memtest2_datain_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(22),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_23_FFY_RST,
      O => memtest2_datain(22)
    );
  memtest2_datain_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_31_FFY_RST
    );
  memtest2_datain_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(31),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_31_FFY_RST,
      O => memtest2_datain(31)
    );
  memtest2_datain_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_25_FFY_RST
    );
  memtest2_datain_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(24),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_25_FFY_RST,
      O => memtest2_datain(24)
    );
  d2_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_11_FFY_RST
    );
  memtest2_MD_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(10),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_11_FFY_RST,
      O => d2(10)
    );
  memtest2_datain_26_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_26_FFY_RST
    );
  memtest2_datain_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(26),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_26_FFY_RST,
      O => memtest2_datain(26)
    );
  memcontroller_qn_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(4),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_4_IFF_RST,
      O => memcontroller_qn(4)
    );
  MD_4_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_4_IFF_RST
    );
  memcontroller_dnout_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_3_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_3_OFF_RST,
      O => memcontroller_dnout(3)
    );
  MD_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_3_OFF_RST
    );
  err_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => err_FFY_RST
    );
  memtest_ERR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_lerr,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => err_FFY_RST,
      O => err
    );
  memcontroller_ts_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_3_TFF_RST,
      O => memcontroller_ts(3)
    );
  MD_3_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_3_TFF_RST
    );
  maccontrol_Mmux_n0023_Result_8_26_2_710 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => maccontrol_phyaddr(8),
      ADR1 => VCC,
      ADR2 => maccontrol_n0069,
      ADR3 => maccontrol_N30162,
      O => maccontrol_Mmux_n0023_Result_8_26_2_FROM
    );
  maccontrol_Mmux_n0023_Result_1_26_2_711 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => maccontrol_n0069,
      ADR1 => VCC,
      ADR2 => maccontrol_phyaddr(1),
      ADR3 => maccontrol_N30162,
      O => maccontrol_Mmux_n0023_Result_8_26_2_GROM
    );
  maccontrol_Mmux_n0023_Result_8_26_2_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_8_26_2_FROM,
      O => maccontrol_Mmux_n0023_Result_8_26_2
    );
  maccontrol_Mmux_n0023_Result_8_26_2_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_8_26_2_GROM,
      O => maccontrol_Mmux_n0023_Result_1_26_2
    );
  maccontrol_PHY_status_MII_Interface_sout273_SW1 : X_LUT4
    generic map(
      INIT => X"BBAB"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_CHOICE784,
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR3 => maccontrol_PHY_status_din(14),
      O => maccontrol_PHY_status_MII_Interface_N46670_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout273 : X_LUT4
    generic map(
      INIT => X"EFE0"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_CHOICE770,
      ADR1 => maccontrol_PHY_status_MII_Interface_N46672,
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(1),
      ADR3 => maccontrol_PHY_status_MII_Interface_N46670,
      O => maccontrol_PHY_status_MII_Interface_N46670_GROM
    );
  maccontrol_PHY_status_MII_Interface_N46670_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_N46670_FROM,
      O => maccontrol_PHY_status_MII_Interface_N46670
    );
  maccontrol_PHY_status_MII_Interface_N46670_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_N46670_GROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE793
    );
  maccontrol_phydo_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_5_FFY_RST
    );
  maccontrol_PHY_status_PHYDOUT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(4),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_5_FFY_RST,
      O => maccontrol_phydo(4)
    );
  MDC_OBUF_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MDC_OBUF_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_mdcint : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt(5),
      CE => maccontrol_PHY_status_MII_Interface_N20226,
      CLK => clk,
      SET => GND,
      RST => MDC_OBUF_FFY_RST,
      O => MDC_OBUF
    );
  addr4_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_1_FFY_RST
    );
  memtest_addrcntll_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(0),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_1_FFY_RST,
      O => addr4(0)
    );
  maccontrol_phydo_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_9_FFY_RST
    );
  maccontrol_PHY_status_PHYDOUT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(8),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_9_FFY_RST,
      O => maccontrol_phydo(8)
    );
  addr4_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_3_FFY_RST
    );
  memtest_addrcntll_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(2),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_3_FFY_RST,
      O => addr4(2)
    );
  addr4_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_7_FFY_RST
    );
  memtest_addrcntll_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(6),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_7_FFY_RST,
      O => addr4(6)
    );
  addr4_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_9_FFY_RST
    );
  memtest_addrcntll_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(8),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_9_FFY_RST,
      O => addr4(8)
    );
  memtest2_ldata_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_1_FFY_RST
    );
  memtest2_ldata_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(0),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_1_FFY_RST,
      O => memtest2_ldata(0)
    );
  memtest2_ldata_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_5_FFY_RST
    );
  memtest2_ldata_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(4),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_5_FFY_RST,
      O => memtest2_ldata(4)
    );
  maccontrol_Mmux_n0023_Result_6_26_2_712 : X_LUT4
    generic map(
      INIT => X"EEAA"
    )
    port map (
      ADR0 => maccontrol_N30162,
      ADR1 => maccontrol_n0069,
      ADR2 => VCC,
      ADR3 => maccontrol_phyaddr(6),
      O => maccontrol_Mmux_n0023_Result_6_26_2_FROM
    );
  maccontrol_Mmux_n0023_Result_2_26_2_713 : X_LUT4
    generic map(
      INIT => X"ECEC"
    )
    port map (
      ADR0 => maccontrol_phyaddr(2),
      ADR1 => maccontrol_N30162,
      ADR2 => maccontrol_n0069,
      ADR3 => VCC,
      O => maccontrol_Mmux_n0023_Result_6_26_2_GROM
    );
  maccontrol_Mmux_n0023_Result_6_26_2_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_6_26_2_FROM,
      O => maccontrol_Mmux_n0023_Result_6_26_2
    );
  maccontrol_Mmux_n0023_Result_6_26_2_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_6_26_2_GROM,
      O => maccontrol_Mmux_n0023_Result_2_26_2
    );
  memcontroller_qn_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(5),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_5_IFF_RST,
      O => memcontroller_qn(5)
    );
  MD_5_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_5_IFF_RST
    );
  memtest2_ldata_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_7_FFY_RST
    );
  memtest2_ldata_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(6),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_7_FFY_RST,
      O => memtest2_ldata(6)
    );
  memcontroller_dnout_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_4_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_4_OFF_RST,
      O => memcontroller_dnout(4)
    );
  MD_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_4_OFF_RST
    );
  q2_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_3_FFY_RST
    );
  memcontroller_Q2_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(2),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_3_FFY_RST,
      O => q2(2)
    );
  memtest2_ldata_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_9_FFY_RST
    );
  memtest2_ldata_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(8),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_9_FFY_RST,
      O => memtest2_ldata(8)
    );
  q2_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_5_FFY_RST
    );
  memcontroller_Q2_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(4),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_5_FFY_RST,
      O => q2(4)
    );
  maccontrol_Ker302831 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_addr(1),
      ADR2 => VCC,
      ADR3 => maccontrol_addr(0),
      O => maccontrol_N30285_FROM
    );
  maccontrol_Ker302261_SW12 : X_LUT4
    generic map(
      INIT => X"0808"
    )
    port map (
      ADR0 => maccontrol_din(0),
      ADR1 => maccontrol_addr(0),
      ADR2 => maccontrol_addr(1),
      ADR3 => VCC,
      O => maccontrol_N30285_GROM
    );
  maccontrol_N30285_XUSED : X_BUF
    port map (
      I => maccontrol_N30285_FROM,
      O => maccontrol_N30285
    );
  maccontrol_N30285_YUSED : X_BUF
    port map (
      I => maccontrol_N30285_GROM,
      O => maccontrol_N46337
    );
  maccontrol_Ker302711 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => clkslen,
      ADR3 => RESET_IBUF,
      O => maccontrol_N30273_FROM
    );
  maccontrol_PHY_status_n00111 : X_LUT4
    generic map(
      INIT => X"0A00"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd4,
      ADR1 => VCC,
      ADR2 => RESET_IBUF,
      ADR3 => clkslen,
      O => maccontrol_N30273_GROM
    );
  maccontrol_N30273_XUSED : X_BUF
    port map (
      I => maccontrol_N30273_FROM,
      O => maccontrol_N30273
    );
  maccontrol_N30273_YUSED : X_BUF
    port map (
      I => maccontrol_N30273_GROM,
      O => maccontrol_PHY_status_n0011
    );
  memcontroller_ts_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_4_TFF_RST,
      O => memcontroller_ts(4)
    );
  MD_4_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_4_TFF_RST
    );
  q4_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_1_FFY_RST
    );
  memcontroller_Q4_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(0),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_1_FFY_RST,
      O => q4(0)
    );
  maccontrol_Mmux_n0023_Result_7_40_SW0 : X_LUT4
    generic map(
      INIT => X"F088"
    )
    port map (
      ADR0 => maccontrol_addr(0),
      ADR1 => maccontrol_lmacaddr(7),
      ADR2 => maccontrol_N46689,
      ADR3 => maccontrol_addr(1),
      O => maccontrol_Mmux_n0023_Result_7_40_SW0_O_FROM
    );
  maccontrol_Mmux_n0023_Result_7_40 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_N30192,
      ADR1 => maccontrol_N30212,
      ADR2 => maccontrol_CHOICE1368,
      ADR3 => maccontrol_Mmux_n0023_Result_7_40_SW0_O,
      O => maccontrol_Mmux_n0023_Result_7_40_SW0_O_GROM
    );
  maccontrol_Mmux_n0023_Result_7_40_SW0_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_7_40_SW0_O_FROM,
      O => maccontrol_Mmux_n0023_Result_7_40_SW0_O
    );
  maccontrol_Mmux_n0023_Result_7_40_SW0_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_7_40_SW0_O_GROM,
      O => maccontrol_CHOICE1376
    );
  maccontrol_Ker302101 : X_LUT4
    generic map(
      INIT => X"000A"
    )
    port map (
      ADR0 => maccontrol_addr(3),
      ADR1 => VCC,
      ADR2 => maccontrol_addr(2),
      ADR3 => maccontrol_addr(4),
      O => maccontrol_N30212_FROM
    );
  maccontrol_Ker302261_SW16 : X_LUT4
    generic map(
      INIT => X"0010"
    )
    port map (
      ADR0 => maccontrol_addr(2),
      ADR1 => maccontrol_addr(3),
      ADR2 => maccontrol_din(0),
      ADR3 => maccontrol_addr(4),
      O => maccontrol_N30212_GROM
    );
  maccontrol_N30212_XUSED : X_BUF
    port map (
      I => maccontrol_N30212_FROM,
      O => maccontrol_N30212
    );
  maccontrol_N30212_YUSED : X_BUF
    port map (
      I => maccontrol_N30212_GROM,
      O => maccontrol_N46356
    );
  maccontrol_PHY_status_n00151_1_714 : X_LUT4
    generic map(
      INIT => X"FF33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => clkslen,
      ADR2 => VCC,
      ADR3 => RESET_IBUF,
      O => maccontrol_PHY_status_n00151_1_FROM
    );
  maccontrol_PHY_status_n00211 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => maccontrol_PHY_status_N23512,
      ADR2 => maccontrol_PHY_status_done,
      ADR3 => clkslen,
      O => maccontrol_PHY_status_n00151_1_GROM
    );
  maccontrol_PHY_status_n00151_1_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_n00151_1_FROM,
      O => maccontrol_PHY_status_n00151_1
    );
  maccontrol_PHY_status_n00151_1_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_n00151_1_GROM,
      O => maccontrol_PHY_status_n0021
    );
  memtest2_Ker226584 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => memtest2_cnt(6),
      ADR1 => memtest2_cnt(3),
      ADR2 => memtest2_cnt(4),
      ADR3 => memtest2_cnt(5),
      O => memtest2_CHOICE1064_GROM
    );
  memtest2_CHOICE1064_YUSED : X_BUF
    port map (
      I => memtest2_CHOICE1064_GROM,
      O => memtest2_CHOICE1064
    );
  memtest2_Ker226589 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => memtest2_cnt(8),
      ADR1 => memtest2_cnt(7),
      ADR2 => memtest2_cs(0),
      ADR3 => memtest2_cnt(9),
      O => memtest2_CHOICE1067_FROM
    );
  memtest2_Ker2265849_2_715 : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_CHOICE1064,
      ADR2 => memtest2_CHOICE1071,
      ADR3 => memtest2_CHOICE1067,
      O => memtest2_CHOICE1067_GROM
    );
  memtest2_CHOICE1067_XUSED : X_BUF
    port map (
      I => memtest2_CHOICE1067_FROM,
      O => memtest2_CHOICE1067
    );
  memtest2_CHOICE1067_YUSED : X_BUF
    port map (
      I => memtest2_CHOICE1067_GROM,
      O => memtest2_Ker2265849_2
    );
  maccontrol_phyaddr_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_2_FFY_RST
    );
  maccontrol_phyaddr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(2),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_2_FFY_RST,
      O => maccontrol_phyaddr(2)
    );
  maccontrol_phyaddr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_5_FFY_RST
    );
  maccontrol_phyaddr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(4),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_5_FFY_RST,
      O => maccontrol_phyaddr(4)
    );
  maccontrol_phyaddr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_7_FFY_RST
    );
  maccontrol_phyaddr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(6),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_7_FFY_RST,
      O => maccontrol_phyaddr(6)
    );
  maccontrol_phyaddr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_9_FFY_RST
    );
  maccontrol_phyaddr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(8),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_9_FFY_RST,
      O => maccontrol_phyaddr(8)
    );
  maccontrol_PHY_status_dout_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_1_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(0),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_1_FFY_RST,
      O => maccontrol_PHY_status_dout(0)
    );
  maccontrol_PHY_status_dout_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_3_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(2),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_3_FFY_RST,
      O => maccontrol_PHY_status_dout(2)
    );
  maccontrol_PHY_status_dout_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_5_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(4),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_5_FFY_RST,
      O => maccontrol_PHY_status_dout(4)
    );
  maccontrol_PHY_status_dout_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_9_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(8),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_9_FFY_RST,
      O => maccontrol_PHY_status_dout(8)
    );
  maccontrol_phydo_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_11_FFY_RST
    );
  maccontrol_PHY_status_PHYDOUT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(10),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_11_FFY_RST,
      O => maccontrol_phydo(10)
    );
  memcontroller_dnout_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_5_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_5_OFF_RST,
      O => memcontroller_dnout(5)
    );
  MD_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_5_OFF_RST
    );
  maccontrol_phydo_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_13_FFY_RST
    );
  maccontrol_PHY_status_PHYDOUT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(12),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_13_FFY_RST,
      O => maccontrol_phydo(12)
    );
  maccontrol_phydo_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_15_FFY_RST
    );
  maccontrol_PHY_status_PHYDOUT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(14),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_15_FFY_RST,
      O => maccontrol_phydo(14)
    );
  addr4_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_11_FFY_RST
    );
  memtest_addrcntll_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(10),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_11_FFY_RST,
      O => addr4(10)
    );
  addr4_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_13_FFY_RST
    );
  memtest_addrcntll_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(12),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_13_FFY_RST,
      O => addr4(12)
    );
  addr4_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_15_FFY_RST
    );
  memtest_addrcntll_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(14),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_15_FFY_RST,
      O => addr4(14)
    );
  maccontrol_Mmux_n0023_Result_10_26_2_716 : X_LUT4
    generic map(
      INIT => X"EECC"
    )
    port map (
      ADR0 => maccontrol_n0069,
      ADR1 => maccontrol_N30162,
      ADR2 => VCC,
      ADR3 => maccontrol_phyaddr(10),
      O => maccontrol_Mmux_n0023_Result_10_26_2_FROM
    );
  maccontrol_Mmux_n0023_Result_5_26_2_717 : X_LUT4
    generic map(
      INIT => X"EAEA"
    )
    port map (
      ADR0 => maccontrol_N30162,
      ADR1 => maccontrol_n0069,
      ADR2 => maccontrol_phyaddr(5),
      ADR3 => VCC,
      O => maccontrol_Mmux_n0023_Result_10_26_2_GROM
    );
  maccontrol_Mmux_n0023_Result_10_26_2_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_10_26_2_FROM,
      O => maccontrol_Mmux_n0023_Result_10_26_2
    );
  maccontrol_Mmux_n0023_Result_10_26_2_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_10_26_2_GROM,
      O => maccontrol_Mmux_n0023_Result_5_26_2
    );
  maccontrol_PHY_status_MII_Interface_n001111 : X_LUT4
    generic map(
      INIT => X"0004"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_mdccnt(3),
      ADR1 => maccontrol_PHY_status_MII_Interface_mdccnt(5),
      ADR2 => maccontrol_PHY_status_MII_Interface_mdccnt(2),
      ADR3 => maccontrol_PHY_status_MII_Interface_mdccnt(4),
      O => maccontrol_PHY_status_MII_Interface_CHOICE920_FROM
    );
  maccontrol_PHY_status_MII_Interface_n001127 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => maccontrol_PHY_status_MII_Interface_CHOICE925,
      ADR2 => clkslen,
      ADR3 => maccontrol_PHY_status_MII_Interface_CHOICE920,
      O => maccontrol_PHY_status_MII_Interface_CHOICE920_GROM
    );
  maccontrol_PHY_status_MII_Interface_CHOICE920_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE920_FROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE920
    );
  maccontrol_PHY_status_MII_Interface_CHOICE920_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE920_GROM,
      O => maccontrol_PHY_status_MII_Interface_n0011
    );
  memcontroller_ts_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_5_TFF_RST,
      O => memcontroller_ts(5)
    );
  MD_5_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_5_TFF_RST
    );
  Q_n0034_2_718 : X_LUT4
    generic map(
      INIT => X"A000"
    )
    port map (
      ADR0 => cnt0(0),
      ADR1 => VCC,
      ADR2 => cnt0(2),
      ADR3 => cnt0(1),
      O => Q_n0034_2_FROM
    );
  Q_n0034_719 : X_LUT4
    generic map(
      INIT => X"7FFF"
    )
    port map (
      ADR0 => cnt0(4),
      ADR1 => Q_n0034_2,
      ADR2 => cnt0(3),
      ADR3 => cnt0(5),
      O => Q_n0034_2_GROM
    );
  Q_n0034_2_XUSED : X_BUF
    port map (
      I => Q_n0034_2_FROM,
      O => Q_n0034_2
    );
  Q_n0034_2_YUSED : X_BUF
    port map (
      I => Q_n0034_2_GROM,
      O => Q_n0034
    );
  memtest2_datalfsr_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(11),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(12)
    );
  memtest2_datalfsr_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(13),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(14)
    );
  memtest2_datalfsr_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(21),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(22)
    );
  memtest2_datalfsr_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(29),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(30)
    );
  memtest2_datalfsr_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(15),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(16)
    );
  memtest2_datalfsr_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(23),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(24)
    );
  memcontroller_qn_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(6),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_6_IFF_RST,
      O => memcontroller_qn(6)
    );
  MD_6_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_6_IFF_RST
    );
  memcontroller_dnl2_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_1_FFY_RST
    );
  memcontroller_dnl2_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(0),
      CE => memcontroller_dnl2_1_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_1_FFY_RST,
      O => memcontroller_dnl2(0)
    );
  memcontroller_dnl2_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_1_CEMUXNOT
    );
  maccontrol_lmacaddr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_11_FFY_RST
    );
  maccontrol_lmacaddr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(10),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_11_FFY_RST,
      O => maccontrol_lmacaddr(10)
    );
  memcontroller_dnl2_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_3_FFY_RST
    );
  memcontroller_dnl2_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(2),
      CE => memcontroller_dnl2_3_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_3_FFY_RST,
      O => memcontroller_dnl2(2)
    );
  memcontroller_dnl2_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_3_CEMUXNOT
    );
  maccontrol_lmacaddr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_13_FFY_RST
    );
  maccontrol_lmacaddr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(12),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_13_FFY_RST,
      O => maccontrol_lmacaddr(12)
    );
  memcontroller_dnl2_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_5_FFY_RST
    );
  memcontroller_dnl2_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(4),
      CE => memcontroller_dnl2_5_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_5_FFY_RST,
      O => memcontroller_dnl2(4)
    );
  memcontroller_dnl2_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_5_CEMUXNOT
    );
  maccontrol_lmacaddr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_15_FFY_RST
    );
  maccontrol_lmacaddr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(14),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_15_FFY_RST,
      O => maccontrol_lmacaddr(14)
    );
  memtest2_ldata_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_11_FFY_RST
    );
  memtest2_ldata_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(10),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_11_FFY_RST,
      O => memtest2_ldata(10)
    );
  memcontroller_dnl2_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_7_CEMUXNOT
    );
  memcontroller_dnout_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_6_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_6_OFF_RST,
      O => memcontroller_dnout(6)
    );
  MD_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_6_OFF_RST
    );
  maccontrol_lmacaddr_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_41_FFY_RST
    );
  maccontrol_lmacaddr_40 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(8),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_41_FFY_RST,
      O => maccontrol_lmacaddr(40)
    );
  maccontrol_lmacaddr_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_17_FFY_RST
    );
  maccontrol_lmacaddr_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(0),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_17_FFY_RST,
      O => maccontrol_lmacaddr(16)
    );
  maccontrol_lmacaddr_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_25_FFY_RST
    );
  maccontrol_lmacaddr_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(8),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_25_FFY_RST,
      O => maccontrol_lmacaddr(24)
    );
  memcontroller_clknum_0_2_BXMUX : X_INV
    port map (
      I => memcontroller_clknum_0_2,
      O => memcontroller_clknum_0_2_BXMUXNOT
    );
  memcontroller_clknum_0_2_BYMUX : X_INV
    port map (
      I => memcontroller_clknum_0_2,
      O => memcontroller_clknum_0_2_BYMUXNOT
    );
  memcontroller_dnl2_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_9_CEMUXNOT
    );
  memcontroller_ts_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_6_TFF_RST,
      O => memcontroller_ts(6)
    );
  MD_6_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_6_TFF_RST
    );
  maccontrol_lmacaddr_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_19_FFY_RST
    );
  maccontrol_lmacaddr_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(2),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_19_FFY_RST,
      O => maccontrol_lmacaddr(18)
    );
  memtest2_ldata_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_31_FFY_RST
    );
  memtest2_ldata_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(30),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_31_FFY_RST,
      O => memtest2_ldata(30)
    );
  memcontroller_qn_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(7),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_7_IFF_RST,
      O => memcontroller_qn(7)
    );
  MD_7_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_7_IFF_RST
    );
  maccontrol_lmacaddr_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_29_FFY_RST
    );
  maccontrol_lmacaddr_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(12),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_29_FFY_RST,
      O => maccontrol_lmacaddr(28)
    );
  maccontrol_lmacaddr_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_47_FFY_RST
    );
  maccontrol_lmacaddr_46 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(14),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_47_FFY_RST,
      O => maccontrol_lmacaddr(46)
    );
  memtest2_ldata_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_27_FFY_RST
    );
  memtest2_ldata_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(26),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_27_FFY_RST,
      O => memtest2_ldata(26)
    );
  memcontroller_qn_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(8),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_8_IFF_RST,
      O => memcontroller_qn(8)
    );
  MD_8_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_8_IFF_RST
    );
  memcontroller_dnout_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_7_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_7_OFF_RST,
      O => memcontroller_dnout(7)
    );
  MD_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_7_OFF_RST
    );
  memtest2_n002184_2_720 : X_LUT4
    generic map(
      INIT => X"8800"
    )
    port map (
      ADR0 => memtest2_CHOICE941,
      ADR1 => memtest2_Mcompar_n0028_inst_lut4_16,
      ADR2 => VCC,
      ADR3 => memtest2_CHOICE948,
      O => memtest2_lfsr_rst_FROM
    );
  memtest2_n002184 : X_LUT4
    generic map(
      INIT => X"0100"
    )
    port map (
      ADR0 => memtest2_n002184_SW0_2,
      ADR1 => memtest2_cnt(7),
      ADR2 => memtest2_cnt(8),
      ADR3 => memtest2_n002184_2,
      O => memtest2_n0021
    );
  memtest2_lfsr_rst_XUSED : X_BUF
    port map (
      I => memtest2_lfsr_rst_FROM,
      O => memtest2_n002184_2
    );
  memcontroller_ts_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_7_TFF_RST,
      O => memcontroller_ts(7)
    );
  MD_7_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_7_TFF_RST
    );
  testrx_n00044 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => testrx_addr(0),
      ADR1 => testrx_addr(2),
      ADR2 => testrx_addr(3),
      ADR3 => testrx_addr(1),
      O => testrx_CHOICE930_GROM
    );
  testrx_CHOICE930_YUSED : X_BUF
    port map (
      I => testrx_CHOICE930_GROM,
      O => testrx_CHOICE930
    );
  maccontrol_PHY_status_MII_Interface_sout12 : X_LUT4
    generic map(
      INIT => X"A088"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      ADR1 => maccontrol_PHY_status_din(11),
      ADR2 => maccontrol_PHY_status_din(3),
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      O => maccontrol_PHY_status_MII_Interface_CHOICE735_FROM
    );
  maccontrol_PHY_status_MII_Interface_sts28_SW0 : X_LUT4
    generic map(
      INIT => X"3FFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(1),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      O => maccontrol_PHY_status_MII_Interface_CHOICE735_GROM
    );
  maccontrol_PHY_status_MII_Interface_CHOICE735_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE735_FROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE735
    );
  maccontrol_PHY_status_MII_Interface_CHOICE735_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE735_GROM,
      O => maccontrol_PHY_status_MII_Interface_N46530
    );
  testrx_n00049 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => testrx_addr(4),
      ADR1 => testrx_addr(7),
      ADR2 => testrx_addr(5),
      ADR3 => testrx_addr(6),
      O => testrx_CHOICE933_GROM
    );
  testrx_CHOICE933_YUSED : X_BUF
    port map (
      I => testrx_CHOICE933_GROM,
      O => testrx_CHOICE933
    );
  maccontrol_Mmux_n0023_Result_23_7 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n00701_1,
      ADR1 => maccontrol_phyaddr(23),
      ADR2 => maccontrol_phydi(23),
      ADR3 => maccontrol_n0069,
      O => maccontrol_CHOICE1204_FROM
    );
  maccontrol_Mmux_n0023_Result_0_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_phydi(0),
      ADR1 => maccontrol_n00701_1,
      ADR2 => maccontrol_n0069,
      ADR3 => maccontrol_phyaddr(0),
      O => maccontrol_CHOICE1204_GROM
    );
  maccontrol_CHOICE1204_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1204_FROM,
      O => maccontrol_CHOICE1204
    );
  maccontrol_CHOICE1204_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1204_GROM,
      O => maccontrol_CHOICE1426
    );
  maccontrol_Mmux_n0023_Result_10_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(42),
      ADR1 => maccontrol_n0085,
      ADR2 => maccontrol_n0083,
      ADR3 => maccontrol_lmacaddr(10),
      O => maccontrol_CHOICE1543_FROM
    );
  maccontrol_Mmux_n0023_Result_1_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(33),
      ADR1 => maccontrol_n0083,
      ADR2 => maccontrol_lmacaddr(1),
      ADR3 => maccontrol_n0085,
      O => maccontrol_CHOICE1543_GROM
    );
  maccontrol_CHOICE1543_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1543_FROM,
      O => maccontrol_CHOICE1543
    );
  maccontrol_CHOICE1543_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1543_GROM,
      O => maccontrol_CHOICE1453
    );
  maccontrol_n00321 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => maccontrol_N30181,
      ADR1 => maccontrol_N30206,
      ADR2 => maccontrol_addr_0_1,
      ADR3 => maccontrol_addr_1_1,
      O => maccontrol_n0032_FROM
    );
  maccontrol_Mmux_n0023_Result_0_8 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_addr_0_1,
      ADR1 => maccontrol_N30206,
      ADR2 => maccontrol_addr(1),
      ADR3 => maccontrol_lrxmcast,
      O => maccontrol_n0032_GROM
    );
  maccontrol_n0032_XUSED : X_BUF
    port map (
      I => maccontrol_n0032_FROM,
      O => maccontrol_n0032
    );
  maccontrol_n0032_YUSED : X_BUF
    port map (
      I => maccontrol_n0032_GROM,
      O => maccontrol_CHOICE1429
    );
  maccontrol_Mmux_n0023_Result_6_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_n0085,
      ADR1 => maccontrol_n0083,
      ADR2 => maccontrol_lmacaddr(6),
      ADR3 => maccontrol_lmacaddr(38),
      O => maccontrol_CHOICE1489_FROM
    );
  maccontrol_Mmux_n0023_Result_2_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n0085,
      ADR1 => maccontrol_lmacaddr(2),
      ADR2 => maccontrol_lmacaddr(34),
      ADR3 => maccontrol_n0083,
      O => maccontrol_CHOICE1489_GROM
    );
  maccontrol_CHOICE1489_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1489_FROM,
      O => maccontrol_CHOICE1489
    );
  maccontrol_CHOICE1489_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1489_GROM,
      O => maccontrol_CHOICE1471
    );
  maccontrol_Mmux_n0023_Result_10_9 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_n0084,
      ADR1 => maccontrol_n0067,
      ADR2 => maccontrol_phystat(10),
      ADR3 => maccontrol_lmacaddr(26),
      O => maccontrol_CHOICE1546_FROM
    );
  maccontrol_Mmux_n0023_Result_1_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(17),
      ADR1 => maccontrol_n0084,
      ADR2 => maccontrol_n0067,
      ADR3 => maccontrol_phystat(1),
      O => maccontrol_CHOICE1546_GROM
    );
  maccontrol_CHOICE1546_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1546_FROM,
      O => maccontrol_CHOICE1546
    );
  maccontrol_CHOICE1546_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1546_GROM,
      O => maccontrol_CHOICE1456
    );
  maccontrol_Mmux_n0023_Result_0_43_SW0 : X_LUT4
    generic map(
      INIT => X"B5BF"
    )
    port map (
      ADR0 => maccontrol_addr(0),
      ADR1 => maccontrol_lrxbcast,
      ADR2 => maccontrol_addr(1),
      ADR3 => maccontrol_lrxallf,
      O => maccontrol_N46676_FROM
    );
  maccontrol_Mmux_n0023_Result_0_43 : X_LUT4
    generic map(
      INIT => X"0020"
    )
    port map (
      ADR0 => maccontrol_addr(3),
      ADR1 => maccontrol_addr(2),
      ADR2 => maccontrol_addr(4),
      ADR3 => maccontrol_N46676,
      O => maccontrol_N46676_GROM
    );
  maccontrol_N46676_XUSED : X_BUF
    port map (
      I => maccontrol_N46676_FROM,
      O => maccontrol_N46676
    );
  maccontrol_N46676_YUSED : X_BUF
    port map (
      I => maccontrol_N46676_GROM,
      O => maccontrol_CHOICE1439
    );
  maccontrol_Mmux_n0023_Result_8_9 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_phystat(8),
      ADR1 => maccontrol_lmacaddr(24),
      ADR2 => maccontrol_n00671_1,
      ADR3 => maccontrol_n0084,
      O => maccontrol_CHOICE1528_FROM
    );
  maccontrol_Mmux_n0023_Result_5_9 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n0084,
      ADR1 => maccontrol_n00671_1,
      ADR2 => maccontrol_lmacaddr(21),
      ADR3 => maccontrol_phystat(5),
      O => maccontrol_CHOICE1528_GROM
    );
  maccontrol_CHOICE1528_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1528_FROM,
      O => maccontrol_CHOICE1528
    );
  maccontrol_CHOICE1528_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1528_GROM,
      O => maccontrol_CHOICE1510
    );
  memtest2_n002125 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(12),
      ADR1 => memtest2_cnt(11),
      ADR2 => memtest2_cnt(13),
      ADR3 => memtest2_cnt(2),
      O => memtest2_CHOICE948_FROM
    );
  memtest2_Ker2265821 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => memtest2_cnt(10),
      ADR1 => memtest2_cnt(11),
      ADR2 => memtest2_cnt(12),
      ADR3 => memtest2_cnt(13),
      O => memtest2_CHOICE948_GROM
    );
  memtest2_CHOICE948_XUSED : X_BUF
    port map (
      I => memtest2_CHOICE948_FROM,
      O => memtest2_CHOICE948
    );
  memtest2_CHOICE948_YUSED : X_BUF
    port map (
      I => memtest2_CHOICE948_GROM,
      O => memtest2_CHOICE1071
    );
  maccontrol_Mmux_n0023_Result_11_6 : X_LUT4
    generic map(
      INIT => X"E000"
    )
    port map (
      ADR0 => maccontrol_phystat(11),
      ADR1 => maccontrol_addr_0_1,
      ADR2 => maccontrol_addr_1_1,
      ADR3 => maccontrol_N30199,
      O => maccontrol_CHOICE1385_FROM
    );
  maccontrol_Mmux_n0023_Result_7_6 : X_LUT4
    generic map(
      INIT => X"8880"
    )
    port map (
      ADR0 => maccontrol_addr_1_1,
      ADR1 => maccontrol_N30199,
      ADR2 => maccontrol_addr_0_1,
      ADR3 => maccontrol_phystat(7),
      O => maccontrol_CHOICE1385_GROM
    );
  maccontrol_CHOICE1385_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1385_FROM,
      O => maccontrol_CHOICE1385
    );
  maccontrol_CHOICE1385_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1385_GROM,
      O => maccontrol_CHOICE1364
    );
  memcontroller_dnout_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_8_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_8_OFF_RST,
      O => memcontroller_dnout(8)
    );
  MD_8_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_8_OFF_RST
    );
  maccontrol_Mmux_n0023_Result_0_56 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(0),
      ADR1 => maccontrol_n0085,
      ADR2 => maccontrol_n0083,
      ADR3 => maccontrol_lmacaddr(32),
      O => maccontrol_CHOICE1443_FROM
    );
  maccontrol_Mmux_n0023_Result_8_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(40),
      ADR1 => maccontrol_n0085,
      ADR2 => maccontrol_n0083,
      ADR3 => maccontrol_lmacaddr(8),
      O => maccontrol_CHOICE1443_GROM
    );
  maccontrol_CHOICE1443_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1443_FROM,
      O => maccontrol_CHOICE1443
    );
  maccontrol_CHOICE1443_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1443_GROM,
      O => maccontrol_CHOICE1525
    );
  maccontrol_Mmux_n0023_Result_13_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n0085,
      ADR1 => maccontrol_n00691_1,
      ADR2 => maccontrol_lmacaddr(45),
      ADR3 => maccontrol_phyaddr(13),
      O => maccontrol_CHOICE1323_FROM
    );
  maccontrol_Mmux_n0023_Result_9_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(41),
      ADR1 => maccontrol_phyaddr(9),
      ADR2 => maccontrol_n0085,
      ADR3 => maccontrol_n00691_1,
      O => maccontrol_CHOICE1323_GROM
    );
  maccontrol_CHOICE1323_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1323_FROM,
      O => maccontrol_CHOICE1323
    );
  maccontrol_CHOICE1323_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1323_GROM,
      O => maccontrol_CHOICE1285
    );
  maccontrol_Mmux_n0023_Result_13_9 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_N30212,
      ADR1 => maccontrol_N30192,
      ADR2 => maccontrol_phydi(13),
      ADR3 => maccontrol_lmacaddr(13),
      O => maccontrol_CHOICE1326_FROM
    );
  maccontrol_Mmux_n0023_Result_9_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_phydi(9),
      ADR1 => maccontrol_N30212,
      ADR2 => maccontrol_lmacaddr(9),
      ADR3 => maccontrol_N30192,
      O => maccontrol_CHOICE1326_GROM
    );
  maccontrol_CHOICE1326_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1326_FROM,
      O => maccontrol_CHOICE1326
    );
  maccontrol_CHOICE1326_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1326_GROM,
      O => maccontrol_CHOICE1288
    );
  maccontrol_PHY_status_miiaddr_1_1 : X_LUT4
    generic map(
      INIT => X"FEFA"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd5,
      ADR1 => maccontrol_PHY_status_N23512,
      ADR2 => maccontrol_PHY_status_cs_FFd6,
      ADR3 => maccontrol_PHY_status_addrl(1),
      O => maccontrol_PHY_status_miiaddr_1_FROM
    );
  maccontrol_PHY_status_miiaddr_0_1 : X_LUT4
    generic map(
      INIT => X"FFEF"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd5,
      ADR1 => maccontrol_PHY_status_addrl(0),
      ADR2 => maccontrol_PHY_status_N23512,
      ADR3 => maccontrol_PHY_status_cs_FFd6,
      O => maccontrol_PHY_status_miiaddr_1_GROM
    );
  maccontrol_PHY_status_miiaddr_1_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_miiaddr_1_FROM,
      O => maccontrol_PHY_status_miiaddr(1)
    );
  maccontrol_PHY_status_miiaddr_1_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_miiaddr_1_GROM,
      O => maccontrol_PHY_status_miiaddr(0)
    );
  maccontrol_PHY_status_miiaddr_2_1 : X_LUT4
    generic map(
      INIT => X"FEEE"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd5,
      ADR1 => maccontrol_PHY_status_cs_FFd6,
      ADR2 => maccontrol_PHY_status_N23512,
      ADR3 => maccontrol_PHY_status_addrl(2),
      O => maccontrol_PHY_status_miiaddr_2_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout178 : X_LUT4
    generic map(
      INIT => X"B080"
    )
    port map (
      ADR0 => maccontrol_PHY_status_din(4),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      ADR3 => maccontrol_PHY_status_miiaddr(2),
      O => maccontrol_PHY_status_miiaddr_2_GROM
    );
  maccontrol_PHY_status_miiaddr_2_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_miiaddr_2_FROM,
      O => maccontrol_PHY_status_miiaddr(2)
    );
  maccontrol_PHY_status_miiaddr_2_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_miiaddr_2_GROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE770
    );
  maccontrol_PHY_status_miiaddr_4_1 : X_LUT4
    generic map(
      INIT => X"0045"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd6,
      ADR1 => maccontrol_PHY_status_addrl(4),
      ADR2 => maccontrol_PHY_status_N23512,
      ADR3 => maccontrol_PHY_status_cs_FFd5,
      O => maccontrol_PHY_status_miiaddr_4_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout222 : X_LUT4
    generic map(
      INIT => X"B380"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR2 => maccontrol_PHY_status_din(6),
      ADR3 => maccontrol_PHY_status_miiaddr(4),
      O => maccontrol_PHY_status_miiaddr_4_GROM
    );
  maccontrol_PHY_status_miiaddr_4_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_miiaddr_4_FROM,
      O => maccontrol_PHY_status_miiaddr(4)
    );
  maccontrol_PHY_status_miiaddr_4_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_miiaddr_4_GROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE784
    );
  memcontroller_ts_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_8_TFF_RST,
      O => memcontroller_ts(8)
    );
  MD_8_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_8_TFF_RST
    );
  maccontrol_sclkll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_sclkll_FFY_RST
    );
  maccontrol_sclkll_721 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_sclkl,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => maccontrol_sclkll_FFY_RST,
      O => maccontrol_sclkll
    );
  maccontrol_phyaddr_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_25_FFY_RST
    );
  maccontrol_phyaddr_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(24),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_25_FFY_RST,
      O => maccontrol_phyaddr(24)
    );
  memcontroller_qn_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(9),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_9_IFF_RST,
      O => memcontroller_qn(9)
    );
  MD_9_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_9_IFF_RST
    );
  maccontrol_phyaddr_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_19_FFY_RST
    );
  maccontrol_phyaddr_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(18),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_19_FFY_RST,
      O => maccontrol_phyaddr(18)
    );
  maccontrol_phyaddr_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_29_FFY_RST
    );
  maccontrol_phyaddr_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(28),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_29_FFY_RST,
      O => maccontrol_phyaddr(28)
    );
  maccontrol_n003918 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_107,
      ADR1 => maccontrol_phyrstcnt_106,
      ADR2 => maccontrol_phyrstcnt_105,
      ADR3 => maccontrol_phyrstcnt_104,
      O => maccontrol_CHOICE1585_FROM
    );
  maccontrol_n0041161_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_107,
      ADR1 => maccontrol_phyrstcnt_98,
      ADR2 => maccontrol_phyrstcnt_99,
      ADR3 => maccontrol_phyrstcnt_106,
      O => maccontrol_CHOICE1585_GROM
    );
  maccontrol_CHOICE1585_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1585_FROM,
      O => maccontrol_CHOICE1585
    );
  maccontrol_CHOICE1585_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1585_GROM,
      O => maccontrol_N46406
    );
  txsim_SF227581 : X_LUT4
    generic map(
      INIT => X"0040"
    )
    port map (
      ADR0 => txsim_counter(5),
      ADR1 => txsim_counter(7),
      ADR2 => txsim_SF22756,
      ADR3 => txsim_counter(6),
      O => txsim_llltx_FROM
    );
  txsim_n0002_722 : X_LUT4
    generic map(
      INIT => X"F7C4"
    )
    port map (
      ADR0 => txsim_SF22756,
      ADR1 => txsim_llltx,
      ADR2 => txsim_N41883,
      ADR3 => txsim_SF22758,
      O => txsim_n0002
    );
  txsim_llltx_XUSED : X_BUF
    port map (
      I => txsim_llltx_FROM,
      O => txsim_SF22758
    );
  maccontrol_Mmux_n0023_Result_15_40_SW0 : X_LUT4
    generic map(
      INIT => X"ACA0"
    )
    port map (
      ADR0 => maccontrol_N46681,
      ADR1 => maccontrol_lmacaddr(15),
      ADR2 => maccontrol_addr(1),
      ADR3 => maccontrol_addr(0),
      O => maccontrol_Mmux_n0023_Result_15_40_SW0_O_FROM
    );
  maccontrol_Mmux_n0023_Result_15_40 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_N30212,
      ADR1 => maccontrol_N30192,
      ADR2 => maccontrol_CHOICE1410,
      ADR3 => maccontrol_Mmux_n0023_Result_15_40_SW0_O,
      O => maccontrol_Mmux_n0023_Result_15_40_SW0_O_GROM
    );
  maccontrol_Mmux_n0023_Result_15_40_SW0_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_15_40_SW0_O_FROM,
      O => maccontrol_Mmux_n0023_Result_15_40_SW0_O
    );
  maccontrol_Mmux_n0023_Result_15_40_SW0_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_15_40_SW0_O_GROM,
      O => maccontrol_CHOICE1418
    );
  memtest_llerr_BXMUX : X_INV
    port map (
      I => memtest_n0002,
      O => memtest_llerr_BXMUXNOT
    );
  memtest2_cs_0_BYMUX : X_INV
    port map (
      I => memtest2_cs(0),
      O => memtest2_cs_0_BYMUXNOT
    );
  memcontroller_dnl2_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_11_CEMUXNOT
    );
  memcontroller_dnout_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_9_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_9_OFF_RST,
      O => memcontroller_dnout(9)
    );
  MD_9_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_9_OFF_RST
    );
  memcontroller_dnl2_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_21_CEMUXNOT
    );
  memcontroller_dnl2_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_13_CEMUXNOT
    );
  memcontroller_dnl2_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_31_CEMUXNOT
    );
  memcontroller_dnl2_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_23_CEMUXNOT
    );
  memcontroller_dnl2_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_15_CEMUXNOT
    );
  memcontroller_ts_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_9_TFF_RST,
      O => memcontroller_ts(9)
    );
  MD_9_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_9_TFF_RST
    );
  memcontroller_dnl2_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_25_CEMUXNOT
    );
  memcontroller_dnl2_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_17_CEMUXNOT
    );
  memcontroller_dnl2_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_27_CEMUXNOT
    );
  memcontroller_dnl2_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_19_CEMUXNOT
    );
  memcontroller_dnl2_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_29_CEMUXNOT
    );
  maccontrol_PHY_status_MII_Interface_Ker202241 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => clkslen,
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => VCC,
      O => maccontrol_PHY_status_MII_Interface_N20226_FROM
    );
  maccontrol_PHY_status_MII_Interface_n00101 : X_LUT4
    generic map(
      INIT => X"F400"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_mdccnt(5),
      ADR1 => MDC_OBUF,
      ADR2 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => maccontrol_PHY_status_MII_Interface_N20226,
      O => maccontrol_PHY_status_MII_Interface_N20226_GROM
    );
  maccontrol_PHY_status_MII_Interface_N20226_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_N20226_FROM,
      O => maccontrol_PHY_status_MII_Interface_N20226
    );
  maccontrol_PHY_status_MII_Interface_N20226_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_N20226_GROM,
      O => maccontrol_PHY_status_MII_Interface_n0010
    );
  maccontrol_PHY_status_MII_Interface_Ker202191 : X_LUT4
    generic map(
      INIT => X"8080"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(1),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      ADR3 => VCC,
      O => maccontrol_PHY_status_MII_Interface_N20221_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout312 : X_LUT4
    generic map(
      INIT => X"B800"
    )
    port map (
      ADR0 => maccontrol_PHY_status_din(0),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      ADR2 => maccontrol_PHY_status_din(8),
      ADR3 => maccontrol_PHY_status_MII_Interface_N20221,
      O => maccontrol_PHY_status_MII_Interface_N20221_GROM
    );
  maccontrol_PHY_status_MII_Interface_N20221_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_N20221_FROM,
      O => maccontrol_PHY_status_MII_Interface_N20221
    );
  maccontrol_PHY_status_MII_Interface_N20221_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_N20221_GROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE800
    );
  LEDACT_723 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDACT_OD,
      CE => LEDACT_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => LEDACT_OFF_RST,
      O => LEDACT_OBUF
    );
  LEDACT_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDACT_OFF_RST
    );
  maccontrol_PHY_status_MII_Interface_n0079_SW0 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(1),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(5),
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      O => maccontrol_PHY_status_MII_Interface_N41816_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout27 : X_LUT4
    generic map(
      INIT => X"3120"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      ADR2 => maccontrol_PHY_status_din(7),
      ADR3 => maccontrol_PHY_status_din(15),
      O => maccontrol_PHY_status_MII_Interface_N41816_GROM
    );
  maccontrol_PHY_status_MII_Interface_N41816_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_N41816_FROM,
      O => maccontrol_PHY_status_MII_Interface_N41816
    );
  maccontrol_PHY_status_MII_Interface_N41816_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_N41816_GROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE741
    );
  maccontrol_PHY_status_MII_Interface_sout63 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      O => maccontrol_PHY_status_MII_Interface_CHOICE749_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout68 : X_LUT4
    generic map(
      INIT => X"AC00"
    )
    port map (
      ADR0 => maccontrol_PHY_status_din(2),
      ADR1 => maccontrol_PHY_status_din(10),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      ADR3 => maccontrol_PHY_status_MII_Interface_CHOICE749,
      O => maccontrol_PHY_status_MII_Interface_CHOICE749_GROM
    );
  maccontrol_PHY_status_MII_Interface_CHOICE749_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE749_FROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE749
    );
  maccontrol_PHY_status_MII_Interface_CHOICE749_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE749_GROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE750
    );
  maccontrol_PHY_status_MII_Interface_sout73 : X_LUT4
    generic map(
      INIT => X"FF54"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(0),
      ADR1 => maccontrol_PHY_status_MII_Interface_CHOICE741,
      ADR2 => maccontrol_PHY_status_MII_Interface_CHOICE735,
      ADR3 => maccontrol_PHY_status_MII_Interface_CHOICE750,
      O => maccontrol_PHY_status_MII_Interface_CHOICE751_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout498_2_724 : X_LUT4
    generic map(
      INIT => X"CFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(1),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR3 => maccontrol_PHY_status_MII_Interface_CHOICE751,
      O => maccontrol_PHY_status_MII_Interface_CHOICE751_GROM
    );
  maccontrol_PHY_status_MII_Interface_CHOICE751_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE751_FROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE751
    );
  maccontrol_PHY_status_MII_Interface_CHOICE751_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE751_GROM,
      O => maccontrol_PHY_status_MII_Interface_sout498_2
    );
  maccontrol_phydi_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_13_FFY_RST
    );
  maccontrol_phydi_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(12),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_13_FFY_RST,
      O => maccontrol_phydi(12)
    );
  maccontrol_phydi_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_15_FFY_RST
    );
  maccontrol_phydi_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(14),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_15_FFY_RST,
      O => maccontrol_phydi(14)
    );
  maccontrol_phydi_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_23_FFY_RST
    );
  maccontrol_phydi_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(23),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_23_FFY_RST,
      O => maccontrol_phydi(23)
    );
  maccontrol_phydi_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_25_FFY_RST
    );
  maccontrol_phydi_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(24),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_25_FFY_RST,
      O => maccontrol_phydi(24)
    );
  maccontrol_phydi_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_19_FFY_RST
    );
  maccontrol_phydi_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(18),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_19_FFY_RST,
      O => maccontrol_phydi(18)
    );
  maccontrol_phydi_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_27_FFY_RST
    );
  maccontrol_phydi_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(26),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_27_FFY_RST,
      O => maccontrol_phydi(26)
    );
  maccontrol_phydi_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_29_FFY_RST
    );
  maccontrol_phydi_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(28),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_29_FFY_RST,
      O => maccontrol_phydi(28)
    );
  maccontrol_phystat_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_1_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(0),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_1_FFY_RST,
      O => maccontrol_phystat(0)
    );
  maccontrol_phystat_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_3_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(2),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_3_FFY_RST,
      O => maccontrol_phystat(2)
    );
  testrx_n000410 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => testrx_CHOICE933,
      ADR3 => testrx_CHOICE930,
      O => testrx_cs_FFd1_FROM
    );
  testrx_cs_FFd1_In_725 : X_LUT4
    generic map(
      INIT => X"F575"
    )
    port map (
      ADR0 => testrx_N41780,
      ADR1 => testrx_rx_dvl,
      ADR2 => testrx_cs_FFd2,
      ADR3 => testrx_n0004,
      O => testrx_cs_FFd1_In
    );
  testrx_cs_FFd1_XUSED : X_BUF
    port map (
      I => testrx_cs_FFd1_FROM,
      O => testrx_n0004
    );
  maccontrol_Mmux_n0023_Result_15_40_SW0_SW0 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(31),
      ADR1 => maccontrol_addr(0),
      ADR2 => VCC,
      ADR3 => maccontrol_lmacaddr(47),
      O => maccontrol_N46681_FROM
    );
  maccontrol_Mmux_n0023_Result_11_40_SW0_SW0 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(43),
      ADR1 => maccontrol_addr(0),
      ADR2 => VCC,
      ADR3 => maccontrol_lmacaddr(27),
      O => maccontrol_N46681_GROM
    );
  maccontrol_N46681_XUSED : X_BUF
    port map (
      I => maccontrol_N46681_FROM,
      O => maccontrol_N46681
    );
  maccontrol_N46681_YUSED : X_BUF
    port map (
      I => maccontrol_N46681_GROM,
      O => maccontrol_N46685
    );
  maccontrol_LEDDPX : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDDPX_OD,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => LEDDPX_OFF_RST,
      O => maccontrol_LEDDPX_OBUF
    );
  LEDDPX_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDDPX_OFF_RST
    );
  txsim_n0002_SW0 : X_LUT4
    generic map(
      INIT => X"FF5F"
    )
    port map (
      ADR0 => txsim_counter(5),
      ADR1 => VCC,
      ADR2 => txsim_counter(6),
      ADR3 => txsim_counter(7),
      O => txsim_N41883_GROM
    );
  txsim_N41883_YUSED : X_BUF
    port map (
      I => txsim_N41883_GROM,
      O => txsim_N41883
    );
  maccontrol_Mmux_n0023_Result_14_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(14),
      ADR1 => maccontrol_lmacaddr(46),
      ADR2 => maccontrol_n0085,
      ADR3 => maccontrol_n0083,
      O => maccontrol_CHOICE1561_FROM
    );
  maccontrol_Mmux_n0023_Result_12_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n00691_1,
      ADR1 => maccontrol_n0085,
      ADR2 => maccontrol_phyaddr(12),
      ADR3 => maccontrol_lmacaddr(44),
      O => maccontrol_CHOICE1561_GROM
    );
  maccontrol_CHOICE1561_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1561_FROM,
      O => maccontrol_CHOICE1561
    );
  maccontrol_CHOICE1561_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1561_GROM,
      O => maccontrol_CHOICE1304
    );
  maccontrol_Mmux_n0023_Result_18_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_phydi(18),
      ADR1 => maccontrol_n0067,
      ADR2 => maccontrol_phystat(18),
      ADR3 => maccontrol_n0070,
      O => maccontrol_CHOICE1111_FROM
    );
  maccontrol_Mmux_n0023_Result_20_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_phydi(20),
      ADR1 => maccontrol_n0070,
      ADR2 => maccontrol_n0067,
      ADR3 => maccontrol_phystat(20),
      O => maccontrol_CHOICE1111_GROM
    );
  maccontrol_CHOICE1111_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1111_FROM,
      O => maccontrol_CHOICE1111
    );
  maccontrol_CHOICE1111_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1111_GROM,
      O => maccontrol_CHOICE1120
    );
  maccontrol_PHY_status_din_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_11_FFY_RST
    );
  maccontrol_PHY_status_din_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(10),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_11_FFY_RST,
      O => maccontrol_PHY_status_din(10)
    );
  maccontrol_PHY_status_din_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_13_FFY_RST
    );
  maccontrol_PHY_status_din_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(12),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_13_FFY_RST,
      O => maccontrol_PHY_status_din(12)
    );
  maccontrol_Mmux_n0023_Result_17_5 : X_LUT4
    generic map(
      INIT => X"3210"
    )
    port map (
      ADR0 => maccontrol_addr_0_1,
      ADR1 => maccontrol_addr_1_1,
      ADR2 => maccontrol_phyaddr(17),
      ADR3 => maccontrol_phydi(17),
      O => maccontrol_CHOICE1234_FROM
    );
  maccontrol_Mmux_n0023_Result_21_5 : X_LUT4
    generic map(
      INIT => X"3022"
    )
    port map (
      ADR0 => maccontrol_phyaddr(21),
      ADR1 => maccontrol_addr_1_1,
      ADR2 => maccontrol_phydi(21),
      ADR3 => maccontrol_addr_0_1,
      O => maccontrol_CHOICE1234_GROM
    );
  maccontrol_CHOICE1234_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1234_FROM,
      O => maccontrol_CHOICE1234
    );
  maccontrol_CHOICE1234_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1234_GROM,
      O => maccontrol_CHOICE1245
    );
  maccontrol_Mmux_n0023_Result_3_40 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_CHOICE1347,
      ADR1 => maccontrol_N46462,
      ADR2 => maccontrol_N30192,
      ADR3 => maccontrol_N30212,
      O => maccontrol_CHOICE1355_FROM
    );
  maccontrol_Mmux_n0023_Result_12_9 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_N30192,
      ADR1 => maccontrol_phydi(12),
      ADR2 => maccontrol_lmacaddr(12),
      ADR3 => maccontrol_N30212,
      O => maccontrol_CHOICE1355_GROM
    );
  maccontrol_CHOICE1355_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1355_FROM,
      O => maccontrol_CHOICE1355
    );
  maccontrol_CHOICE1355_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1355_GROM,
      O => maccontrol_CHOICE1307
    );
  maccontrol_Mmux_n0023_Result_29_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n00701_1,
      ADR1 => maccontrol_n0067,
      ADR2 => maccontrol_phydi(29),
      ADR3 => maccontrol_phystat(29),
      O => maccontrol_CHOICE1174_FROM
    );
  maccontrol_Mmux_n0023_Result_30_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_phystat(30),
      ADR1 => maccontrol_n00701_1,
      ADR2 => maccontrol_n00671_1,
      ADR3 => maccontrol_phydi(30),
      O => maccontrol_CHOICE1174_GROM
    );
  maccontrol_CHOICE1174_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1174_FROM,
      O => maccontrol_CHOICE1174
    );
  maccontrol_CHOICE1174_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1174_GROM,
      O => maccontrol_CHOICE1165
    );
  LEDRX_726 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDRX_LOGIC_ONE,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => LEDRX_N1683,
      O => LEDRX_OBUF
    );
  maccontrol_Mmux_n0023_Result_26_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n00701_1,
      ADR1 => maccontrol_phystat(26),
      ADR2 => maccontrol_phydi(26),
      ADR3 => maccontrol_n0067,
      O => maccontrol_CHOICE1147_FROM
    );
  maccontrol_Mmux_n0023_Result_22_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_phystat(22),
      ADR1 => maccontrol_phydi(22),
      ADR2 => maccontrol_n00701_1,
      ADR3 => maccontrol_n0067,
      O => maccontrol_CHOICE1147_GROM
    );
  maccontrol_CHOICE1147_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1147_FROM,
      O => maccontrol_CHOICE1147
    );
  maccontrol_CHOICE1147_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1147_GROM,
      O => maccontrol_CHOICE1129
    );
  maccontrol_Mmux_n0023_Result_16_5 : X_LUT4
    generic map(
      INIT => X"00CA"
    )
    port map (
      ADR0 => maccontrol_phyaddr(16),
      ADR1 => maccontrol_phydi(16),
      ADR2 => maccontrol_addr_0_1,
      ADR3 => maccontrol_addr_1_1,
      O => maccontrol_CHOICE1223_FROM
    );
  maccontrol_Mmux_n0023_Result_15_6 : X_LUT4
    generic map(
      INIT => X"8880"
    )
    port map (
      ADR0 => maccontrol_N30199,
      ADR1 => maccontrol_addr_1_1,
      ADR2 => maccontrol_addr_0_1,
      ADR3 => maccontrol_phystat(15),
      O => maccontrol_CHOICE1223_GROM
    );
  maccontrol_CHOICE1223_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1223_FROM,
      O => maccontrol_CHOICE1223
    );
  maccontrol_CHOICE1223_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1223_GROM,
      O => maccontrol_CHOICE1406
    );
  maccontrol_Mmux_n0023_Result_10_26_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_n0071,
      ADR1 => maccontrol_phydo(10),
      ADR2 => maccontrol_phydi(10),
      ADR3 => maccontrol_n0070,
      O => maccontrol_Mmux_n0023_Result_10_26_SW0_O_FROM
    );
  maccontrol_Mmux_n0023_Result_2_26_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n0070,
      ADR1 => maccontrol_phydo(2),
      ADR2 => maccontrol_phydi(2),
      ADR3 => maccontrol_n0071,
      O => maccontrol_Mmux_n0023_Result_10_26_SW0_O_GROM
    );
  maccontrol_Mmux_n0023_Result_10_26_SW0_O_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_10_26_SW0_O_FROM,
      O => maccontrol_Mmux_n0023_Result_10_26_SW0_O
    );
  maccontrol_Mmux_n0023_Result_10_26_SW0_O_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_10_26_SW0_O_GROM,
      O => maccontrol_Mmux_n0023_Result_2_26_SW0_O
    );
  memtest2_Mshreg_data4_13_srl_50 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_47,
      A1 => GLOBAL_LOGIC1_18,
      A2 => GLOBAL_LOGIC0_47,
      A3 => GLOBAL_LOGIC0_49,
      D => memtest2_ldata(13),
      CE => memtest2_n00511_3,
      CLK => clk,
      Q => memtest2_Mshreg_data4_13_net101_GSHIFT
    );
  memtest2_Mshreg_data4_13_net101_YUSED : X_BUF
    port map (
      I => memtest2_Mshreg_data4_13_net101_GSHIFT,
      O => memtest2_Mshreg_data4_13_net101
    );
  memtest2_Mshreg_data4_21_srl_42 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_27,
      A1 => GLOBAL_LOGIC1_17,
      A2 => GLOBAL_LOGIC0_25,
      A3 => GLOBAL_LOGIC0_25,
      D => memtest2_ldata(21),
      CE => memtest2_n00511_2,
      CLK => clk,
      Q => memtest2_Mshreg_data4_21_net85_GSHIFT
    );
  memtest2_Mshreg_data4_21_net85_YUSED : X_BUF
    port map (
      I => memtest2_Mshreg_data4_21_net85_GSHIFT,
      O => memtest2_Mshreg_data4_21_net85
    );
  maccontrol_Mmux_n0023_Result_24_5 : X_LUT4
    generic map(
      INIT => X"00CA"
    )
    port map (
      ADR0 => maccontrol_phyaddr(24),
      ADR1 => maccontrol_phydi(24),
      ADR2 => maccontrol_addr_0_1,
      ADR3 => maccontrol_addr_1_1,
      O => maccontrol_CHOICE1256_GROM
    );
  maccontrol_CHOICE1256_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1256_GROM,
      O => maccontrol_CHOICE1256
    );
  maccontrol_n00361 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_N30273,
      ADR1 => maccontrol_addr(7),
      ADR2 => maccontrol_n0084,
      ADR3 => maccontrol_newcmd,
      O => maccontrol_n0036_FROM
    );
  maccontrol_Mmux_n0023_Result_0_61 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(16),
      ADR1 => maccontrol_n0067,
      ADR2 => maccontrol_n0084,
      ADR3 => maccontrol_phystat(0),
      O => maccontrol_n0036_GROM
    );
  maccontrol_n0036_XUSED : X_BUF
    port map (
      I => maccontrol_n0036_FROM,
      O => maccontrol_n0036
    );
  maccontrol_n0036_YUSED : X_BUF
    port map (
      I => maccontrol_n0036_GROM,
      O => maccontrol_CHOICE1446
    );
  maccontrol_Mmux_n0023_Result_28_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_n0067,
      ADR1 => maccontrol_phystat(28),
      ADR2 => maccontrol_phydi(28),
      ADR3 => maccontrol_n00701_1,
      O => maccontrol_CHOICE1156_FROM
    );
  maccontrol_Mmux_n0023_Result_25_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => maccontrol_n0067,
      ADR1 => maccontrol_phystat(25),
      ADR2 => maccontrol_n00701_1,
      ADR3 => maccontrol_phydi(25),
      O => maccontrol_CHOICE1156_GROM
    );
  maccontrol_CHOICE1156_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1156_FROM,
      O => maccontrol_CHOICE1156
    );
  maccontrol_CHOICE1156_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1156_GROM,
      O => maccontrol_CHOICE1138
    );
  maccontrol_Mmux_n0023_Result_11_16 : X_LUT4
    generic map(
      INIT => X"3088"
    )
    port map (
      ADR0 => maccontrol_phydo(11),
      ADR1 => maccontrol_addr(1),
      ADR2 => maccontrol_phydi(11),
      ADR3 => maccontrol_addr(0),
      O => maccontrol_CHOICE1389_FROM
    );
  maccontrol_Mmux_n0023_Result_7_40_SW0_SW0 : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => maccontrol_lmacaddr(23),
      ADR1 => maccontrol_lmacaddr(39),
      ADR2 => maccontrol_addr(0),
      ADR3 => VCC,
      O => maccontrol_CHOICE1389_GROM
    );
  maccontrol_CHOICE1389_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1389_FROM,
      O => maccontrol_CHOICE1389
    );
  maccontrol_CHOICE1389_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1389_GROM,
      O => maccontrol_N46689
    );
  maccontrol_Mmux_n0023_Result_14_26_2_727 : X_LUT4
    generic map(
      INIT => X"ECEC"
    )
    port map (
      ADR0 => maccontrol_n0069,
      ADR1 => maccontrol_N30162,
      ADR2 => maccontrol_phyaddr(14),
      ADR3 => VCC,
      O => maccontrol_Mmux_n0023_Result_14_26_2_FROM
    );
  maccontrol_Mmux_n0023_Result_27_7 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_n00701_1,
      ADR1 => maccontrol_n0069,
      ADR2 => maccontrol_phyaddr(27),
      ADR3 => maccontrol_phydi(27),
      O => maccontrol_Mmux_n0023_Result_14_26_2_GROM
    );
  maccontrol_Mmux_n0023_Result_14_26_2_XUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_14_26_2_FROM,
      O => maccontrol_Mmux_n0023_Result_14_26_2
    );
  maccontrol_Mmux_n0023_Result_14_26_2_YUSED : X_BUF
    port map (
      I => maccontrol_Mmux_n0023_Result_14_26_2_GROM,
      O => maccontrol_CHOICE1214
    );
  maccontrol_n003977_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_113,
      ADR1 => maccontrol_phyrstcnt_114,
      ADR2 => maccontrol_phyrstcnt_112,
      ADR3 => maccontrol_phyrstcnt_111,
      O => maccontrol_N46402_FROM
    );
  maccontrol_n003977 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_n003963_O,
      ADR1 => maccontrol_CHOICE1603,
      ADR2 => maccontrol_CHOICE1596,
      ADR3 => maccontrol_N46402,
      O => maccontrol_N46402_GROM
    );
  maccontrol_N46402_XUSED : X_BUF
    port map (
      I => maccontrol_N46402_FROM,
      O => maccontrol_N46402
    );
  maccontrol_N46402_YUSED : X_BUF
    port map (
      I => maccontrol_N46402_GROM,
      O => maccontrol_CHOICE1605
    );
  maccontrol_Mmux_n0023_Result_15_16 : X_LUT4
    generic map(
      INIT => X"2C20"
    )
    port map (
      ADR0 => maccontrol_phydo(15),
      ADR1 => maccontrol_addr(0),
      ADR2 => maccontrol_addr(1),
      ADR3 => maccontrol_phydi(15),
      O => maccontrol_CHOICE1410_FROM
    );
  maccontrol_Mmux_n0023_Result_3_16 : X_LUT4
    generic map(
      INIT => X"3088"
    )
    port map (
      ADR0 => maccontrol_phydi(3),
      ADR1 => maccontrol_addr(0),
      ADR2 => maccontrol_phydo(3),
      ADR3 => maccontrol_addr(1),
      O => maccontrol_CHOICE1410_GROM
    );
  maccontrol_CHOICE1410_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1410_FROM,
      O => maccontrol_CHOICE1410
    );
  maccontrol_CHOICE1410_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1410_GROM,
      O => maccontrol_CHOICE1347
    );
  maccontrol_PHY_status_MII_Interface_sout330 : X_LUT4
    generic map(
      INIT => X"CE00"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_CHOICE793,
      ADR1 => maccontrol_PHY_status_MII_Interface_CHOICE800,
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(0),
      O => maccontrol_PHY_status_MII_Interface_CHOICE802_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout498 : X_LUT4
    generic map(
      INIT => X"FFEF"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_CHOICE831,
      ADR1 => maccontrol_PHY_status_MII_Interface_CHOICE764,
      ADR2 => maccontrol_PHY_status_MII_Interface_sout498_2,
      ADR3 => maccontrol_PHY_status_MII_Interface_CHOICE802,
      O => maccontrol_PHY_status_MII_Interface_CHOICE802_GROM
    );
  maccontrol_PHY_status_MII_Interface_CHOICE802_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE802_FROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE802
    );
  maccontrol_PHY_status_MII_Interface_CHOICE802_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE802_GROM,
      O => maccontrol_PHY_status_MII_Interface_sout
    );
  maccontrol_PHY_status_MII_Interface_sout361 : X_LUT4
    generic map(
      INIT => X"30B8"
    )
    port map (
      ADR0 => maccontrol_PHY_status_din(5),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR2 => maccontrol_PHY_status_miiaddr(3),
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      O => maccontrol_PHY_status_MII_Interface_CHOICE812_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout365 : X_LUT4
    generic map(
      INIT => X"FFA2"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR2 => maccontrol_PHY_status_din(1),
      ADR3 => maccontrol_PHY_status_MII_Interface_CHOICE812,
      O => maccontrol_PHY_status_MII_Interface_CHOICE812_GROM
    );
  maccontrol_PHY_status_MII_Interface_CHOICE812_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE812_FROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE812
    );
  maccontrol_PHY_status_MII_Interface_CHOICE812_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE812_GROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE813
    );
  maccontrol_PHY_status_MII_Interface_sout442 : X_LUT4
    generic map(
      INIT => X"0E0C"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      ADR1 => maccontrol_PHY_status_MII_Interface_CHOICE826,
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(0),
      ADR3 => maccontrol_PHY_status_MII_Interface_CHOICE813,
      O => maccontrol_PHY_status_MII_Interface_CHOICE829_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout472 : X_LUT4
    generic map(
      INIT => X"F333"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(5),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(1),
      ADR3 => maccontrol_PHY_status_MII_Interface_CHOICE829,
      O => maccontrol_PHY_status_MII_Interface_CHOICE829_GROM
    );
  maccontrol_PHY_status_MII_Interface_CHOICE829_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE829_FROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE829
    );
  maccontrol_PHY_status_MII_Interface_CHOICE829_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE829_GROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE831
    );
  maccontrol_Mmux_n0023_Result_12_65 : X_LUT4
    generic map(
      INIT => X"F070"
    )
    port map (
      ADR0 => maccontrol_sclkdeltall,
      ADR1 => maccontrol_N30218,
      ADR2 => maccontrol_dout(11),
      ADR3 => maccontrol_bitcnt_90,
      O => maccontrol_CHOICE1319_FROM
    );
  maccontrol_Mmux_n0023_Result_4_65 : X_LUT4
    generic map(
      INIT => X"F070"
    )
    port map (
      ADR0 => maccontrol_N30218,
      ADR1 => maccontrol_sclkdeltall,
      ADR2 => maccontrol_dout(3),
      ADR3 => maccontrol_bitcnt_90,
      O => maccontrol_CHOICE1319_GROM
    );
  maccontrol_CHOICE1319_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1319_FROM,
      O => maccontrol_CHOICE1319
    );
  maccontrol_CHOICE1319_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1319_GROM,
      O => maccontrol_CHOICE1281
    );
  maccontrol_Mmux_n0023_Result_7_16 : X_LUT4
    generic map(
      INIT => X"2C20"
    )
    port map (
      ADR0 => maccontrol_phydi(7),
      ADR1 => maccontrol_addr(1),
      ADR2 => maccontrol_addr(0),
      ADR3 => maccontrol_phydo(7),
      O => maccontrol_CHOICE1368_GROM
    );
  maccontrol_CHOICE1368_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1368_GROM,
      O => maccontrol_CHOICE1368
    );
  maccontrol_PHY_status_Ker235101 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd2,
      ADR1 => maccontrol_PHY_status_cs_FFd4,
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_cs_FFd3,
      O => maccontrol_PHY_status_N23512_FROM
    );
  maccontrol_PHY_status_miiaddr_3_1 : X_LUT4
    generic map(
      INIT => X"FEFC"
    )
    port map (
      ADR0 => maccontrol_PHY_status_addrl(3),
      ADR1 => maccontrol_PHY_status_cs_FFd5,
      ADR2 => maccontrol_PHY_status_cs_FFd6,
      ADR3 => maccontrol_PHY_status_N23512,
      O => maccontrol_PHY_status_N23512_GROM
    );
  maccontrol_PHY_status_N23512_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_N23512_FROM,
      O => maccontrol_PHY_status_N23512
    );
  maccontrol_PHY_status_N23512_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_N23512_GROM,
      O => maccontrol_PHY_status_miiaddr(3)
    );
  maccontrol_Mmux_n0023_Result_17_33 : X_LUT4
    generic map(
      INIT => X"CC4C"
    )
    port map (
      ADR0 => maccontrol_N30218,
      ADR1 => maccontrol_dout(16),
      ADR2 => maccontrol_sclkdeltall,
      ADR3 => maccontrol_bitcnt_90,
      O => maccontrol_CHOICE1240_FROM
    );
  maccontrol_Mmux_n0023_Result_9_65 : X_LUT4
    generic map(
      INIT => X"DF00"
    )
    port map (
      ADR0 => maccontrol_sclkdeltall,
      ADR1 => maccontrol_bitcnt_90,
      ADR2 => maccontrol_N30218,
      ADR3 => maccontrol_dout(8),
      O => maccontrol_CHOICE1240_GROM
    );
  maccontrol_CHOICE1240_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1240_FROM,
      O => maccontrol_CHOICE1240
    );
  maccontrol_CHOICE1240_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1240_GROM,
      O => maccontrol_CHOICE1300
    );
  maccontrol_PHY_status_Ker235181 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_cs_FFd6,
      ADR2 => maccontrol_PHY_status_cs_FFd5,
      ADR3 => VCC,
      O => maccontrol_PHY_status_N23520_FROM
    );
  maccontrol_PHY_status_n00201 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => clkslen,
      ADR1 => maccontrol_PHY_status_done,
      ADR2 => RESET_IBUF,
      ADR3 => maccontrol_PHY_status_N23520,
      O => maccontrol_PHY_status_N23520_GROM
    );
  maccontrol_PHY_status_N23520_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_N23520_FROM,
      O => maccontrol_PHY_status_N23520
    );
  maccontrol_PHY_status_N23520_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_N23520_GROM,
      O => maccontrol_PHY_status_n0020
    );
  memcontroller_addr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_10_OD,
      CE => MA_10_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_10_OFF_RST,
      O => memcontroller_ADDREXT(10)
    );
  MA_10_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_10_OFF_RST
    );
  maccontrol_PHY_status_MII_Interface_n00131 : X_LUT4
    generic map(
      INIT => X"AAA8"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_N20226,
      ADR1 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      ADR2 => maccontrol_PHY_status_MII_Interface_cs_FFd4,
      ADR3 => maccontrol_PHY_status_MII_Interface_cs_FFd3,
      O => maccontrol_PHY_status_MII_Interface_n0013_GROM
    );
  maccontrol_PHY_status_MII_Interface_n0013_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0013_GROM,
      O => maccontrol_PHY_status_MII_Interface_n0013
    );
  clken_n00051 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => clken_clkcnt(0),
      ADR2 => clken_clkcnt(2),
      ADR3 => clken_clkcnt(1),
      O => clken_clkcnt_0_FROM
    );
  clken_clkcnt_Madd_n0000_Mxor_Result_1_Result1 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => clken_clkcnt(0),
      ADR1 => VCC,
      ADR2 => clken_clkcnt(1),
      ADR3 => VCC,
      O => clken_clkcnt_n0000(1)
    );
  clken_clkcnt_0_BXMUX : X_INV
    port map (
      I => clken_clkcnt(0),
      O => clken_clkcnt_0_BXMUXNOT
    );
  clken_clkcnt_0_XUSED : X_BUF
    port map (
      I => clken_clkcnt_0_FROM,
      O => clken_n0005
    );
  maccontrol_n001223_1_728 : X_LUT4
    generic map(
      INIT => X"00A2"
    )
    port map (
      ADR0 => clkslen,
      ADR1 => maccontrol_N46628,
      ADR2 => maccontrol_CHOICE1055,
      ADR3 => RESET_IBUF,
      O => maccontrol_n001223_1_FROM
    );
  maccontrol_PHY_status_MII_Interface_n00161 : X_LUT4
    generic map(
      INIT => X"2020"
    )
    port map (
      ADR0 => clkslen,
      ADR1 => RESET_IBUF,
      ADR2 => maccontrol_PHY_status_MII_Interface_cs_FFd2,
      ADR3 => VCC,
      O => maccontrol_n001223_1_GROM
    );
  maccontrol_n001223_1_XUSED : X_BUF
    port map (
      I => maccontrol_n001223_1_FROM,
      O => maccontrol_n001223_1
    );
  maccontrol_n001223_1_YUSED : X_BUF
    port map (
      I => maccontrol_n001223_1_GROM,
      O => maccontrol_PHY_status_MII_Interface_n0016
    );
  maccontrol_PHY_status_MII_Interface_sts28 : X_LUT4
    generic map(
      INIT => X"4457"
    )
    port map (
      ADR0 => maccontrol_PHY_status_miirw,
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(0),
      ADR3 => maccontrol_PHY_status_MII_Interface_N46530,
      O => maccontrol_PHY_status_MII_Interface_CHOICE729_FROM
    );
  maccontrol_PHY_status_MII_Interface_sts35 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(5),
      ADR2 => VCC,
      ADR3 => maccontrol_PHY_status_MII_Interface_CHOICE729,
      O => maccontrol_PHY_status_MII_Interface_CHOICE729_GROM
    );
  maccontrol_PHY_status_MII_Interface_CHOICE729_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE729_FROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE729
    );
  maccontrol_PHY_status_MII_Interface_CHOICE729_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_CHOICE729_GROM,
      O => maccontrol_PHY_status_MII_Interface_sts
    );
  maccontrol_Mmux_n0023_Result_13_65 : X_LUT4
    generic map(
      INIT => X"C4CC"
    )
    port map (
      ADR0 => maccontrol_N30218,
      ADR1 => maccontrol_dout(12),
      ADR2 => maccontrol_bitcnt_90,
      ADR3 => maccontrol_sclkdeltall,
      O => maccontrol_CHOICE1338_FROM
    );
  maccontrol_Mmux_n0023_Result_21_33 : X_LUT4
    generic map(
      INIT => X"F700"
    )
    port map (
      ADR0 => maccontrol_N30218,
      ADR1 => maccontrol_sclkdeltall,
      ADR2 => maccontrol_bitcnt_90,
      ADR3 => maccontrol_dout(20),
      O => maccontrol_CHOICE1338_GROM
    );
  maccontrol_CHOICE1338_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1338_FROM,
      O => maccontrol_CHOICE1338
    );
  maccontrol_CHOICE1338_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1338_GROM,
      O => maccontrol_CHOICE1251
    );
  memcontroller_addr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_11_OD,
      CE => MA_11_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_11_OFF_RST,
      O => memcontroller_ADDREXT(11)
    );
  MA_11_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_11_OFF_RST
    );
  maccontrol_Mmux_n0023_Result_24_33 : X_LUT4
    generic map(
      INIT => X"BF00"
    )
    port map (
      ADR0 => maccontrol_bitcnt_90,
      ADR1 => maccontrol_sclkdeltall,
      ADR2 => maccontrol_N30218,
      ADR3 => maccontrol_dout(23),
      O => maccontrol_CHOICE1262_FROM
    );
  maccontrol_Mmux_n0023_Result_16_33 : X_LUT4
    generic map(
      INIT => X"8CCC"
    )
    port map (
      ADR0 => maccontrol_bitcnt_90,
      ADR1 => maccontrol_dout(15),
      ADR2 => maccontrol_N30218,
      ADR3 => maccontrol_sclkdeltall,
      O => maccontrol_CHOICE1262_GROM
    );
  maccontrol_CHOICE1262_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1262_FROM,
      O => maccontrol_CHOICE1262
    );
  maccontrol_CHOICE1262_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1262_GROM,
      O => maccontrol_CHOICE1229
    );
  memtest2_n0030_SW0 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memtest2_deql(2),
      ADR3 => memtest2_deql(3),
      O => memtest2_N41527_FROM
    );
  memtest2_n0030_729 : X_LUT4
    generic map(
      INIT => X"1333"
    )
    port map (
      ADR0 => memtest2_deql(1),
      ADR1 => memtest2_cs(0),
      ADR2 => memtest2_deql(0),
      ADR3 => memtest2_N41527,
      O => memtest2_N41527_GROM
    );
  memtest2_N41527_XUSED : X_BUF
    port map (
      I => memtest2_N41527_FROM,
      O => memtest2_N41527
    );
  memtest2_N41527_YUSED : X_BUF
    port map (
      I => memtest2_N41527_GROM,
      O => memtest2_n0030
    );
  maccontrol_PHY_status_n0019_SW0 : X_LUT4
    generic map(
      INIT => X"FFFB"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => maccontrol_PHY_status_done,
      ADR2 => maccontrol_PHY_status_cs_FFd4,
      ADR3 => maccontrol_PHY_status_cs_FFd2,
      O => maccontrol_PHY_status_N42089_GROM
    );
  maccontrol_PHY_status_N42089_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_N42089_GROM,
      O => maccontrol_PHY_status_N42089
    );
  txsim_SF2275642 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => txsim_counter(8),
      ADR1 => txsim_counter(16),
      ADR2 => txsim_counter(14),
      ADR3 => txsim_counter(13),
      O => txsim_CHOICE1098_GROM
    );
  txsim_CHOICE1098_YUSED : X_BUF
    port map (
      I => txsim_CHOICE1098_GROM,
      O => txsim_CHOICE1098
    );
  txsim_SF2275619 : X_LUT4
    generic map(
      INIT => X"0004"
    )
    port map (
      ADR0 => txsim_counter(10),
      ADR1 => txsim_counter(3),
      ADR2 => txsim_counter(0),
      ADR3 => txsim_counter(1),
      O => txsim_CHOICE1090_FROM
    );
  txsim_SF2275667 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => txsim_CHOICE1105,
      ADR1 => txsim_CHOICE1098,
      ADR2 => txsim_N46398,
      ADR3 => txsim_CHOICE1090,
      O => txsim_CHOICE1090_GROM
    );
  txsim_CHOICE1090_XUSED : X_BUF
    port map (
      I => txsim_CHOICE1090_FROM,
      O => txsim_CHOICE1090
    );
  txsim_CHOICE1090_YUSED : X_BUF
    port map (
      I => txsim_CHOICE1090_GROM,
      O => txsim_SF22756
    );
  txsim_SF2275655 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => txsim_counter(17),
      ADR1 => txsim_counter(11),
      ADR2 => txsim_counter(12),
      ADR3 => txsim_counter(15),
      O => txsim_CHOICE1105_GROM
    );
  txsim_CHOICE1105_YUSED : X_BUF
    port map (
      I => txsim_CHOICE1105_GROM,
      O => txsim_CHOICE1105
    );
  memtest2_MD_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(20),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_0_FFY_RST,
      O => d2(20)
    );
  d2_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_0_FFY_RST
    );
  memtest2_MD_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(0),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_0_FFX_RST,
      O => d2(0)
    );
  d2_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_0_FFX_RST
    );
  memtest2_MD_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(23),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_3_FFY_RST,
      O => d2(23)
    );
  d2_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_3_FFY_RST
    );
  memtest2_MD_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(3),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_3_FFX_RST,
      O => d2(3)
    );
  d2_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_3_FFX_RST
    );
  memtest2_Mshreg_data4_13_56_730 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_13_net101,
      CE => memtest2_n00511_3,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_13_56_FFX_RST,
      O => memtest2_Mshreg_data4_13_56
    );
  memtest2_Mshreg_data4_13_56_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_13_56_FFX_RST
    );
  memtest2_Mshreg_data4_21_48_731 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_21_net85,
      CE => memtest2_n00511_2,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_21_48_FFX_RST,
      O => memtest2_Mshreg_data4_21_48
    );
  memtest2_Mshreg_data4_21_48_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_21_48_FFX_RST
    );
  maccontrol_PHY_status_cs_FFd6_732 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_cs_FFd6_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_cs_FFd6_FFX_RST,
      O => maccontrol_PHY_status_cs_FFd6
    );
  maccontrol_PHY_status_cs_FFd6_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_cs_FFd6_FFX_RST
    );
  maccontrol_PHY_status_cs_FFd8_733 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => maccontrol_PHY_status_cs_FFd8_In,
      CE => clkslen,
      CLK => clk,
      SET => maccontrol_PHY_status_cs_FFd8_FFX_SET,
      RST => GND,
      O => maccontrol_PHY_status_cs_FFd8
    );
  maccontrol_PHY_status_cs_FFd8_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => maccontrol_PHY_status_cs_FFd8_FFX_SET
    );
  memtest2_Mshreg_data4_0_69_734 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_0_net127,
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_0_69_FFY_RST,
      O => memtest2_Mshreg_data4_0_69
    );
  memtest2_Mshreg_data4_0_69_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_0_69_FFY_RST
    );
  memtest2_Mshreg_data4_1_68_735 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_1_net125,
      CE => memtest2_n00511_3,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_1_68_FFY_RST,
      O => memtest2_Mshreg_data4_1_68
    );
  memtest2_Mshreg_data4_1_68_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_1_68_FFY_RST
    );
  maccontrol_Mshreg_sinlll_83_736 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mshreg_sinlll_net279,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => maccontrol_Mshreg_sinlll_83_FFY_RST,
      O => maccontrol_Mshreg_sinlll_83
    );
  maccontrol_Mshreg_sinlll_83_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_Mshreg_sinlll_83_FFY_RST
    );
  memtest_Mshreg_dataw4_10_27_737 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_10_net43,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_10_27_FFY_RST,
      O => memtest_Mshreg_dataw4_10_27
    );
  memtest_Mshreg_dataw4_10_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_10_27_FFY_RST
    );
  memtest2_Mshreg_data4_3_66_738 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_3_net121,
      CE => memtest2_n00511_1,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_3_66_FFY_RST,
      O => memtest2_Mshreg_data4_3_66
    );
  memtest2_Mshreg_data4_3_66_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_3_66_FFY_RST
    );
  memtest2_Mshreg_data4_2_67_739 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_2_net123,
      CE => memtest2_n00511_2,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_2_67_FFY_RST,
      O => memtest2_Mshreg_data4_2_67
    );
  memtest2_Mshreg_data4_2_67_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_2_67_FFY_RST
    );
  memtest_Mshreg_dataw4_11_26_740 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_11_net41,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_11_26_FFY_RST,
      O => memtest_Mshreg_dataw4_11_26
    );
  memtest_Mshreg_dataw4_11_26_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_11_26_FFY_RST
    );
  memtest_Mshreg_dataw4_12_25_741 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_12_net39,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_12_25_FFY_RST,
      O => memtest_Mshreg_dataw4_12_25
    );
  memtest_Mshreg_dataw4_12_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_12_25_FFY_RST
    );
  memcontroller_dnl1_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(19),
      CE => memcontroller_dnl1_19_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_19_FFX_RST,
      O => memcontroller_dnl1(19)
    );
  memcontroller_dnl1_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_19_FFX_RST
    );
  memcontroller_dnl1_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(29),
      CE => memcontroller_dnl1_29_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_29_FFX_RST,
      O => memcontroller_dnl1(29)
    );
  memcontroller_dnl1_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_29_FFX_RST
    );
  memtest2_datalfsr_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(0),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(1)
    );
  maccontrol_PHY_status_cs_FFd1_742 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_cs_FFd1_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_cs_FFd2_FFY_RST,
      O => maccontrol_PHY_status_cs_FFd1
    );
  maccontrol_PHY_status_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_cs_FFd2_FFY_RST
    );
  maccontrol_PHY_status_cs_FFd7_743 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_cs_FFd7_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_cs_FFd8_FFY_RST,
      O => maccontrol_PHY_status_cs_FFd7
    );
  maccontrol_PHY_status_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_cs_FFd8_FFY_RST
    );
  maccontrol_PHY_status_cs_FFd2_744 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_cs_FFd2_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_cs_FFd2_FFX_RST,
      O => maccontrol_PHY_status_cs_FFd2
    );
  maccontrol_PHY_status_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_cs_FFd2_FFX_RST
    );
  maccontrol_PHY_status_cs_FFd3_745 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_cs_FFd3_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_cs_FFd4_FFY_RST,
      O => maccontrol_PHY_status_cs_FFd3
    );
  maccontrol_PHY_status_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_cs_FFd4_FFY_RST
    );
  maccontrol_PHY_status_cs_FFd4_746 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_cs_FFd4_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_cs_FFd4_FFX_RST,
      O => maccontrol_PHY_status_cs_FFd4
    );
  maccontrol_PHY_status_cs_FFd4_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_cs_FFd4_FFX_RST
    );
  maccontrol_PHY_status_cs_FFd5_747 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_cs_FFd5_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_cs_FFd6_FFY_RST,
      O => maccontrol_PHY_status_cs_FFd5
    );
  maccontrol_PHY_status_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_cs_FFd6_FFY_RST
    );
  maccontrol_PHY_status_phyaddrws_748 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_phyaddrws_BYMUXNOT,
      CE => maccontrol_PHY_status_n00151_O,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_phyaddrws_FFY_RST,
      O => maccontrol_PHY_status_phyaddrws
    );
  maccontrol_PHY_status_phyaddrws_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_phyaddrws_FFY_RST
    );
  maccontrol_dout_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_12_68_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_12_FFY_RST,
      O => maccontrol_dout(12)
    );
  maccontrol_dout_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_12_FFY_RST
    );
  maccontrol_dout_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_20_22_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_20_FFY_RST,
      O => maccontrol_dout(20)
    );
  maccontrol_dout_20_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_20_FFY_RST
    );
  maccontrol_dout_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_21_36_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_21_FFY_RST,
      O => maccontrol_dout(21)
    );
  maccontrol_dout_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_21_FFY_RST
    );
  maccontrol_dout_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_22_22_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_22_FFY_RST,
      O => maccontrol_dout(22)
    );
  maccontrol_dout_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_22_FFY_RST
    );
  maccontrol_dout_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_13_68_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_13_FFY_RST,
      O => maccontrol_dout(13)
    );
  maccontrol_dout_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_13_FFY_RST
    );
  maccontrol_dout_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_30_22_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_30_FFY_RST,
      O => maccontrol_dout(30)
    );
  maccontrol_dout_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_30_FFY_RST
    );
  memcontroller_addr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_14_OD,
      CE => MA_14_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_14_OFF_RST,
      O => memcontroller_ADDREXT(14)
    );
  MA_14_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_14_OFF_RST
    );
  memtest2_addrlfsr_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(5),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(6)
    );
  memtest2_addrlfsr_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(7),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(8)
    );
  maccontrol_n00131_1_749 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_addr(7),
      ADR1 => maccontrol_n0070,
      ADR2 => maccontrol_N30273,
      ADR3 => maccontrol_newcmd,
      O => maccontrol_n00131_1_FROM
    );
  maccontrol_Mmux_n0023_Result_5_26_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => maccontrol_n0070,
      ADR1 => maccontrol_n0071,
      ADR2 => maccontrol_phydi(5),
      ADR3 => maccontrol_phydo(5),
      O => maccontrol_n00131_1_GROM
    );
  maccontrol_n00131_1_XUSED : X_BUF
    port map (
      I => maccontrol_n00131_1_FROM,
      O => maccontrol_n00131_1
    );
  maccontrol_n00131_1_YUSED : X_BUF
    port map (
      I => maccontrol_n00131_1_GROM,
      O => maccontrol_Mmux_n0023_Result_5_26_SW0_O
    );
  maccontrol_n0041111 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_110,
      ADR1 => maccontrol_phyrstcnt_108,
      ADR2 => maccontrol_phyrstcnt_92,
      ADR3 => maccontrol_phyrstcnt_109,
      O => maccontrol_CHOICE1033_GROM
    );
  maccontrol_CHOICE1033_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1033_GROM,
      O => maccontrol_CHOICE1033
    );
  maccontrol_PHY_status_MII_Interface_sout142_SW0 : X_LUT4
    generic map(
      INIT => X"C4F7"
    )
    port map (
      ADR0 => maccontrol_PHY_status_miiaddr(0),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(0),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(1),
      ADR3 => maccontrol_PHY_status_miiaddr(1),
      O => maccontrol_PHY_status_MII_Interface_N46538_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout142 : X_LUT4
    generic map(
      INIT => X"0200"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(2),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR2 => maccontrol_PHY_status_MII_Interface_N46538,
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      O => maccontrol_PHY_status_MII_Interface_N46538_GROM
    );
  maccontrol_PHY_status_MII_Interface_N46538_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_N46538_FROM,
      O => maccontrol_PHY_status_MII_Interface_N46538
    );
  maccontrol_PHY_status_MII_Interface_N46538_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_N46538_GROM,
      O => maccontrol_PHY_status_MII_Interface_CHOICE764
    );
  maccontrol_n0041135 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_103,
      ADR1 => maccontrol_phyrstcnt_102,
      ADR2 => maccontrol_phyrstcnt_112,
      ADR3 => maccontrol_phyrstcnt_111,
      O => maccontrol_CHOICE1041_GROM
    );
  maccontrol_CHOICE1041_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1041_GROM,
      O => maccontrol_CHOICE1041
    );
  maccontrol_n0041161 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => maccontrol_N46406,
      ADR1 => maccontrol_CHOICE1033,
      ADR2 => maccontrol_CHOICE1048,
      ADR3 => maccontrol_CHOICE1041,
      O => maccontrol_CHOICE1050_FROM
    );
  maccontrol_n0041194 : X_LUT4
    generic map(
      INIT => X"ECCC"
    )
    port map (
      ADR0 => maccontrol_CHOICE1003,
      ADR1 => maccontrol_phyrstcnt_122,
      ADR2 => maccontrol_CHOICE1018,
      ADR3 => maccontrol_CHOICE1050,
      O => maccontrol_CHOICE1050_GROM
    );
  maccontrol_CHOICE1050_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1050_FROM,
      O => maccontrol_CHOICE1050
    );
  maccontrol_CHOICE1050_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1050_GROM,
      O => maccontrol_n0041
    );
  maccontrol_Ker302041 : X_LUT4
    generic map(
      INIT => X"4040"
    )
    port map (
      ADR0 => maccontrol_addr(2),
      ADR1 => maccontrol_addr(3),
      ADR2 => maccontrol_addr(4),
      ADR3 => VCC,
      O => maccontrol_N30206_FROM
    );
  maccontrol_n00331 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_addr_0_1,
      ADR1 => maccontrol_addr_1_1,
      ADR2 => maccontrol_N30181,
      ADR3 => maccontrol_N30206,
      O => maccontrol_N30206_GROM
    );
  maccontrol_N30206_XUSED : X_BUF
    port map (
      I => maccontrol_N30206_FROM,
      O => maccontrol_N30206
    );
  maccontrol_N30206_YUSED : X_BUF
    port map (
      I => maccontrol_N30206_GROM,
      O => maccontrol_n0033
    );
  maccontrol_n0041148 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_105,
      ADR1 => maccontrol_phyrstcnt_100,
      ADR2 => maccontrol_phyrstcnt_104,
      ADR3 => maccontrol_phyrstcnt_91,
      O => maccontrol_CHOICE1048_GROM
    );
  maccontrol_CHOICE1048_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1048_GROM,
      O => maccontrol_CHOICE1048
    );
  maccontrol_Ker303031 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_addr(0),
      ADR2 => maccontrol_addr(1),
      ADR3 => VCC,
      O => maccontrol_N30305_FROM
    );
  maccontrol_n00691 : X_LUT4
    generic map(
      INIT => X"0200"
    )
    port map (
      ADR0 => maccontrol_addr(3),
      ADR1 => maccontrol_addr(4),
      ADR2 => maccontrol_addr(2),
      ADR3 => maccontrol_N30305,
      O => maccontrol_N30305_GROM
    );
  maccontrol_N30305_XUSED : X_BUF
    port map (
      I => maccontrol_N30305_FROM,
      O => maccontrol_N30305
    );
  maccontrol_N30305_YUSED : X_BUF
    port map (
      I => maccontrol_N30305_GROM,
      O => maccontrol_n0069
    );
  maccontrol_Ker302261 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_N30316,
      ADR1 => maccontrol_N30285,
      ADR2 => maccontrol_N30199,
      ADR3 => maccontrol_din(0),
      O => maccontrol_N30228_FROM
    );
  maccontrol_n00401 : X_LUT4
    generic map(
      INIT => X"0044"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => clkslen,
      ADR2 => VCC,
      ADR3 => maccontrol_N30228,
      O => maccontrol_N30228_GROM
    );
  maccontrol_N30228_XUSED : X_BUF
    port map (
      I => maccontrol_N30228_FROM,
      O => maccontrol_N30228
    );
  maccontrol_N30228_YUSED : X_BUF
    port map (
      I => maccontrol_N30228_GROM,
      O => maccontrol_n0040
    );
  memcontroller_addr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_15_OD,
      CE => MA_15_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_15_OFF_RST,
      O => memcontroller_ADDREXT(15)
    );
  MA_15_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_15_OFF_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_4_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(3),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_4_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(4)
    );
  maccontrol_PHY_status_MII_Interface_dreg_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_6_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(5),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_6_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(6)
    );
  maccontrol_PHY_status_MII_Interface_dreg_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_8_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(7),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_8_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(8)
    );
  maccontrol_PHY_status_MII_Interface_dreg_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_8_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(6),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_8_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(7)
    );
  maccontrol_PHY_status_MII_Interface_dreg_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_10_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(9),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_10_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(10)
    );
  maccontrol_PHY_status_MII_Interface_dreg_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_10_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(8),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_10_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(9)
    );
  memtest_addrcntl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_11_FFX_RST
    );
  memtest_addrcntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(11),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_11_FFX_RST,
      O => memtest_addrcntl(11)
    );
  memtest_addrcntl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_11_FFY_RST
    );
  memtest_addrcntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(10),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_11_FFY_RST,
      O => memtest_addrcntl(10)
    );
  memtest_addrcntl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_13_FFX_RST
    );
  memtest_addrcntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(13),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_13_FFX_RST,
      O => memtest_addrcntl(13)
    );
  memtest_addrcntl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_13_FFY_RST
    );
  memtest_addrcntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(12),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_13_FFY_RST,
      O => memtest_addrcntl(12)
    );
  maccontrol_n004121 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_116,
      ADR1 => maccontrol_phyrstcnt_118,
      ADR2 => maccontrol_phyrstcnt_115,
      ADR3 => maccontrol_phyrstcnt_117,
      O => maccontrol_CHOICE1002_FROM
    );
  maccontrol_n004126 : X_LUT4
    generic map(
      INIT => X"0100"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_101,
      ADR1 => maccontrol_phyrstcnt_114,
      ADR2 => maccontrol_phyrstcnt_113,
      ADR3 => maccontrol_CHOICE1002,
      O => maccontrol_CHOICE1002_GROM
    );
  maccontrol_CHOICE1002_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1002_FROM,
      O => maccontrol_CHOICE1002
    );
  maccontrol_CHOICE1002_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1002_GROM,
      O => maccontrol_CHOICE1003
    );
  memtest_addrcntl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_15_FFX_RST
    );
  memtest_addrcntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(15),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_15_FFX_RST,
      O => memtest_addrcntl(15)
    );
  memtest_addrcntl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_15_FFY_RST
    );
  memtest_addrcntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(14),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_15_FFY_RST,
      O => memtest_addrcntl(14)
    );
  maccontrol_n0039102 : X_LUT4
    generic map(
      INIT => X"00FE"
    )
    port map (
      ADR0 => maccontrol_CHOICE1605,
      ADR1 => maccontrol_CHOICE1589,
      ADR2 => maccontrol_CHOICE1582,
      ADR3 => maccontrol_phyrstcnt_122,
      O => maccontrol_CHOICE1608_FROM
    );
  maccontrol_n0039124 : X_LUT4
    generic map(
      INIT => X"5040"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => maccontrol_N30228,
      ADR2 => clkslen,
      ADR3 => maccontrol_CHOICE1608,
      O => maccontrol_CHOICE1608_GROM
    );
  maccontrol_CHOICE1608_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1608_FROM,
      O => maccontrol_CHOICE1608
    );
  maccontrol_CHOICE1608_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1608_GROM,
      O => maccontrol_n0039
    );
  memcontroller_n00081 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => memcontroller_clknum_0_1,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => VCC,
      O => clken1_FROM
    );
  memcontroller_n00011 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => memcontroller_clknum_0_1,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => VCC,
      O => clken1_GROM
    );
  clken1_XUSED : X_BUF
    port map (
      I => clken1_FROM,
      O => clken1
    );
  clken1_YUSED : X_BUF
    port map (
      I => clken1_GROM,
      O => clken4
    );
  maccontrol_PHY_status_dout_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_11_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(10),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_11_FFY_RST,
      O => maccontrol_PHY_status_dout(10)
    );
  maccontrol_n00111 : X_LUT4
    generic map(
      INIT => X"0020"
    )
    port map (
      ADR0 => maccontrol_sclkdelta,
      ADR1 => RESET_IBUF,
      ADR2 => clkslen,
      ADR3 => maccontrol_N30311,
      O => maccontrol_n0011_FROM
    );
  maccontrol_n00101 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => maccontrol_sclkdelta,
      ADR1 => RESET_IBUF,
      ADR2 => clkslen,
      ADR3 => maccontrol_N30311,
      O => maccontrol_n0011_GROM
    );
  maccontrol_n0011_XUSED : X_BUF
    port map (
      I => maccontrol_n0011_FROM,
      O => maccontrol_n0011
    );
  maccontrol_n0011_YUSED : X_BUF
    port map (
      I => maccontrol_n0011_GROM,
      O => maccontrol_n0010
    );
  maccontrol_n003963 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_121,
      ADR1 => maccontrol_phyrstcnt_93,
      ADR2 => maccontrol_phyrstcnt_120,
      ADR3 => maccontrol_phyrstcnt_119,
      O => maccontrol_n003963_O_FROM
    );
  maccontrol_n004144 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_121,
      ADR1 => maccontrol_phyrstcnt_93,
      ADR2 => maccontrol_phyrstcnt_120,
      ADR3 => maccontrol_phyrstcnt_119,
      O => maccontrol_n003963_O_GROM
    );
  maccontrol_n003963_O_XUSED : X_BUF
    port map (
      I => maccontrol_n003963_O_FROM,
      O => maccontrol_n003963_O
    );
  maccontrol_n003963_O_YUSED : X_BUF
    port map (
      I => maccontrol_n003963_O_GROM,
      O => maccontrol_CHOICE1010
    );
  maccontrol_PHY_status_miirw1 : X_LUT4
    generic map(
      INIT => X"0040"
    )
    port map (
      ADR0 => maccontrol_PHY_status_cs_FFd5,
      ADR1 => maccontrol_PHY_status_rwl,
      ADR2 => maccontrol_PHY_status_N23512,
      ADR3 => maccontrol_PHY_status_cs_FFd6,
      O => maccontrol_PHY_status_miirw_FROM
    );
  maccontrol_PHY_status_MII_Interface_sout273_SW2 : X_LUT4
    generic map(
      INIT => X"0B08"
    )
    port map (
      ADR0 => maccontrol_PHY_status_din(12),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR2 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      ADR3 => maccontrol_PHY_status_miirw,
      O => maccontrol_PHY_status_miirw_GROM
    );
  maccontrol_PHY_status_miirw_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_miirw_FROM,
      O => maccontrol_PHY_status_miirw
    );
  maccontrol_PHY_status_miirw_YUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_miirw_GROM,
      O => maccontrol_PHY_status_MII_Interface_N46672
    );
  memcontroller_n00071 : X_LUT4
    generic map(
      INIT => X"5000"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_n0007_FROM
    );
  memcontroller_n00051 : X_LUT4
    generic map(
      INIT => X"0050"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_0_2,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_n0007_GROM
    );
  memcontroller_n0007_XUSED : X_BUF
    port map (
      I => memcontroller_n0007_FROM,
      O => memcontroller_n0007
    );
  memcontroller_n0007_YUSED : X_BUF
    port map (
      I => memcontroller_n0007_GROM,
      O => memcontroller_n0005
    );
  maccontrol_n004157 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_95,
      ADR1 => maccontrol_phyrstcnt_96,
      ADR2 => maccontrol_phyrstcnt_97,
      ADR3 => maccontrol_phyrstcnt_94,
      O => maccontrol_CHOICE1017_FROM
    );
  maccontrol_n004158 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => maccontrol_CHOICE1010,
      ADR3 => maccontrol_CHOICE1017,
      O => maccontrol_CHOICE1017_GROM
    );
  maccontrol_CHOICE1017_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1017_FROM,
      O => maccontrol_CHOICE1017
    );
  maccontrol_CHOICE1017_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1017_GROM,
      O => maccontrol_CHOICE1018
    );
  memcontroller_addr_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_16_OD,
      CE => MA_16_OCEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => MA_16_OFF_RST,
      O => memcontroller_ADDREXT(16)
    );
  MA_16_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MA_16_OFF_RST
    );
  maccontrol_n00311_1_750 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_newcmd,
      ADR1 => maccontrol_addr(7),
      ADR2 => maccontrol_N30273,
      ADR3 => maccontrol_n0069,
      O => maccontrol_n00311_1_FROM
    );
  maccontrol_n00311 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_addr(7),
      ADR1 => maccontrol_n0069,
      ADR2 => maccontrol_newcmd,
      ADR3 => maccontrol_N30273,
      O => maccontrol_n00311_1_GROM
    );
  maccontrol_n00311_1_XUSED : X_BUF
    port map (
      I => maccontrol_n00311_1_FROM,
      O => maccontrol_n00311_1
    );
  maccontrol_n00311_1_YUSED : X_BUF
    port map (
      I => maccontrol_n00311_1_GROM,
      O => maccontrol_n0031
    );
  maccontrol_SOUT : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => SOUT_OD,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => SOUT_OFF_RST,
      O => maccontrol_SOUT_OBUF
    );
  SOUT_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => SOUT_OFF_RST
    );
  maccontrol_n00431 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => maccontrol_phystat(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_phystat(4),
      O => maccontrol_n0043_FROM
    );
  maccontrol_n00421 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => maccontrol_phystat(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => maccontrol_phystat(4),
      O => maccontrol_n0043_GROM
    );
  maccontrol_n0043_XUSED : X_BUF
    port map (
      I => maccontrol_n0043_FROM,
      O => maccontrol_n0043
    );
  maccontrol_n0043_YUSED : X_BUF
    port map (
      I => maccontrol_n0043_GROM,
      O => maccontrol_n0042
    );
  maccontrol_n00371 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_n0085,
      ADR1 => maccontrol_newcmd,
      ADR2 => maccontrol_addr(7),
      ADR3 => maccontrol_N30273,
      O => maccontrol_n0037_FROM
    );
  maccontrol_n00351 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_n0083,
      ADR1 => maccontrol_newcmd,
      ADR2 => maccontrol_addr(7),
      ADR3 => maccontrol_N30273,
      O => maccontrol_n0037_GROM
    );
  maccontrol_n0037_XUSED : X_BUF
    port map (
      I => maccontrol_n0037_FROM,
      O => maccontrol_n0037
    );
  maccontrol_n0037_YUSED : X_BUF
    port map (
      I => maccontrol_n0037_GROM,
      O => maccontrol_n0035
    );
  maccontrol_n00521 : X_LUT4
    generic map(
      INIT => X"8080"
    )
    port map (
      ADR0 => maccontrol_bitcnt_90,
      ADR1 => maccontrol_sclkdeltal,
      ADR2 => maccontrol_N30218,
      ADR3 => VCC,
      O => maccontrol_newcmd_FROM
    );
  maccontrol_n00131 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_addr(7),
      ADR1 => maccontrol_n0070,
      ADR2 => maccontrol_N30273,
      ADR3 => maccontrol_newcmd,
      O => maccontrol_newcmd_GROM
    );
  maccontrol_newcmd_XUSED : X_BUF
    port map (
      I => maccontrol_newcmd_FROM,
      O => maccontrol_newcmd
    );
  maccontrol_newcmd_YUSED : X_BUF
    port map (
      I => maccontrol_newcmd_GROM,
      O => maccontrol_n0013
    );
  maccontrol_n006412 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => maccontrol_ledtx_cnt_133,
      ADR1 => maccontrol_ledtx_cnt_132,
      ADR2 => maccontrol_ledtx_cnt_131,
      ADR3 => maccontrol_ledtx_cnt_134,
      O => maccontrol_CHOICE974_GROM
    );
  maccontrol_CHOICE974_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE974_GROM,
      O => maccontrol_CHOICE974
    );
  maccontrol_n00541 : X_LUT4
    generic map(
      INIT => X"3000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => maccontrol_bitcnt_90,
      ADR2 => maccontrol_N30218,
      ADR3 => maccontrol_sclkdeltall,
      O => maccontrol_CHOICE1055_FROM
    );
  maccontrol_n001223 : X_LUT4
    generic map(
      INIT => X"5010"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => maccontrol_N46628,
      ADR2 => clkslen,
      ADR3 => maccontrol_CHOICE1055,
      O => maccontrol_CHOICE1055_GROM
    );
  maccontrol_CHOICE1055_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1055_FROM,
      O => maccontrol_CHOICE1055
    );
  maccontrol_CHOICE1055_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1055_GROM,
      O => maccontrol_n0012
    );
  testrx_MACDATA_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_0_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_0_OFF_RST,
      O => testrx_MACDATA_0_OBUF
    );
  MACDATA_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_0_OFF_RST
    );
  maccontrol_n003951 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_115,
      ADR1 => maccontrol_phyrstcnt_117,
      ADR2 => maccontrol_phyrstcnt_116,
      ADR3 => maccontrol_phyrstcnt_118,
      O => maccontrol_CHOICE1596_GROM
    );
  maccontrol_CHOICE1596_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1596_GROM,
      O => maccontrol_CHOICE1596
    );
  maccontrol_n00701 : X_LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      ADR0 => maccontrol_addr(4),
      ADR1 => maccontrol_addr(2),
      ADR2 => maccontrol_N30285,
      ADR3 => maccontrol_addr(3),
      O => maccontrol_n0070_FROM
    );
  maccontrol_Mmux_n0023_Result_19_7 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => maccontrol_phydi(19),
      ADR1 => maccontrol_n0069,
      ADR2 => maccontrol_phyaddr(19),
      ADR3 => maccontrol_n0070,
      O => maccontrol_n0070_GROM
    );
  maccontrol_n0070_XUSED : X_BUF
    port map (
      I => maccontrol_n0070_FROM,
      O => maccontrol_n0070
    );
  maccontrol_n0070_YUSED : X_BUF
    port map (
      I => maccontrol_n0070_GROM,
      O => maccontrol_CHOICE1194
    );
  maccontrol_n006425 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => maccontrol_ledtx_cnt_123,
      ADR1 => maccontrol_ledtx_cnt_126,
      ADR2 => maccontrol_ledtx_cnt_125,
      ADR3 => maccontrol_ledtx_cnt_124,
      O => maccontrol_CHOICE981_FROM
    );
  maccontrol_n00451 : X_LUT4
    generic map(
      INIT => X"5FFF"
    )
    port map (
      ADR0 => maccontrol_CHOICE974,
      ADR1 => VCC,
      ADR2 => maccontrol_CHOICE988,
      ADR3 => maccontrol_CHOICE981,
      O => maccontrol_CHOICE981_GROM
    );
  maccontrol_CHOICE981_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE981_FROM,
      O => maccontrol_CHOICE981
    );
  maccontrol_CHOICE981_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE981_GROM,
      O => maccontrol_n0045
    );
  maccontrol_PHY_status_MII_Interface_n0004_751 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(4),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(5),
      ADR2 => maccontrol_PHY_status_MII_Interface_n0004_2,
      ADR3 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      O => maccontrol_PHY_status_MII_Interface_cs_FFd2_FROM
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => maccontrol_PHY_status_MII_Interface_cs_FFd3,
      ADR3 => maccontrol_PHY_status_MII_Interface_n0004,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd2_In
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd2_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_cs_FFd2_FROM,
      O => maccontrol_PHY_status_MII_Interface_n0004
    );
  maccontrol_n006438 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => maccontrol_ledtx_cnt_130,
      ADR1 => maccontrol_ledtx_cnt_128,
      ADR2 => maccontrol_ledtx_cnt_127,
      ADR3 => maccontrol_ledtx_cnt_129,
      O => maccontrol_CHOICE988_FROM
    );
  maccontrol_n00441 : X_LUT4
    generic map(
      INIT => X"7F00"
    )
    port map (
      ADR0 => maccontrol_CHOICE981,
      ADR1 => maccontrol_CHOICE988,
      ADR2 => maccontrol_CHOICE974,
      ADR3 => maccontrol_N30273,
      O => maccontrol_CHOICE988_GROM
    );
  maccontrol_CHOICE988_XUSED : X_BUF
    port map (
      I => maccontrol_CHOICE988_FROM,
      O => maccontrol_CHOICE988
    );
  maccontrol_CHOICE988_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE988_GROM,
      O => maccontrol_n0044
    );
  maccontrol_n02341 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => maccontrol_N30285,
      ADR1 => maccontrol_Ker303141_2,
      ADR2 => clkslen,
      ADR3 => maccontrol_N30206,
      O => maccontrol_n0234_GROM
    );
  maccontrol_n0234_YUSED : X_BUF
    port map (
      I => maccontrol_n0234_GROM,
      O => maccontrol_n0234
    );
  maccontrol_n003968 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => maccontrol_phyrstcnt_97,
      ADR1 => maccontrol_phyrstcnt_94,
      ADR2 => maccontrol_phyrstcnt_96,
      ADR3 => maccontrol_phyrstcnt_95,
      O => maccontrol_CHOICE1603_GROM
    );
  maccontrol_CHOICE1603_YUSED : X_BUF
    port map (
      I => maccontrol_CHOICE1603_GROM,
      O => maccontrol_CHOICE1603
    );
  maccontrol_n00681 : X_LUT4
    generic map(
      INIT => X"0004"
    )
    port map (
      ADR0 => maccontrol_addr(2),
      ADR1 => maccontrol_N30299,
      ADR2 => maccontrol_addr(3),
      ADR3 => maccontrol_addr(4),
      O => maccontrol_n0068_GROM
    );
  maccontrol_n0068_YUSED : X_BUF
    port map (
      I => maccontrol_n0068_GROM,
      O => maccontrol_n0068
    );
  memtest2_laddr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_3_FFY_RST
    );
  memtest2_laddr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(2),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_3_FFY_RST,
      O => memtest2_laddr(2)
    );
  memtest2_n01171 : X_LUT4
    generic map(
      INIT => X"C0D0"
    )
    port map (
      ADR0 => memtest2_cs(0),
      ADR1 => memtest2_N22660,
      ADR2 => memcontroller_Ker256691_O,
      ADR3 => memtest2_n0025,
      O => memtest2_n0117_FROM
    );
  memtest2_n00111 : X_LUT4
    generic map(
      INIT => X"F040"
    )
    port map (
      ADR0 => memtest2_cs(0),
      ADR1 => memtest2_n0027,
      ADR2 => memcontroller_Ker256691_O,
      ADR3 => memtest2_N22660,
      O => memtest2_n0117_GROM
    );
  memtest2_n0117_XUSED : X_BUF
    port map (
      I => memtest2_n0117_FROM,
      O => memtest2_n0117
    );
  memtest2_n0117_YUSED : X_BUF
    port map (
      I => memtest2_n0117_GROM,
      O => memtest2_n0011
    );
  memtest2_laddr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_5_FFY_RST
    );
  memtest2_laddr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(4),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_5_FFY_RST,
      O => memtest2_laddr(4)
    );
  memtest2_laddr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_13_FFY_RST
    );
  memtest2_laddr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(12),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_13_FFY_RST,
      O => memtest2_laddr(12)
    );
  memtest2_laddr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_15_FFY_RST
    );
  memtest2_laddr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(14),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_15_FFY_RST,
      O => memtest2_laddr(14)
    );
  maccontrol_PHY_status_MII_Interface_statecnt_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_statecnt_1_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_statecnt_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0014(1),
      CE => maccontrol_PHY_status_MII_Interface_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_statecnt_1_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_statecnt(1)
    );
  maccontrol_PHY_status_MII_Interface_n0079_752 : X_LUT4
    generic map(
      INIT => X"070F"
    )
    port map (
      ADR0 => maccontrol_PHY_status_MII_Interface_statecnt(3),
      ADR1 => maccontrol_PHY_status_MII_Interface_statecnt(0),
      ADR2 => maccontrol_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => maccontrol_PHY_status_MII_Interface_N41816,
      O => maccontrol_PHY_status_MII_Interface_statecnt_1_FROM
    );
  maccontrol_PHY_status_MII_Interface_n0014_1_1 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => maccontrol_PHY_status_MII_Interface_n0078(1),
      ADR3 => maccontrol_PHY_status_MII_Interface_n0079,
      O => maccontrol_PHY_status_MII_Interface_n0014(1)
    );
  maccontrol_PHY_status_MII_Interface_statecnt_1_XUSED : X_BUF
    port map (
      I => maccontrol_PHY_status_MII_Interface_statecnt_1_FROM,
      O => maccontrol_PHY_status_MII_Interface_n0079
    );
  memtest2_n002112 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => memtest2_cnt(10),
      ADR1 => memtest2_cnt(15),
      ADR2 => memtest2_cnt(1),
      ADR3 => memtest2_cnt(14),
      O => memtest2_CHOICE941_GROM
    );
  memtest2_CHOICE941_YUSED : X_BUF
    port map (
      I => memtest2_CHOICE941_GROM,
      O => memtest2_CHOICE941
    );
  testrx_MACDATA_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_1_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_1_OFF_RST,
      O => testrx_MACDATA_1_OBUF
    );
  MACDATA_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_1_OFF_RST
    );
  LEDRX_Sclr_INV1 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => RX_ER_IBUF,
      ADR1 => VCC,
      ADR2 => RX_DV_IBUF,
      ADR3 => VCC,
      O => LEDRX_N1683_GROM
    );
  LEDRX_N1683_YUSED : X_BUF
    port map (
      I => LEDRX_N1683_GROM,
      O => LEDRX_N1683
    );
  memtest2_n01191 : X_LUT4
    generic map(
      INIT => X"C0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memtest2_cs(0),
      ADR2 => memcontroller_Ker256691_O,
      ADR3 => memtest2_n0028,
      O => memtest2_n0119_GROM
    );
  memtest2_n0119_YUSED : X_BUF
    port map (
      I => memtest2_n0119_GROM,
      O => memtest2_n0119
    );
  memcontroller_clknum_1_BYMUX : X_INV
    port map (
      I => memcontroller_clknum_0_2,
      O => memcontroller_clknum_1_BYMUXNOT
    );
  maccontrol_Ker30216_SW1 : X_LUT4
    generic map(
      INIT => X"BFFF"
    )
    port map (
      ADR0 => maccontrol_bitcnt_86,
      ADR1 => maccontrol_sclkdeltal,
      ADR2 => maccontrol_addr(7),
      ADR3 => maccontrol_bitcnt_90,
      O => maccontrol_N46368_FROM
    );
  maccontrol_Ker303141 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => maccontrol_bitcnt_88,
      ADR1 => maccontrol_bitcnt_89,
      ADR2 => maccontrol_N42043,
      ADR3 => maccontrol_N46368,
      O => maccontrol_N46368_GROM
    );
  maccontrol_N46368_XUSED : X_BUF
    port map (
      I => maccontrol_N46368_FROM,
      O => maccontrol_N46368
    );
  maccontrol_N46368_YUSED : X_BUF
    port map (
      I => maccontrol_N46368_GROM,
      O => maccontrol_N30316
    );
  clken_lclken_LOGIC_ONE_753 : X_ONE
    port map (
      O => clken_lclken_LOGIC_ONE
    );
  testrx_MACDATA_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_2_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_2_OFF_RST,
      O => testrx_MACDATA_2_OBUF
    );
  MACDATA_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_2_OFF_RST
    );
  testrx_MACDATA_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_3_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_3_OFF_RST,
      O => testrx_MACDATA_3_OBUF
    );
  MACDATA_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_3_OFF_RST
    );
  testrx_MACDATA_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_4_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_4_OFF_RST,
      O => testrx_MACDATA_4_OBUF
    );
  MACDATA_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_4_OFF_RST
    );
  testrx_MACDATA_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_5_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_5_OFF_RST,
      O => testrx_MACDATA_5_OBUF
    );
  MACDATA_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_5_OFF_RST
    );
  testrx_MACDATA_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_6_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_6_OFF_RST,
      O => testrx_MACDATA_6_OBUF
    );
  MACDATA_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_6_OFF_RST
    );
  testrx_MACDATA_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_7_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_7_OFF_RST,
      O => testrx_MACDATA_7_OBUF
    );
  MACDATA_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_7_OFF_RST
    );
  testrx_MACDATA_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_8_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_8_OFF_RST,
      O => testrx_MACDATA_8_OBUF
    );
  MACDATA_8_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_8_OFF_RST
    );
  memcontroller_qn_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(10),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_10_IFF_RST,
      O => memcontroller_qn(10)
    );
  MD_10_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_10_IFF_RST
    );
  memcontroller_ts_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_31_TFF_RST,
      O => memcontroller_ts(31)
    );
  MD_31_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_31_TFF_RST
    );
  memcontroller_dnout_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_24_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_24_OFF_RST,
      O => memcontroller_dnout(24)
    );
  MD_24_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_24_OFF_RST
    );
  memcontroller_ts_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_24_TFF_RST,
      O => memcontroller_ts(24)
    );
  MD_24_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_24_TFF_RST
    );
  memcontroller_qn_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(16),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_16_IFF_RST,
      O => memcontroller_qn(16)
    );
  MD_16_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_16_IFF_RST
    );
  memcontroller_dnout_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_16_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_16_OFF_RST,
      O => memcontroller_dnout(16)
    );
  MD_16_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_16_OFF_RST
    );
  memcontroller_ts_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_16_TFF_RST,
      O => memcontroller_ts(16)
    );
  MD_16_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_16_TFF_RST
    );
  memcontroller_qn_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(17),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_17_IFF_RST,
      O => memcontroller_qn(17)
    );
  MD_17_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_17_IFF_RST
    );
  memcontroller_qn_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(25),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_25_IFF_RST,
      O => memcontroller_qn(25)
    );
  MD_25_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_25_IFF_RST
    );
  memcontroller_dnout_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_17_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_17_OFF_RST,
      O => memcontroller_dnout(17)
    );
  MD_17_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_17_OFF_RST
    );
  memcontroller_dnout_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_10_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_10_OFF_RST,
      O => memcontroller_dnout(10)
    );
  MD_10_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_10_OFF_RST
    );
  memcontroller_ts_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_10_TFF_RST,
      O => memcontroller_ts(10)
    );
  MD_10_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_10_TFF_RST
    );
  testrx_MACDATA_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_9_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_9_OFF_RST,
      O => testrx_MACDATA_9_OBUF
    );
  MACDATA_9_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_9_OFF_RST
    );
  memcontroller_qn_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(11),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_11_IFF_RST,
      O => memcontroller_qn(11)
    );
  MD_11_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_11_IFF_RST
    );
  memcontroller_dnout_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_11_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_11_OFF_RST,
      O => memcontroller_dnout(11)
    );
  MD_11_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_11_OFF_RST
    );
  memcontroller_ts_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_11_TFF_RST,
      O => memcontroller_ts(11)
    );
  MD_11_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_11_TFF_RST
    );
  memcontroller_qn_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(20),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_20_IFF_RST,
      O => memcontroller_qn(20)
    );
  MD_20_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_20_IFF_RST
    );
  memcontroller_qn_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(12),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_12_IFF_RST,
      O => memcontroller_qn(12)
    );
  MD_12_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_12_IFF_RST
    );
  memcontroller_dnout_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_20_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_20_OFF_RST,
      O => memcontroller_dnout(20)
    );
  MD_20_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_20_OFF_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_sin,
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => MDIO_IFF_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(0)
    );
  MDIO_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MDIO_IFF_RST
    );
  testrx_rxdl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_RXD_0_IBUF,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => RXD_0_IFF_RST,
      O => testrx_rxdl(0)
    );
  RXD_0_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_0_IFF_RST
    );
  testrx_rxdl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_RXD_1_IBUF,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => RXD_1_IFF_RST,
      O => testrx_rxdl(1)
    );
  RXD_1_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_1_IFF_RST
    );
  testrx_rxdl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_RXD_2_IBUF,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => RXD_2_IFF_RST,
      O => testrx_rxdl(2)
    );
  RXD_2_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_2_IFF_RST
    );
  testrx_rxdl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_RXD_3_IBUF,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => RXD_3_IFF_RST,
      O => testrx_rxdl(3)
    );
  RXD_3_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_3_IFF_RST
    );
  testrx_rxdl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_RXD_4_IBUF,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => RXD_4_IFF_RST,
      O => testrx_rxdl(4)
    );
  RXD_4_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_4_IFF_RST
    );
  testrx_rxdl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_RXD_5_IBUF,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => RXD_5_IFF_RST,
      O => testrx_rxdl(5)
    );
  RXD_5_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_5_IFF_RST
    );
  memcontroller_dnout_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_28_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_28_OFF_RST,
      O => memcontroller_dnout(28)
    );
  MD_28_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_28_OFF_RST
    );
  memcontroller_ts_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_28_TFF_RST,
      O => memcontroller_ts(28)
    );
  MD_28_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_28_TFF_RST
    );
  memcontroller_qn_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(29),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_29_IFF_RST,
      O => memcontroller_qn(29)
    );
  MD_29_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_29_IFF_RST
    );
  memcontroller_dnout_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_29_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_29_OFF_RST,
      O => memcontroller_dnout(29)
    );
  MD_29_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_29_OFF_RST
    );
  memcontroller_ts_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_29_TFF_RST,
      O => memcontroller_ts(29)
    );
  MD_29_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_29_TFF_RST
    );
  maccontrol_LED100 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LED100_OD,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => LED100_OFF_RST,
      O => maccontrol_LED100_OBUF
    );
  LED100_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LED100_OFF_RST
    );
  testrx_nextfl_754 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => NEXTF_IBUF_0,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => NEXTF_IFF_RST,
      O => testrx_nextfl
    );
  NEXTF_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => NEXTF_IFF_RST
    );
  memcontroller_ts_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_30_TFF_RST,
      O => memcontroller_ts(30)
    );
  MD_30_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_30_TFF_RST
    );
  memcontroller_dnout_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_23_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_23_OFF_RST,
      O => memcontroller_dnout(23)
    );
  MD_23_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_23_OFF_RST
    );
  memcontroller_ts_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_23_TFF_RST,
      O => memcontroller_ts(23)
    );
  MD_23_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_23_TFF_RST
    );
  memcontroller_qn_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(15),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_15_IFF_RST,
      O => memcontroller_qn(15)
    );
  MD_15_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_15_IFF_RST
    );
  memcontroller_dnout_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_15_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_15_OFF_RST,
      O => memcontroller_dnout(15)
    );
  MD_15_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_15_OFF_RST
    );
  memcontroller_ts_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_15_TFF_RST,
      O => memcontroller_ts(15)
    );
  MD_15_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_15_TFF_RST
    );
  memcontroller_qn_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(31),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_31_IFF_RST,
      O => memcontroller_qn(31)
    );
  MD_31_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_31_IFF_RST
    );
  memcontroller_qn_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(24),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_24_IFF_RST,
      O => memcontroller_qn(24)
    );
  MD_24_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_24_IFF_RST
    );
  memcontroller_dnout_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_31_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_31_OFF_RST,
      O => memcontroller_dnout(31)
    );
  MD_31_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_31_OFF_RST
    );
  memcontroller_we : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => MWE_OD,
      CE => MWE_OCEMUXNOT,
      CLK => clk,
      SET => MWE_OFF_SET,
      RST => GND,
      O => memcontroller_WEEXT
    );
  MWE_OFF_SETOR : X_BUF
    port map (
      I => GSR,
      O => MWE_OFF_SET
    );
  testrx_rxdl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_RXD_6_IBUF,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => RXD_6_IFF_RST,
      O => testrx_rxdl(6)
    );
  RXD_6_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_6_IFF_RST
    );
  testrx_rxdl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_RXD_7_IBUF,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => RXD_7_IFF_RST,
      O => testrx_rxdl(7)
    );
  RXD_7_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_7_IFF_RST
    );
  maccontrol_LED1000 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LED1000_OD,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => LED1000_OFF_RST,
      O => maccontrol_LED1000_OBUF
    );
  LED1000_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LED1000_OFF_RST
    );
  testrx_rx_dvl_755 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => RX_DV_IBUF_5,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => RX_DV_IFF_RST,
      O => testrx_rx_dvl
    );
  RX_DV_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RX_DV_IFF_RST
    );
  testrx_MACDATA_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_10_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_10_OFF_RST,
      O => testrx_MACDATA_10_OBUF
    );
  MACDATA_10_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_10_OFF_RST
    );
  memtest_datacnt_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(1),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_0_FFY_RST,
      O => d1(1)
    );
  d1_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_0_FFY_RST
    );
  memtest_datacnt_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(3),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_2_FFY_RST,
      O => d1(3)
    );
  d1_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_2_FFY_RST
    );
  memtest_datacnt_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_Madd_n0000_inst_lut2_38,
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_0_FFX_RST,
      O => d1(0)
    );
  d1_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_0_FFX_RST
    );
  memtest_datacnt_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(5),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_4_FFY_RST,
      O => d1(5)
    );
  d1_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_4_FFY_RST
    );
  maccontrol_ledtx_cnt_124_756 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_178,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_123_FFY_RST,
      O => maccontrol_ledtx_cnt_124
    );
  maccontrol_ledtx_cnt_123_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_123_FFY_RST
    );
  maccontrol_ledtx_cnt_126_757 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_180,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_125_FFY_RST,
      O => maccontrol_ledtx_cnt_126
    );
  maccontrol_ledtx_cnt_125_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_125_FFY_RST
    );
  maccontrol_ledtx_cnt_128_758 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_182,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_127_FFY_RST,
      O => maccontrol_ledtx_cnt_128
    );
  maccontrol_ledtx_cnt_127_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_127_FFY_RST
    );
  maccontrol_ledtx_cnt_123_759 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_lut3_155,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_123_FFX_RST,
      O => maccontrol_ledtx_cnt_123
    );
  maccontrol_ledtx_cnt_123_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_123_FFX_RST
    );
  testrx_MACDATA_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_11_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_11_OFF_RST,
      O => testrx_MACDATA_11_OBUF
    );
  MACDATA_11_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_11_OFF_RST
    );
  testrx_MACDATA_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_12_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_12_OFF_RST,
      O => testrx_MACDATA_12_OBUF
    );
  MACDATA_12_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_12_OFF_RST
    );
  testrx_MACDATA_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_13_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_13_OFF_RST,
      O => testrx_MACDATA_13_OBUF
    );
  MACDATA_13_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_13_OFF_RST
    );
  testrx_MACDATA_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_14_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_14_OFF_RST,
      O => testrx_MACDATA_14_OBUF
    );
  MACDATA_14_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_14_OFF_RST
    );
  maccontrol_ledtx_cnt_125_760 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_179,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_125_FFX_RST,
      O => maccontrol_ledtx_cnt_125
    );
  maccontrol_ledtx_cnt_125_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_125_FFX_RST
    );
  maccontrol_ledtx_cnt_127_761 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_181,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_127_FFX_RST,
      O => maccontrol_ledtx_cnt_127
    );
  maccontrol_ledtx_cnt_127_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_127_FFX_RST
    );
  maccontrol_ledtx_cnt_130_762 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_184,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_129_FFY_RST,
      O => maccontrol_ledtx_cnt_130
    );
  maccontrol_ledtx_cnt_129_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_129_FFY_RST
    );
  maccontrol_ledtx_cnt_129_763 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_183,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_129_FFX_RST,
      O => maccontrol_ledtx_cnt_129
    );
  maccontrol_ledtx_cnt_129_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_129_FFX_RST
    );
  maccontrol_ledtx_cnt_132_764 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_186,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_131_FFY_RST,
      O => maccontrol_ledtx_cnt_132
    );
  maccontrol_ledtx_cnt_131_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_131_FFY_RST
    );
  maccontrol_bitcnt_86_765 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_bitcnt_inst_sum_140,
      CE => maccontrol_n0022,
      CLK => clk,
      SET => GND,
      RST => maccontrol_bitcnt_86_FFX_RST,
      O => maccontrol_bitcnt_86
    );
  maccontrol_bitcnt_86_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_bitcnt_86_FFX_RST
    );
  maccontrol_bitcnt_89_766 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_bitcnt_inst_sum_143,
      CE => maccontrol_n0022,
      CLK => clk,
      SET => GND,
      RST => maccontrol_bitcnt_88_FFY_RST,
      O => maccontrol_bitcnt_89
    );
  maccontrol_bitcnt_88_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_bitcnt_88_FFY_RST
    );
  maccontrol_phyrstcnt_91_767 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_145,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_91_FFY_RST,
      O => maccontrol_phyrstcnt_91
    );
  maccontrol_phyrstcnt_91_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_91_FFY_RST
    );
  maccontrol_bitcnt_90_768 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_bitcnt_inst_sum_144,
      CE => maccontrol_n0022,
      CLK => clk,
      SET => GND,
      RST => maccontrol_bitcnt_90_FFX_RST,
      O => maccontrol_bitcnt_90
    );
  maccontrol_bitcnt_90_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_bitcnt_90_FFX_RST
    );
  maccontrol_bitcnt_88_769 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_bitcnt_inst_sum_142,
      CE => maccontrol_n0022,
      CLK => clk,
      SET => GND,
      RST => maccontrol_bitcnt_88_FFX_RST,
      O => maccontrol_bitcnt_88
    );
  maccontrol_bitcnt_88_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_bitcnt_88_FFX_RST
    );
  maccontrol_phyrstcnt_93_770 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_147,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_92_FFY_RST,
      O => maccontrol_phyrstcnt_93
    );
  maccontrol_phyrstcnt_92_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_92_FFY_RST
    );
  memcontroller_ts_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_26_TFF_RST,
      O => memcontroller_ts(26)
    );
  MD_26_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_26_TFF_RST
    );
  memcontroller_dnout_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_19_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_19_OFF_RST,
      O => memcontroller_dnout(19)
    );
  MD_19_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_19_OFF_RST
    );
  memcontroller_ts_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_19_TFF_RST,
      O => memcontroller_ts(19)
    );
  MD_19_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_19_TFF_RST
    );
  memcontroller_qn_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(27),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_27_IFF_RST,
      O => memcontroller_qn(27)
    );
  MD_27_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_27_IFF_RST
    );
  memcontroller_dnout_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_27_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_27_OFF_RST,
      O => memcontroller_dnout(27)
    );
  MD_27_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_27_OFF_RST
    );
  memcontroller_ts_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_27_TFF_RST,
      O => memcontroller_ts(27)
    );
  MD_27_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_27_TFF_RST
    );
  maccontrol_PHYRESET : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => PHYRESET_OD,
      CE => maccontrol_n0040,
      CLK => clk,
      SET => GND,
      RST => PHYRESET_OFF_RST,
      O => maccontrol_PHYRESET_OBUF
    );
  PHYRESET_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => PHYRESET_OFF_RST
    );
  memcontroller_qn_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(28),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_28_IFF_RST,
      O => memcontroller_qn(28)
    );
  MD_28_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_28_IFF_RST
    );
  memcontroller_ts_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_13_TFF_RST,
      O => memcontroller_ts(13)
    );
  MD_13_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_13_TFF_RST
    );
  memcontroller_dnout_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_22_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_22_OFF_RST,
      O => memcontroller_dnout(22)
    );
  MD_22_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_22_OFF_RST
    );
  memcontroller_ts_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_22_TFF_RST,
      O => memcontroller_ts(22)
    );
  MD_22_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_22_TFF_RST
    );
  memcontroller_qn_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(14),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_14_IFF_RST,
      O => memcontroller_qn(14)
    );
  MD_14_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_14_IFF_RST
    );
  memcontroller_dnout_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_14_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_14_OFF_RST,
      O => memcontroller_dnout(14)
    );
  MD_14_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_14_OFF_RST
    );
  memcontroller_ts_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_14_TFF_RST,
      O => memcontroller_ts(14)
    );
  MD_14_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_14_TFF_RST
    );
  memcontroller_qn_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(30),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_30_IFF_RST,
      O => memcontroller_qn(30)
    );
  MD_30_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_30_IFF_RST
    );
  memcontroller_qn_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(23),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_23_IFF_RST,
      O => memcontroller_qn(23)
    );
  MD_23_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_23_IFF_RST
    );
  memcontroller_dnout_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_30_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_30_OFF_RST,
      O => memcontroller_dnout(30)
    );
  MD_30_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_30_OFF_RST
    );
  cnt_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(2),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_2_FFX_RST,
      O => cnt(2)
    );
  cnt_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_2_FFX_RST
    );
  cnt_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(5),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_4_FFY_RST,
      O => cnt(5)
    );
  cnt_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_4_FFY_RST
    );
  cnt_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(9),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_8_FFY_RST,
      O => cnt(9)
    );
  cnt_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_8_FFY_RST
    );
  cnt_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(4),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_4_FFX_RST,
      O => cnt(4)
    );
  cnt_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_4_FFX_RST
    );
  cnt_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(7),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_6_FFY_RST,
      O => cnt(7)
    );
  cnt_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_6_FFY_RST
    );
  memcontroller_ts_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_20_TFF_RST,
      O => memcontroller_ts(20)
    );
  MD_20_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_20_TFF_RST
    );
  memcontroller_dnout_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_12_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_12_OFF_RST,
      O => memcontroller_dnout(12)
    );
  MD_12_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_12_OFF_RST
    );
  memcontroller_ts_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_12_TFF_RST,
      O => memcontroller_ts(12)
    );
  MD_12_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_12_TFF_RST
    );
  memcontroller_qn_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(21),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_21_IFF_RST,
      O => memcontroller_qn(21)
    );
  MD_21_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_21_IFF_RST
    );
  memcontroller_dnout_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_21_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_21_OFF_RST,
      O => memcontroller_dnout(21)
    );
  MD_21_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_21_OFF_RST
    );
  memcontroller_ts_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_21_TFF_RST,
      O => memcontroller_ts(21)
    );
  MD_21_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_21_TFF_RST
    );
  memcontroller_qn_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(13),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_13_IFF_RST,
      O => memcontroller_qn(13)
    );
  MD_13_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_13_IFF_RST
    );
  memcontroller_qn_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(22),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_22_IFF_RST,
      O => memcontroller_qn(22)
    );
  MD_22_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_22_IFF_RST
    );
  memcontroller_dnout_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_13_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_13_OFF_RST,
      O => memcontroller_dnout(13)
    );
  MD_13_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_13_OFF_RST
    );
  testrx_addr_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_addr_n0000(7),
      CE => testrx_cs_FFd2,
      CLK => rx_clk_int,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => testrx_n0008,
      O => testrx_addr(7)
    );
  testrx_addr_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_addr_n0000(2),
      CE => testrx_cs_FFd2,
      CLK => rx_clk_int,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => testrx_n0008,
      O => testrx_addr(2)
    );
  testrx_addr_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_addr_n0000(4),
      CE => testrx_cs_FFd2,
      CLK => rx_clk_int,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => testrx_n0008,
      O => testrx_addr(4)
    );
  testrx_addr_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_addr_n0000(6),
      CE => testrx_cs_FFd2,
      CLK => rx_clk_int,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => testrx_n0008,
      O => testrx_addr(6)
    );
  memtest2_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(1),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(1)
    );
  memtest2_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(3),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(3)
    );
  cnt_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(6),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_6_FFX_RST,
      O => cnt(6)
    );
  cnt_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_6_FFX_RST
    );
  cnt_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(8),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_8_FFX_RST,
      O => cnt(8)
    );
  cnt_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_8_FFX_RST
    );
  cnt_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(11),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_10_FFY_RST,
      O => cnt(11)
    );
  cnt_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_10_FFY_RST
    );
  cnt_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(15),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_14_FFY_RST,
      O => cnt(15)
    );
  cnt_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_14_FFY_RST
    );
  cnt_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(10),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_10_FFX_RST,
      O => cnt(10)
    );
  cnt_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_10_FFX_RST
    );
  cnt_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(13),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_12_FFY_RST,
      O => cnt(13)
    );
  cnt_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_12_FFY_RST
    );
  memcontroller_ts_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_17_TFF_RST,
      O => memcontroller_ts(17)
    );
  MD_17_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_17_TFF_RST
    );
  memcontroller_dnout_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_25_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_25_OFF_RST,
      O => memcontroller_dnout(25)
    );
  MD_25_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_25_OFF_RST
    );
  memcontroller_ts_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_25_TFF_RST,
      O => memcontroller_ts(25)
    );
  MD_25_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_25_TFF_RST
    );
  memcontroller_qn_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(18),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_18_IFF_RST,
      O => memcontroller_qn(18)
    );
  MD_18_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_18_IFF_RST
    );
  memcontroller_dnout_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_18_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_18_OFF_RST,
      O => memcontroller_dnout(18)
    );
  MD_18_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_18_OFF_RST
    );
  memcontroller_ts_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_18_TFF_RST,
      O => memcontroller_ts(18)
    );
  MD_18_TFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_18_TFF_RST
    );
  memcontroller_qn_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(26),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_26_IFF_RST,
      O => memcontroller_qn(26)
    );
  MD_26_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_26_IFF_RST
    );
  memcontroller_qn_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(19),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_19_IFF_RST,
      O => memcontroller_qn(19)
    );
  MD_19_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_19_IFF_RST
    );
  memcontroller_dnout_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_26_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => MD_26_OFF_RST,
      O => memcontroller_dnout(26)
    );
  MD_26_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_26_OFF_RST
    );
  maccontrol_phyrstcnt_110_771 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_164,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_110_FFX_RST,
      O => maccontrol_phyrstcnt_110
    );
  maccontrol_phyrstcnt_110_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_110_FFX_RST
    );
  maccontrol_phyrstcnt_113_772 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_167,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_112_FFY_RST,
      O => maccontrol_phyrstcnt_113
    );
  maccontrol_phyrstcnt_112_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_112_FFY_RST
    );
  maccontrol_phyrstcnt_117_773 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_171,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_116_FFY_RST,
      O => maccontrol_phyrstcnt_117
    );
  maccontrol_phyrstcnt_116_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_116_FFY_RST
    );
  maccontrol_phyrstcnt_112_774 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_166,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_112_FFX_RST,
      O => maccontrol_phyrstcnt_112
    );
  maccontrol_phyrstcnt_112_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_112_FFX_RST
    );
  maccontrol_phyrstcnt_115_775 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_169,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_114_FFY_RST,
      O => maccontrol_phyrstcnt_115
    );
  maccontrol_phyrstcnt_114_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_114_FFY_RST
    );
  maccontrol_phyrstcnt_114_776 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_168,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_114_FFX_RST,
      O => maccontrol_phyrstcnt_114
    );
  maccontrol_phyrstcnt_114_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_114_FFX_RST
    );
  testrx_MACDATA_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MACDATA_15_OD,
      CE => VCC,
      CLK => ifclk_int,
      SET => GND,
      RST => MACDATA_15_OFF_RST,
      O => testrx_MACDATA_15_OBUF
    );
  MACDATA_15_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MACDATA_15_OFF_RST
    );
  maccontrol_LEDTX : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDTX_OD,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => LEDTX_OFF_RST,
      O => maccontrol_LEDTX_OBUF
    );
  LEDTX_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDTX_OFF_RST
    );
  LEDPOWER_777 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDPOWER_OD,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => LEDPOWER_OFF_RST,
      O => LEDPOWER_OBUF
    );
  LEDPOWER_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDPOWER_OFF_RST
    );
  maccontrol_phyrstcnt_96_778 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_150,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_96_FFX_RST,
      O => maccontrol_phyrstcnt_96
    );
  maccontrol_phyrstcnt_96_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_96_FFX_RST
    );
  maccontrol_phyrstcnt_98_779 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_152,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_98_FFX_RST,
      O => maccontrol_phyrstcnt_98
    );
  maccontrol_phyrstcnt_98_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_98_FFX_RST
    );
  maccontrol_phyrstcnt_101_780 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_155,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_100_FFY_RST,
      O => maccontrol_phyrstcnt_101
    );
  maccontrol_phyrstcnt_100_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_100_FFY_RST
    );
  maccontrol_phyrstcnt_103_781 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_157,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_102_FFY_RST,
      O => maccontrol_phyrstcnt_103
    );
  maccontrol_phyrstcnt_102_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_102_FFY_RST
    );
  maccontrol_phyrstcnt_100_782 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_154,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_100_FFX_RST,
      O => maccontrol_phyrstcnt_100
    );
  maccontrol_phyrstcnt_100_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_100_FFX_RST
    );
  maccontrol_phyrstcnt_105_783 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_159,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_104_FFY_RST,
      O => maccontrol_phyrstcnt_105
    );
  maccontrol_phyrstcnt_104_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_104_FFY_RST
    );
  maccontrol_ledtx_cnt_131_784 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_185,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_131_FFX_RST,
      O => maccontrol_ledtx_cnt_131
    );
  maccontrol_ledtx_cnt_131_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_131_FFX_RST
    );
  maccontrol_ledtx_cnt_134_785 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_188,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_133_FFY_RST,
      O => maccontrol_ledtx_cnt_134
    );
  maccontrol_ledtx_cnt_133_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_133_FFY_RST
    );
  maccontrol_bitcnt_87_786 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_bitcnt_inst_sum_141,
      CE => maccontrol_n0022,
      CLK => clk,
      SET => GND,
      RST => maccontrol_bitcnt_86_FFY_RST,
      O => maccontrol_bitcnt_87
    );
  maccontrol_bitcnt_86_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_bitcnt_86_FFY_RST
    );
  maccontrol_ledtx_cnt_133_787 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_ledtx_cnt_inst_sum_187,
      CE => maccontrol_n0044,
      CLK => clk,
      SET => GND,
      RST => maccontrol_ledtx_cnt_133_FFX_RST,
      O => maccontrol_ledtx_cnt_133
    );
  maccontrol_ledtx_cnt_133_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_ledtx_cnt_133_FFX_RST
    );
  maccontrol_bitcnt_85_788 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_bitcnt_inst_sum_139,
      CE => maccontrol_n0022,
      CLK => clk,
      SET => GND,
      RST => maccontrol_bitcnt_85_FFY_RST,
      O => maccontrol_bitcnt_85
    );
  maccontrol_bitcnt_85_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_bitcnt_85_FFY_RST
    );
  memtest_Mshreg_dataw4_27_10_789 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_27_net9,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_27_10_FFY_RST,
      O => memtest_Mshreg_dataw4_27_10
    );
  memtest_Mshreg_dataw4_27_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_27_10_FFY_RST
    );
  memcontroller_oe_790 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_wen,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memcontroller_oe_FFY_RST,
      O => memcontroller_oe
    );
  memcontroller_oe_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_oe_FFY_RST
    );
  memtest_Mshreg_dataw4_19_18_791 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_19_net25,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_19_18_FFY_RST,
      O => memtest_Mshreg_dataw4_19_18
    );
  memtest_Mshreg_dataw4_19_18_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_19_18_FFY_RST
    );
  maccontrol_sclkdelta_792 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_lsclkdelta,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => maccontrol_sclkdelta_FFY_RST,
      O => maccontrol_sclkdelta
    );
  maccontrol_sclkdelta_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_sclkdelta_FFY_RST
    );
  memtest_Mshreg_dataw4_30_7_793 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_30_net3,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_30_7_FFY_RST,
      O => memtest_Mshreg_dataw4_30_7
    );
  memtest_Mshreg_dataw4_30_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_30_7_FFY_RST
    );
  memtest2_addrlfsr_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(0),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(1)
    );
  memtest2_addrlfsr_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_n0150,
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(0)
    );
  memtest_Mshreg_dataw4_0_37_794 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_0_net63,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_0_37_FFY_RST,
      O => memtest_Mshreg_dataw4_0_37
    );
  memtest_Mshreg_dataw4_0_37_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_0_37_FFY_RST
    );
  memtest_Mshreg_dataw4_28_9_795 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_28_net7,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_28_9_FFY_RST,
      O => memtest_Mshreg_dataw4_28_9
    );
  memtest_Mshreg_dataw4_28_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_28_9_FFY_RST
    );
  memtest_Mshreg_dataw4_29_8_796 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_29_net5,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_29_8_FFY_RST,
      O => memtest_Mshreg_dataw4_29_8
    );
  memtest_Mshreg_dataw4_29_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_29_8_FFY_RST
    );
  maccontrol_phyrstcnt_92_797 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_146,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_92_FFX_RST,
      O => maccontrol_phyrstcnt_92
    );
  maccontrol_phyrstcnt_92_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_92_FFX_RST
    );
  maccontrol_phyrstcnt_95_798 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_149,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_94_FFY_RST,
      O => maccontrol_phyrstcnt_95
    );
  maccontrol_phyrstcnt_94_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_94_FFY_RST
    );
  maccontrol_phyrstcnt_94_799 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_148,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_94_FFX_RST,
      O => maccontrol_phyrstcnt_94
    );
  maccontrol_phyrstcnt_94_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_94_FFX_RST
    );
  maccontrol_phyrstcnt_97_800 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_151,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_96_FFY_RST,
      O => maccontrol_phyrstcnt_97
    );
  maccontrol_phyrstcnt_96_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_96_FFY_RST
    );
  maccontrol_phyrstcnt_99_801 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_153,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_98_FFY_RST,
      O => maccontrol_phyrstcnt_99
    );
  maccontrol_phyrstcnt_98_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_98_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_124,
      CE => maccontrol_PHY_status_MII_Interface_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_mdccnt_3_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_mdccnt(3)
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_3_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_126,
      CE => maccontrol_PHY_status_MII_Interface_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_mdccnt_5_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_mdccnt(5)
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_5_FFX_RST
    );
  maccontrol_phyrstcnt_102_802 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_156,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_102_FFX_RST,
      O => maccontrol_phyrstcnt_102
    );
  maccontrol_phyrstcnt_102_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_102_FFX_RST
    );
  maccontrol_phyrstcnt_104_803 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_158,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_104_FFX_RST,
      O => maccontrol_phyrstcnt_104
    );
  maccontrol_phyrstcnt_104_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_104_FFX_RST
    );
  maccontrol_phyrstcnt_107_804 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_161,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_106_FFY_RST,
      O => maccontrol_phyrstcnt_107
    );
  maccontrol_phyrstcnt_106_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_106_FFY_RST
    );
  maccontrol_phyrstcnt_106_805 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_160,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_106_FFX_RST,
      O => maccontrol_phyrstcnt_106
    );
  maccontrol_phyrstcnt_106_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_106_FFX_RST
    );
  maccontrol_phyrstcnt_109_806 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_163,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_108_FFY_RST,
      O => maccontrol_phyrstcnt_109
    );
  maccontrol_phyrstcnt_108_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_108_FFY_RST
    );
  maccontrol_phyrstcnt_108_807 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_162,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_108_FFX_RST,
      O => maccontrol_phyrstcnt_108
    );
  maccontrol_phyrstcnt_108_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_108_FFX_RST
    );
  maccontrol_phyrstcnt_111_808 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_165,
      CE => maccontrol_n0039,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_110_FFY_RST,
      O => maccontrol_phyrstcnt_111
    );
  maccontrol_phyrstcnt_110_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_110_FFY_RST
    );
  cnt0_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => cnt0_n0000(4),
      CE => Q_n0034,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => err,
      O => cnt0(4)
    );
  cnt_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(1),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_0_FFY_RST,
      O => cnt(1)
    );
  cnt_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_0_FFY_RST
    );
  cnt_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Madd_n0000_inst_lut2_0,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_0_FFX_RST,
      O => cnt(0)
    );
  cnt_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_0_FFX_RST
    );
  cnt_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(3),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_2_FFY_RST,
      O => cnt(3)
    );
  cnt_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_2_FFY_RST
    );
  cnt_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(12),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_12_FFX_RST,
      O => cnt(12)
    );
  cnt_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_12_FFX_RST
    );
  cnt_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(14),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_14_FFX_RST,
      O => cnt(14)
    );
  cnt_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_14_FFX_RST
    );
  cnt_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(17),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_16_FFY_RST,
      O => cnt(17)
    );
  cnt_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_16_FFY_RST
    );
  cnt_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(16),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_16_FFX_RST,
      O => cnt(16)
    );
  cnt_16_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_16_FFX_RST
    );
  cnt_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(19),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_18_FFY_RST,
      O => cnt(19)
    );
  cnt_18_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_18_FFY_RST
    );
  memtest_datacnt_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(8),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_8_FFX_RST,
      O => d1(8)
    );
  d1_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_8_FFX_RST
    );
  memtest_datacnt_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(10),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_10_FFX_RST,
      O => d1(10)
    );
  d1_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_10_FFX_RST
    );
  memtest_datacnt_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(13),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_12_FFY_RST,
      O => d1(13)
    );
  d1_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_12_FFY_RST
    );
  memtest_datacnt_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(12),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_12_FFX_RST,
      O => d1(12)
    );
  d1_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_12_FFX_RST
    );
  memtest_datacnt_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(15),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_14_FFY_RST,
      O => d1(15)
    );
  d1_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_14_FFY_RST
    );
  maccontrol_phyrstcnt_120_809 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_174,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_120_FFX_RST,
      O => maccontrol_phyrstcnt_120
    );
  maccontrol_phyrstcnt_120_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_120_FFX_RST
    );
  maccontrol_phyrstcnt_122_810 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_176,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_122_FFX_RST,
      O => maccontrol_phyrstcnt_122
    );
  maccontrol_phyrstcnt_122_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_122_FFX_RST
    );
  cnt0_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => cnt0_n0000(1),
      CE => Q_n0034,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => err,
      O => cnt0(1)
    );
  cnt0_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => cnt0_Madd_n0000_inst_lut2_24,
      CE => Q_n0034,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => err,
      O => cnt0(0)
    );
  cnt0_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => cnt0_n0000(2),
      CE => Q_n0034,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => err,
      O => cnt0(2)
    );
  cnt0_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => cnt0_n0000(5),
      CE => Q_n0034,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => err,
      O => cnt0(5)
    );
  maccontrol_phyrstcnt_116_811 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_170,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_116_FFX_RST,
      O => maccontrol_phyrstcnt_116
    );
  maccontrol_phyrstcnt_116_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_116_FFX_RST
    );
  maccontrol_phyrstcnt_119_812 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_173,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_118_FFY_RST,
      O => maccontrol_phyrstcnt_119
    );
  maccontrol_phyrstcnt_118_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_118_FFY_RST
    );
  maccontrol_phyrstcnt_118_813 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_172,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_118_FFX_RST,
      O => maccontrol_phyrstcnt_118
    );
  maccontrol_phyrstcnt_118_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_118_FFX_RST
    );
  maccontrol_phyrstcnt_121_814 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyrstcnt_inst_sum_175,
      CE => maccontrol_n0039124_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyrstcnt_120_FFY_RST,
      O => maccontrol_phyrstcnt_121
    );
  maccontrol_phyrstcnt_120_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyrstcnt_120_FFY_RST
    );
  txsim_counter_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(14),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(14)
    );
  txsim_counter_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(16),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(16)
    );
  testrx_addr_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_addr_n0000(3),
      CE => testrx_cs_FFd2,
      CLK => rx_clk_int,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => testrx_n0008,
      O => testrx_addr(3)
    );
  testrx_addr_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_addr_n0000(1),
      CE => testrx_cs_FFd2,
      CLK => rx_clk_int,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => testrx_n0008,
      O => testrx_addr(1)
    );
  testrx_addr_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_addr_Madd_n0000_inst_lut2_30,
      CE => testrx_cs_FFd2,
      CLK => rx_clk_int,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => testrx_n0008,
      O => testrx_addr(0)
    );
  testrx_addr_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_addr_n0000(5),
      CE => testrx_cs_FFd2,
      CLK => rx_clk_int,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => testrx_n0008,
      O => testrx_addr(5)
    );
  txsim_counter_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(1),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(1)
    );
  txsim_counter_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(3),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(3)
    );
  txsim_counter_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_Madd_n0000_inst_lut2_103,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(0)
    );
  txsim_counter_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(5),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(5)
    );
  txsim_counter_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(2),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(2)
    );
  txsim_counter_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(4),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(4)
    );
  txsim_counter_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(7),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(7)
    );
  txsim_counter_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(11),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(11)
    );
  txsim_counter_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(6),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(6)
    );
  txsim_counter_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(9),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(9)
    );
  memtest_datacnt_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(18),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_18_FFX_RST,
      O => d1(18)
    );
  d1_18_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_18_FFX_RST
    );
  memtest_datacnt_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(20),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_20_FFX_RST,
      O => d1(20)
    );
  d1_20_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_20_FFX_RST
    );
  memtest_datacnt_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(23),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_22_FFY_RST,
      O => d1(23)
    );
  d1_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_22_FFY_RST
    );
  memtest_datacnt_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(27),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_26_FFY_RST,
      O => d1(27)
    );
  d1_26_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_26_FFY_RST
    );
  memtest_datacnt_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(22),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_22_FFX_RST,
      O => d1(22)
    );
  d1_22_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_22_FFX_RST
    );
  memtest_datacnt_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(25),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_24_FFY_RST,
      O => d1(25)
    );
  d1_24_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_24_FFY_RST
    );
  memtest_datacnt_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(2),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_2_FFX_RST,
      O => d1(2)
    );
  d1_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_2_FFX_RST
    );
  memtest_datacnt_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(4),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_4_FFX_RST,
      O => d1(4)
    );
  d1_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_4_FFX_RST
    );
  memtest_datacnt_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(7),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_6_FFY_RST,
      O => d1(7)
    );
  d1_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_6_FFY_RST
    );
  memtest_datacnt_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(11),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_10_FFY_RST,
      O => d1(11)
    );
  d1_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_10_FFY_RST
    );
  memtest_datacnt_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(6),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_6_FFX_RST,
      O => d1(6)
    );
  d1_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_6_FFX_RST
    );
  memtest_datacnt_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(9),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_8_FFY_RST,
      O => d1(9)
    );
  d1_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_8_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_122,
      CE => maccontrol_PHY_status_MII_Interface_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_mdccnt_1_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_mdccnt(1)
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_1_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_125,
      CE => maccontrol_PHY_status_MII_Interface_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_mdccnt_3_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_mdccnt(4)
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_3_FFY_RST
    );
  cnt_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(18),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_18_FFX_RST,
      O => cnt(18)
    );
  cnt_18_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_18_FFX_RST
    );
  cnt_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(21),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_20_FFY_RST,
      O => cnt(21)
    );
  cnt_20_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_20_FFY_RST
    );
  cnt_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(20),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_20_FFX_RST,
      O => cnt(20)
    );
  cnt_20_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_20_FFX_RST
    );
  cnt_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => cnt_22_XORG,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_22_FFY_RST,
      O => cnt(23)
    );
  cnt_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_22_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_mdccnt_inst_sum_121,
      CE => maccontrol_PHY_status_MII_Interface_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_mdccnt_0_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_mdccnt(0)
    );
  maccontrol_PHY_status_MII_Interface_mdccnt_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_mdccnt_0_FFY_RST
    );
  cnt_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => Q_n0000(22),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => cnt_22_FFX_RST,
      O => cnt(22)
    );
  cnt_22_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => cnt_22_FFX_RST
    );
  memtest2_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(12),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(12)
    );
  memtest2_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(16),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(16)
    );
  memtest2_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(14),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(14)
    );
  memtest2_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_Madd_n0000_inst_lut2_86,
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(0)
    );
  memtest2_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(5),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(5)
    );
  memtest2_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(2),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(2)
    );
  memtest2_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(9),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(9)
    );
  memtest2_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(4),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(4)
    );
  memtest2_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(7),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(7)
    );
  memtest2_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(11),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(11)
    );
  memtest2_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(6),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(6)
    );
  memtest2_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(8),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(8)
    );
  memtest2_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(15),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(15)
    );
  memtest2_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(10),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(10)
    );
  memtest2_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cnt_n0000(13),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_n0011,
      O => memtest2_cnt(13)
    );
  txsim_counter_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(8),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(8)
    );
  txsim_counter_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(10),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(10)
    );
  txsim_counter_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(13),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(13)
    );
  txsim_counter_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(17),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(17)
    );
  txsim_counter_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(12),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(12)
    );
  txsim_counter_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_counter_n0000(15),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => txsim_SF22758,
      O => txsim_counter(15)
    );
  memtest_datacnt_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(14),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_14_FFX_RST,
      O => d1(14)
    );
  d1_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_14_FFX_RST
    );
  memtest_datacnt_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(17),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_16_FFY_RST,
      O => d1(17)
    );
  d1_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_16_FFY_RST
    );
  memtest_datacnt_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(21),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_20_FFY_RST,
      O => d1(21)
    );
  d1_20_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_20_FFY_RST
    );
  memtest_datacnt_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(16),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_16_FFX_RST,
      O => d1(16)
    );
  d1_16_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_16_FFX_RST
    );
  memtest_datacnt_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(19),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_18_FFY_RST,
      O => d1(19)
    );
  d1_18_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_18_FFY_RST
    );
  memtest_datacnt_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(30),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_30_FFX_RST,
      O => d1(30)
    );
  d1_30_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_30_FFX_RST
    );
  memtest_addrcnt_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(1),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_0_FFY_RST,
      O => addr1(1)
    );
  addr1_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_0_FFY_RST
    );
  memtest_addrcnt_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(5),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_4_FFY_RST,
      O => addr1(5)
    );
  addr1_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_4_FFY_RST
    );
  memtest_addrcnt_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_Madd_n0000_inst_lut2_70,
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_0_FFX_RST,
      O => addr1(0)
    );
  addr1_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_0_FFX_RST
    );
  memtest_addrcnt_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(3),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_2_FFY_RST,
      O => addr1(3)
    );
  addr1_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_2_FFY_RST
    );
  maccontrol_dout_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_14_58_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_14_FFX_RST,
      O => maccontrol_dout(14)
    );
  maccontrol_dout_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_14_FFX_RST
    );
  maccontrol_dout_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_3_76_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_3_FFY_RST,
      O => maccontrol_dout(3)
    );
  maccontrol_dout_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_3_FFY_RST
    );
  maccontrol_dout_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_5_58_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_5_FFY_RST,
      O => maccontrol_dout(5)
    );
  maccontrol_dout_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_5_FFY_RST
    );
  maccontrol_dout_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_6_58_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_8_FFY_RST,
      O => maccontrol_dout(6)
    );
  maccontrol_dout_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_8_FFY_RST
    );
  maccontrol_dout_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_8_58_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_8_FFX_RST,
      O => maccontrol_dout(8)
    );
  maccontrol_dout_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_8_FFX_RST
    );
  memtest_addrcnt_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(8),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_8_FFX_RST,
      O => addr1(8)
    );
  addr1_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_8_FFX_RST
    );
  memtest_addrcnt_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(10),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_10_FFX_RST,
      O => addr1(10)
    );
  addr1_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_10_FFX_RST
    );
  memtest_addrcnt_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(13),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_12_FFY_RST,
      O => addr1(13)
    );
  addr1_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_12_FFY_RST
    );
  memtest_addrcnt_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(12),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_12_FFX_RST,
      O => addr1(12)
    );
  addr1_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_12_FFX_RST
    );
  memtest_addrcnt_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(15),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_14_FFY_RST,
      O => addr1(15)
    );
  addr1_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_14_FFY_RST
    );
  memtest_addrcnt_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(14),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_14_FFX_RST,
      O => addr1(14)
    );
  addr1_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_14_FFX_RST
    );
  memtest2_MA_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(12),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_13_FFY_RST,
      O => addr2(12)
    );
  addr2_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_13_FFY_RST
    );
  memtest2_MA_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(13),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_13_FFX_RST,
      O => addr2(13)
    );
  addr2_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_13_FFX_RST
    );
  memtest2_datain_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(11),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_11_FFX_RST,
      O => memtest2_datain(11)
    );
  memtest2_datain_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_11_FFX_RST
    );
  memtest2_datain_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(30),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_30_FFX_RST,
      O => memtest2_datain(30)
    );
  memtest2_datain_30_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_30_FFX_RST
    );
  maccontrol_dout_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_0_92_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_0_FFY_RST,
      O => maccontrol_dout(0)
    );
  maccontrol_dout_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_0_FFY_RST
    );
  maccontrol_dout_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_26_22_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_26_FFY_RST,
      O => maccontrol_dout(26)
    );
  maccontrol_dout_26_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_26_FFY_RST
    );
  maccontrol_dout_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_27_25_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_27_FFY_RST,
      O => maccontrol_dout(27)
    );
  maccontrol_dout_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_27_FFY_RST
    );
  maccontrol_dout_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_19_25_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_19_FFY_RST,
      O => maccontrol_dout(19)
    );
  maccontrol_dout_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_19_FFY_RST
    );
  maccontrol_dout_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_28_22_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_28_FFY_RST,
      O => maccontrol_dout(28)
    );
  maccontrol_dout_28_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_28_FFY_RST
    );
  maccontrol_dout_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_29_22_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_29_FFY_RST,
      O => maccontrol_dout(29)
    );
  maccontrol_dout_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_29_FFY_RST
    );
  maccontrol_lmacaddr_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(11),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_27_FFX_RST,
      O => maccontrol_lmacaddr(27)
    );
  maccontrol_lmacaddr_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_27_FFX_RST
    );
  memtest2_ldata_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(31),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_31_FFX_RST,
      O => memtest2_ldata(31)
    );
  memtest2_ldata_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_31_FFX_RST
    );
  memtest2_ldata_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(22),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_23_FFY_RST,
      O => memtest2_ldata(22)
    );
  memtest2_ldata_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_23_FFY_RST
    );
  memtest2_ldata_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(23),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_23_FFX_RST,
      O => memtest2_ldata(23)
    );
  memtest2_ldata_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_23_FFX_RST
    );
  memtest2_ldata_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(14),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_15_FFY_RST,
      O => memtest2_ldata(14)
    );
  memtest2_ldata_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_15_FFY_RST
    );
  memtest2_ldata_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(15),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_15_FFX_RST,
      O => memtest2_ldata(15)
    );
  memtest2_ldata_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_15_FFX_RST
    );
  maccontrol_lmacaddr_36 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(4),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_37_FFY_RST,
      O => maccontrol_lmacaddr(36)
    );
  maccontrol_lmacaddr_37_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_37_FFY_RST
    );
  maccontrol_lmacaddr_37 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(5),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_37_FFX_RST,
      O => maccontrol_lmacaddr(37)
    );
  maccontrol_lmacaddr_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_37_FFX_RST
    );
  maccontrol_lmacaddr_44 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(12),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_45_FFY_RST,
      O => maccontrol_lmacaddr(44)
    );
  maccontrol_lmacaddr_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_45_FFY_RST
    );
  maccontrol_lmacaddr_45 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(13),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_45_FFX_RST,
      O => maccontrol_lmacaddr(45)
    );
  maccontrol_lmacaddr_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_45_FFX_RST
    );
  maccontrol_lmacaddr_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(13),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_29_FFX_RST,
      O => maccontrol_lmacaddr(29)
    );
  maccontrol_lmacaddr_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_29_FFX_RST
    );
  memtest2_ldata_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(24),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_25_FFY_RST,
      O => memtest2_ldata(24)
    );
  memtest2_ldata_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_25_FFY_RST
    );
  memtest2_ldata_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(25),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_25_FFX_RST,
      O => memtest2_ldata(25)
    );
  memtest2_ldata_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_25_FFX_RST
    );
  memtest2_ldata_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(16),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_17_FFY_RST,
      O => memtest2_ldata(16)
    );
  memtest2_ldata_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_17_FFY_RST
    );
  maccontrol_lmacaddr_38 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(6),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_39_FFY_RST,
      O => maccontrol_lmacaddr(38)
    );
  maccontrol_lmacaddr_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_39_FFY_RST
    );
  memtest2_Mshreg_data4_30_39_815 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_30_net67,
      CE => memtest2_n00511_1,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_30_39_FFY_RST,
      O => memtest2_Mshreg_data4_30_39
    );
  memtest2_Mshreg_data4_30_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_30_39_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd4_816 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_cs_FFd4_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_cs_FFd5_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd4
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd5_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd5_817 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_cs_FFd5_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_cs_FFd5_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd5
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd5_FFX_RST
    );
  memtest_Mshreg_dataw4_9_28_818 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_9_net45,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_9_28_FFY_RST,
      O => memtest_Mshreg_dataw4_9_28
    );
  memtest_Mshreg_dataw4_9_28_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_9_28_FFY_RST
    );
  memtest2_Mshreg_data4_15_54_819 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_15_net97,
      CE => memtest2_n00511_3,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_15_54_FFY_RST,
      O => memtest2_Mshreg_data4_15_54
    );
  memtest2_Mshreg_data4_15_54_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_15_54_FFY_RST
    );
  memtest2_Mshreg_data4_23_46_820 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_23_net81,
      CE => memtest2_n00511_2,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_23_46_FFY_RST,
      O => memtest2_Mshreg_data4_23_46
    );
  memtest2_Mshreg_data4_23_46_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_23_46_FFY_RST
    );
  memtest2_Mshreg_data4_31_38_821 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_31_net65,
      CE => memtest2_n00511_1,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_31_38_FFY_RST,
      O => memtest2_Mshreg_data4_31_38
    );
  memtest2_Mshreg_data4_31_38_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_31_38_FFY_RST
    );
  memtest2_Mshreg_data4_16_53_822 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_16_net95,
      CE => memtest2_n00511_3,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_16_53_FFY_RST,
      O => memtest2_Mshreg_data4_16_53
    );
  memtest2_Mshreg_data4_16_53_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_16_53_FFY_RST
    );
  memtest2_Mshreg_data4_18_51_823 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_18_net91,
      CE => memtest2_n00511_3,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_18_51_FFY_RST,
      O => memtest2_Mshreg_data4_18_51
    );
  memtest2_Mshreg_data4_18_51_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_18_51_FFY_RST
    );
  memtest2_Mshreg_data4_17_52_824 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_17_net93,
      CE => memtest2_n00511_3,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_17_52_FFY_RST,
      O => memtest2_Mshreg_data4_17_52
    );
  memtest2_Mshreg_data4_17_52_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_17_52_FFY_RST
    );
  memtest2_Mshreg_data4_25_44_825 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_25_net77,
      CE => memtest2_n00511_2,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_25_44_FFY_RST,
      O => memtest2_Mshreg_data4_25_44
    );
  memtest2_Mshreg_data4_25_44_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_25_44_FFY_RST
    );
  memtest_datacnt_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(24),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_24_FFX_RST,
      O => d1(24)
    );
  d1_24_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_24_FFX_RST
    );
  memtest_datacnt_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(31),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_30_FFY_RST,
      O => d1(31)
    );
  d1_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_30_FFY_RST
    );
  memtest_datacnt_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(26),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_26_FFX_RST,
      O => d1(26)
    );
  d1_26_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_26_FFX_RST
    );
  memtest_datacnt_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(29),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_28_FFY_RST,
      O => d1(29)
    );
  d1_28_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_28_FFY_RST
    );
  memtest_datacnt_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_datacnt_n0000(28),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => d1_28_FFX_RST,
      O => d1(28)
    );
  d1_28_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d1_28_FFX_RST
    );
  memtest_Mshreg_dataw4_1_36_826 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_1_net61,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_1_36_FFY_RST,
      O => memtest_Mshreg_dataw4_1_36
    );
  memtest_Mshreg_dataw4_1_36_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_1_36_FFY_RST
    );
  memtest_Mshreg_dataw4_2_35_827 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_2_net59,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_2_35_FFY_RST,
      O => memtest_Mshreg_dataw4_2_35
    );
  memtest_Mshreg_dataw4_2_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_2_35_FFY_RST
    );
  memtest_Mshreg_dataw4_3_34_828 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_3_net57,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_3_34_FFY_RST,
      O => memtest_Mshreg_dataw4_3_34
    );
  memtest_Mshreg_dataw4_3_34_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_3_34_FFY_RST
    );
  memtest2_MA_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(14),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_15_FFY_RST,
      O => addr2(14)
    );
  addr2_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_15_FFY_RST
    );
  memtest2_MA_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(15),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_15_FFX_RST,
      O => addr2(15)
    );
  addr2_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_15_FFX_RST
    );
  memtest2_datain_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(13),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_13_FFX_RST,
      O => memtest2_datain(13)
    );
  memtest2_datain_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_13_FFX_RST
    );
  memtest2_datain_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(21),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_21_FFX_RST,
      O => memtest2_datain(21)
    );
  memtest2_datain_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_21_FFX_RST
    );
  memtest2_datain_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(15),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_15_FFX_RST,
      O => memtest2_datain(15)
    );
  memtest2_datain_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_15_FFX_RST
    );
  memtest2_datain_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(23),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_23_FFX_RST,
      O => memtest2_datain(23)
    );
  memtest2_datain_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_23_FFX_RST
    );
  memtest2_datain_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(16),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_17_FFY_RST,
      O => memtest2_datain(16)
    );
  memtest2_datain_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_17_FFY_RST
    );
  memtest_addrcnt_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(2),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_2_FFX_RST,
      O => addr1(2)
    );
  addr1_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_2_FFX_RST
    );
  memtest_addrcnt_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(4),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_4_FFX_RST,
      O => addr1(4)
    );
  addr1_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_4_FFX_RST
    );
  memtest_addrcnt_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(7),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_6_FFY_RST,
      O => addr1(7)
    );
  addr1_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_6_FFY_RST
    );
  memtest_addrcnt_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(11),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_10_FFY_RST,
      O => addr1(11)
    );
  addr1_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_10_FFY_RST
    );
  memtest_addrcnt_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(6),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_6_FFX_RST,
      O => addr1(6)
    );
  addr1_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_6_FFX_RST
    );
  memtest_addrcnt_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcnt_n0000(9),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => addr1_8_FFY_RST,
      O => addr1(9)
    );
  addr1_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr1_8_FFY_RST
    );
  memtest2_deql_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_deq(3),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_deql_2_FFY_RST,
      O => memtest2_deql(3)
    );
  memtest2_deql_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_deql_2_FFY_RST
    );
  memtest2_deql_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_deq_2_rt,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_deql_2_FFX_RST,
      O => memtest2_deql(2)
    );
  memtest2_deql_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_deql_2_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd6_829 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_cs_FFd6_In,
      CE => clkslen,
      CLK => clk,
      SET => maccontrol_PHY_status_MII_Interface_cs_FFd6_FFY_SET,
      RST => GND,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd6
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd6_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd6_FFY_SET
    );
  maccontrol_din_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(0),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_1_FFX_RST,
      O => maccontrol_din(1)
    );
  maccontrol_din_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_1_FFX_RST
    );
  maccontrol_din_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mshreg_sinlll_83,
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_1_FFY_RST,
      O => maccontrol_din(0)
    );
  maccontrol_din_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_1_FFY_RST
    );
  maccontrol_din_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(1),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_3_FFY_RST,
      O => maccontrol_din(2)
    );
  maccontrol_din_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_3_FFY_RST
    );
  maccontrol_lrxmcast_830 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(0),
      CE => maccontrol_n0033,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lrxmcast_FFY_RST,
      O => maccontrol_lrxmcast
    );
  maccontrol_lrxmcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lrxmcast_FFY_RST
    );
  maccontrol_din_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(2),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_3_FFX_RST,
      O => maccontrol_din(3)
    );
  maccontrol_din_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_3_FFX_RST
    );
  maccontrol_din_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(3),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_5_FFY_RST,
      O => maccontrol_din(4)
    );
  maccontrol_din_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_5_FFY_RST
    );
  maccontrol_din_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(5),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_7_FFY_RST,
      O => maccontrol_din(6)
    );
  maccontrol_din_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_7_FFY_RST
    );
  maccontrol_dout_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_23_25_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_23_FFY_RST,
      O => maccontrol_dout(23)
    );
  maccontrol_dout_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_23_FFY_RST
    );
  maccontrol_dout_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_31_25_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_31_FFY_RST,
      O => maccontrol_dout(31)
    );
  maccontrol_dout_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_31_FFY_RST
    );
  maccontrol_dout_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_15_76_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_15_FFY_RST,
      O => maccontrol_dout(15)
    );
  maccontrol_dout_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_15_FFY_RST
    );
  maccontrol_dout_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_24_36_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_24_FFY_RST,
      O => maccontrol_dout(24)
    );
  maccontrol_dout_24_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_24_FFY_RST
    );
  maccontrol_dout_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_16_36_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_16_FFY_RST,
      O => maccontrol_dout(16)
    );
  maccontrol_dout_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_16_FFY_RST
    );
  maccontrol_dout_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_18_22_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_18_FFY_RST,
      O => maccontrol_dout(18)
    );
  maccontrol_dout_18_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_18_FFY_RST
    );
  maccontrol_dout_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_17_36_O,
      CE => maccontrol_n0012,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_17_FFY_RST,
      O => maccontrol_dout(17)
    );
  maccontrol_dout_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_17_FFY_RST
    );
  maccontrol_dout_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mmux_n0023_Result_25_22_O,
      CE => maccontrol_n001223_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_dout_25_FFY_RST,
      O => maccontrol_dout(25)
    );
  maccontrol_dout_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_dout_25_FFY_RST
    );
  memcontroller_Q2_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(29),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_29_FFX_RST,
      O => q2(29)
    );
  q2_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_29_FFX_RST
    );
  memcontroller_Q4_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(10),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_11_FFY_RST,
      O => q4(10)
    );
  q4_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_11_FFY_RST
    );
  memcontroller_Q4_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(11),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_11_FFX_RST,
      O => q4(11)
    );
  q4_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_11_FFX_RST
    );
  memcontroller_Q4_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(20),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_21_FFY_RST,
      O => q4(20)
    );
  q4_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_21_FFY_RST
    );
  memcontroller_Q4_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(21),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_21_FFX_RST,
      O => q4(21)
    );
  q4_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_21_FFX_RST
    );
  memcontroller_Q4_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(12),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_13_FFY_RST,
      O => q4(12)
    );
  q4_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_13_FFY_RST
    );
  memcontroller_Q4_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(13),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_13_FFX_RST,
      O => q4(13)
    );
  q4_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_13_FFX_RST
    );
  memcontroller_Q4_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(30),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_31_FFY_RST,
      O => q4(30)
    );
  q4_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_31_FFY_RST
    );
  memcontroller_Q4_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(31),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_31_FFX_RST,
      O => q4(31)
    );
  q4_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_31_FFX_RST
    );
  memcontroller_Q4_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(22),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_23_FFY_RST,
      O => q4(22)
    );
  q4_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_23_FFY_RST
    );
  memcontroller_Q4_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(23),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_23_FFX_RST,
      O => q4(23)
    );
  q4_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_23_FFX_RST
    );
  memcontroller_Q4_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(14),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_15_FFY_RST,
      O => q4(14)
    );
  q4_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_15_FFY_RST
    );
  memcontroller_Q4_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(15),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_15_FFX_RST,
      O => q4(15)
    );
  q4_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_15_FFX_RST
    );
  memcontroller_Q4_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(24),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_25_FFY_RST,
      O => q4(24)
    );
  q4_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_25_FFY_RST
    );
  memtest2_Mshreg_data4_26_43_831 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_26_net75,
      CE => memtest2_n00511_2,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_26_43_FFY_RST,
      O => memtest2_Mshreg_data4_26_43
    );
  memtest2_Mshreg_data4_26_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_26_43_FFY_RST
    );
  memtest2_Mshreg_data4_19_50_832 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_19_net89,
      CE => memtest2_n00511_3,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_19_50_FFY_RST,
      O => memtest2_Mshreg_data4_19_50
    );
  memtest2_Mshreg_data4_19_50_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_19_50_FFY_RST
    );
  memtest2_Mshreg_data4_27_42_833 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_27_net73,
      CE => memtest2_n00511_2,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_27_42_FFY_RST,
      O => memtest2_Mshreg_data4_27_42
    );
  memtest2_Mshreg_data4_27_42_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_27_42_FFY_RST
    );
  memcontroller_dnl1_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(0),
      CE => memcontroller_dnl1_1_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_1_FFY_RST,
      O => memcontroller_dnl1(0)
    );
  memcontroller_dnl1_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_1_FFY_RST
    );
  memcontroller_dnl1_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(1),
      CE => memcontroller_dnl1_1_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_1_FFX_RST,
      O => memcontroller_dnl1(1)
    );
  memcontroller_dnl1_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_1_FFX_RST
    );
  memcontroller_dnl1_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(2),
      CE => memcontroller_dnl1_3_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_3_FFY_RST,
      O => memcontroller_dnl1(2)
    );
  memcontroller_dnl1_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_3_FFY_RST
    );
  memcontroller_dnl1_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(3),
      CE => memcontroller_dnl1_3_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_3_FFX_RST,
      O => memcontroller_dnl1(3)
    );
  memcontroller_dnl1_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_3_FFX_RST
    );
  memcontroller_dnl1_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(5),
      CE => memcontroller_dnl1_5_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_5_FFX_RST,
      O => memcontroller_dnl1(5)
    );
  memcontroller_dnl1_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_5_FFX_RST
    );
  memcontroller_dnl1_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(7),
      CE => memcontroller_dnl1_7_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_7_FFX_RST,
      O => memcontroller_dnl1(7)
    );
  memcontroller_dnl1_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_7_FFX_RST
    );
  memcontroller_dnl1_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(9),
      CE => memcontroller_dnl1_9_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_9_FFX_RST,
      O => memcontroller_dnl1(9)
    );
  memcontroller_dnl1_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_9_FFX_RST
    );
  memcontroller_clknum_1_2_834 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_n0001(1),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memcontroller_clknum_1_2_FFX_RST,
      O => memcontroller_clknum_1_2
    );
  memcontroller_clknum_1_2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_1_2_FFX_RST
    );
  maccontrol_Mshreg_scslll_84_835 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mshreg_scslll_net281,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => maccontrol_Mshreg_scslll_84_FFY_RST,
      O => maccontrol_Mshreg_scslll_84
    );
  maccontrol_Mshreg_scslll_84_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_Mshreg_scslll_84_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_statecnt_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0014(2),
      CE => maccontrol_PHY_status_MII_Interface_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_statecnt_3_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_statecnt(2)
    );
  maccontrol_PHY_status_MII_Interface_statecnt_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_statecnt_3_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_statecnt_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0014(0),
      CE => maccontrol_PHY_status_MII_Interface_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_statecnt_0_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_statecnt(0)
    );
  maccontrol_PHY_status_MII_Interface_statecnt_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_statecnt_0_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_statecnt_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0014(4),
      CE => maccontrol_PHY_status_MII_Interface_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_statecnt_5_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_statecnt(4)
    );
  maccontrol_PHY_status_MII_Interface_statecnt_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_statecnt_5_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_statecnt_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0014(3),
      CE => maccontrol_PHY_status_MII_Interface_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_statecnt_3_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_statecnt(3)
    );
  maccontrol_PHY_status_MII_Interface_statecnt_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_statecnt_3_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_statecnt_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_n0014(5),
      CE => maccontrol_PHY_status_MII_Interface_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_statecnt_5_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_statecnt(5)
    );
  maccontrol_PHY_status_MII_Interface_statecnt_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_statecnt_5_FFX_RST
    );
  memcontroller_dnl1_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(10),
      CE => memcontroller_dnl1_11_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_11_FFY_RST,
      O => memcontroller_dnl1(10)
    );
  memcontroller_dnl1_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_11_FFY_RST
    );
  memcontroller_dnl1_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(11),
      CE => memcontroller_dnl1_11_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_11_FFX_RST,
      O => memcontroller_dnl1(11)
    );
  memcontroller_dnl1_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_11_FFX_RST
    );
  memcontroller_dnl1_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(21),
      CE => memcontroller_dnl1_21_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_21_FFX_RST,
      O => memcontroller_dnl1(21)
    );
  memcontroller_dnl1_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_21_FFX_RST
    );
  memcontroller_dnl1_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(13),
      CE => memcontroller_dnl1_13_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_13_FFX_RST,
      O => memcontroller_dnl1(13)
    );
  memcontroller_dnl1_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_13_FFX_RST
    );
  memcontroller_dnl1_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(31),
      CE => memcontroller_dnl1_31_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_31_FFX_RST,
      O => memcontroller_dnl1(31)
    );
  memcontroller_dnl1_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_31_FFX_RST
    );
  memtest_Mshreg_dataw4_4_33_836 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_4_net55,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_4_33_FFY_RST,
      O => memtest_Mshreg_dataw4_4_33
    );
  memtest_Mshreg_dataw4_4_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_4_33_FFY_RST
    );
  maccontrol_PHY_status_PHYADDRSTATUS : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyaddr_31_FROM,
      CE => maccontrol_PHY_status_n00171_O,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_31_FFX_RST,
      O => maccontrol_phyaddr(31)
    );
  maccontrol_phyaddr_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_31_FFX_RST
    );
  memtest_Mshreg_dataw4_5_32_837 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_5_net53,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_5_32_FFY_RST,
      O => memtest_Mshreg_dataw4_5_32
    );
  memtest_Mshreg_dataw4_5_32_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_5_32_FFY_RST
    );
  memtest2_Mshreg_data4_11_58_838 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_11_net105,
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_11_58_FFY_RST,
      O => memtest2_Mshreg_data4_11_58
    );
  memtest2_Mshreg_data4_11_58_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_11_58_FFY_RST
    );
  memtest_Mshreg_dataw4_6_31_839 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_6_net51,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_6_31_FFY_RST,
      O => memtest_Mshreg_dataw4_6_31
    );
  memtest_Mshreg_dataw4_6_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_6_31_FFY_RST
    );
  memtest2_Mshreg_data4_12_57_840 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_12_net103,
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_12_57_FFY_RST,
      O => memtest2_Mshreg_data4_12_57
    );
  memtest2_Mshreg_data4_12_57_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_12_57_FFY_RST
    );
  memtest_Mshreg_dataw4_7_30_841 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_7_net49,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_7_30_FFY_RST,
      O => memtest_Mshreg_dataw4_7_30
    );
  memtest_Mshreg_dataw4_7_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_7_30_FFY_RST
    );
  memtest_Mshreg_dataw4_8_29_842 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_8_net47,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_8_29_FFY_RST,
      O => memtest_Mshreg_dataw4_8_29
    );
  memtest_Mshreg_dataw4_8_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_8_29_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd3_843 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_cs_FFd3_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_cs_FFd3_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd3
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd3_FFY_RST
    );
  memtest2_Mshreg_data4_14_55_844 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_14_net99,
      CE => memtest2_n00511_3,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_14_55_FFY_RST,
      O => memtest2_Mshreg_data4_14_55
    );
  memtest2_Mshreg_data4_14_55_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_14_55_FFY_RST
    );
  memtest2_Mshreg_data4_22_47_845 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_22_net83,
      CE => memtest2_n00511_2,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_22_47_FFY_RST,
      O => memtest2_Mshreg_data4_22_47
    );
  memtest2_Mshreg_data4_22_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_22_47_FFY_RST
    );
  maccontrol_phyaddr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(3),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_3_FFY_RST,
      O => maccontrol_phyaddr(3)
    );
  maccontrol_phyaddr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_3_FFY_RST
    );
  maccontrol_phyaddr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(1),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_1_FFX_RST,
      O => maccontrol_phyaddr(1)
    );
  maccontrol_phyaddr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_1_FFX_RST
    );
  maccontrol_phyaddr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(5),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_5_FFX_RST,
      O => maccontrol_phyaddr(5)
    );
  maccontrol_phyaddr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_5_FFX_RST
    );
  maccontrol_phyaddr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(7),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_7_FFX_RST,
      O => maccontrol_phyaddr(7)
    );
  maccontrol_phyaddr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_7_FFX_RST
    );
  maccontrol_phyaddr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(9),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_9_FFX_RST,
      O => maccontrol_phyaddr(9)
    );
  maccontrol_phyaddr_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_9_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(1),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_1_FFX_RST,
      O => maccontrol_PHY_status_dout(1)
    );
  maccontrol_PHY_status_dout_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_1_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(3),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_3_FFX_RST,
      O => maccontrol_PHY_status_dout(3)
    );
  maccontrol_PHY_status_dout_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_3_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(6),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_7_FFY_RST,
      O => maccontrol_PHY_status_dout(6)
    );
  maccontrol_PHY_status_dout_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_7_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(5),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_5_FFX_RST,
      O => maccontrol_PHY_status_dout(5)
    );
  maccontrol_PHY_status_dout_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_5_FFX_RST
    );
  memcontroller_dnl1_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(23),
      CE => memcontroller_dnl1_23_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_23_FFX_RST,
      O => memcontroller_dnl1(23)
    );
  memcontroller_dnl1_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_23_FFX_RST
    );
  memcontroller_dnl1_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(15),
      CE => memcontroller_dnl1_15_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_15_FFX_RST,
      O => memcontroller_dnl1(15)
    );
  memcontroller_dnl1_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_15_FFX_RST
    );
  memcontroller_dnl1_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(25),
      CE => memcontroller_dnl1_25_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_25_FFX_RST,
      O => memcontroller_dnl1(25)
    );
  memcontroller_dnl1_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_25_FFX_RST
    );
  memcontroller_dnl1_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(17),
      CE => memcontroller_dnl1_17_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_17_FFX_RST,
      O => memcontroller_dnl1(17)
    );
  memcontroller_dnl1_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_17_FFX_RST
    );
  memcontroller_dnl1_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(27),
      CE => memcontroller_dnl1_27_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl1_27_FFX_RST,
      O => memcontroller_dnl1(27)
    );
  memcontroller_dnl1_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_27_FFX_RST
    );
  memtest_Mshreg_dataw4_20_17_846 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_20_net23,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_20_17_FFY_RST,
      O => memtest_Mshreg_dataw4_20_17
    );
  memtest_Mshreg_dataw4_20_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_20_17_FFY_RST
    );
  memtest2_Mshreg_data4_4_65_847 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_4_net119,
      CE => memtest2_n00511_1,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_4_65_FFY_RST,
      O => memtest2_Mshreg_data4_4_65
    );
  memtest2_Mshreg_data4_4_65_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_4_65_FFY_RST
    );
  memtest_Mshreg_dataw4_13_24_848 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_13_net37,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_13_24_FFY_RST,
      O => memtest_Mshreg_dataw4_13_24
    );
  memtest_Mshreg_dataw4_13_24_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_13_24_FFY_RST
    );
  memtest_Mshreg_dataw4_21_16_849 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_21_net21,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_21_16_FFY_RST,
      O => memtest_Mshreg_dataw4_21_16
    );
  memtest_Mshreg_dataw4_21_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_21_16_FFY_RST
    );
  memtest2_Mshreg_data4_5_64_850 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_5_net117,
      CE => memtest2_n00511_1,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_5_64_FFY_RST,
      O => memtest2_Mshreg_data4_5_64
    );
  memtest2_Mshreg_data4_5_64_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_5_64_FFY_RST
    );
  testrx_cs_FFd2_851 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_cs_FFd2_In,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => testrx_cs_FFd2_FFY_RST,
      O => testrx_cs_FFd2
    );
  testrx_cs_FFd2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => testrx_cs_FFd2_FFY_RST
    );
  memtest_Mshreg_dataw4_14_23_852 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_14_net35,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_14_23_FFY_RST,
      O => memtest_Mshreg_dataw4_14_23
    );
  memtest_Mshreg_dataw4_14_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_14_23_FFY_RST
    );
  memtest_Mshreg_dataw4_22_15_853 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_22_net19,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_22_15_FFY_RST,
      O => memtest_Mshreg_dataw4_22_15
    );
  memtest_Mshreg_dataw4_22_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_22_15_FFY_RST
    );
  testrx_cs_FFd3_854 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => testrx_cs_FFd3_In,
      CE => VCC,
      CLK => rx_clk_int,
      SET => testrx_cs_FFd3_FFY_SET,
      RST => GND,
      O => testrx_cs_FFd3
    );
  testrx_cs_FFd3_FFY_SETOR : X_BUF
    port map (
      I => GSR,
      O => testrx_cs_FFd3_FFY_SET
    );
  memtest2_Mshreg_data4_6_63_855 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_6_net115,
      CE => memtest2_n00511_1,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_6_63_FFY_RST,
      O => memtest2_Mshreg_data4_6_63
    );
  memtest2_Mshreg_data4_6_63_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_6_63_FFY_RST
    );
  maccontrol_PHY_status_PHYDOUT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(2),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_3_FFY_RST,
      O => maccontrol_phydo(2)
    );
  maccontrol_phydo_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_3_FFY_RST
    );
  maccontrol_PHY_status_PHYDOUT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(1),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_1_FFX_RST,
      O => maccontrol_phydo(1)
    );
  maccontrol_phydo_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_1_FFX_RST
    );
  maccontrol_PHY_status_PHYDOUT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(3),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_3_FFX_RST,
      O => maccontrol_phydo(3)
    );
  maccontrol_phydo_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_3_FFX_RST
    );
  maccontrol_PHY_status_PHYDOUT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(6),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_7_FFY_RST,
      O => maccontrol_phydo(6)
    );
  maccontrol_phydo_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_7_FFY_RST
    );
  maccontrol_PHY_status_PHYDOUT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(5),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_5_FFX_RST,
      O => maccontrol_phydo(5)
    );
  maccontrol_phydo_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_5_FFX_RST
    );
  maccontrol_PHY_status_PHYDOUT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(7),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_7_FFX_RST,
      O => maccontrol_phydo(7)
    );
  maccontrol_phydo_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_7_FFX_RST
    );
  memtest_addrcntll_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(1),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_1_FFX_RST,
      O => addr4(1)
    );
  addr4_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_1_FFX_RST
    );
  maccontrol_PHY_status_PHYDOUT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(9),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_9_FFX_RST,
      O => maccontrol_phydo(9)
    );
  maccontrol_phydo_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_9_FFX_RST
    );
  memtest_addrcntll_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(4),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_5_FFY_RST,
      O => addr4(4)
    );
  addr4_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_5_FFY_RST
    );
  maccontrol_din_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(10),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_11_FFX_RST,
      O => maccontrol_din(11)
    );
  maccontrol_din_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_11_FFX_RST
    );
  maccontrol_phydi_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(5),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_5_FFX_RST,
      O => maccontrol_phydi(5)
    );
  maccontrol_phydi_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_5_FFX_RST
    );
  maccontrol_din_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(12),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_13_FFX_RST,
      O => maccontrol_din(13)
    );
  maccontrol_din_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_13_FFX_RST
    );
  maccontrol_din_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(19),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_21_FFY_RST,
      O => maccontrol_din(20)
    );
  maccontrol_din_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_21_FFY_RST
    );
  maccontrol_din_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(20),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_21_FFX_RST,
      O => maccontrol_din(21)
    );
  maccontrol_din_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_21_FFX_RST
    );
  maccontrol_phydi_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(6),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_7_FFY_RST,
      O => maccontrol_phydi(6)
    );
  maccontrol_phydi_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_7_FFY_RST
    );
  maccontrol_phydi_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(7),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_7_FFX_RST,
      O => maccontrol_phydi(7)
    );
  maccontrol_phydi_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_7_FFX_RST
    );
  maccontrol_din_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(13),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_15_FFY_RST,
      O => maccontrol_din(14)
    );
  maccontrol_din_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_15_FFY_RST
    );
  maccontrol_din_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(14),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_15_FFX_RST,
      O => maccontrol_din(15)
    );
  maccontrol_din_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_15_FFX_RST
    );
  maccontrol_din_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(21),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_23_FFY_RST,
      O => maccontrol_din(22)
    );
  maccontrol_din_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_23_FFY_RST
    );
  maccontrol_din_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(22),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_23_FFX_RST,
      O => maccontrol_din(23)
    );
  maccontrol_din_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_23_FFX_RST
    );
  maccontrol_din_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(29),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_31_FFY_RST,
      O => maccontrol_din(30)
    );
  maccontrol_din_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_31_FFY_RST
    );
  maccontrol_din_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(30),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_31_FFX_RST,
      O => maccontrol_din(31)
    );
  maccontrol_din_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_31_FFX_RST
    );
  maccontrol_phydi_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(8),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_9_FFY_RST,
      O => maccontrol_phydi(8)
    );
  maccontrol_phydi_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_9_FFY_RST
    );
  maccontrol_din_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(15),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_17_FFY_RST,
      O => maccontrol_din(16)
    );
  maccontrol_din_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_17_FFY_RST
    );
  maccontrol_phydi_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(9),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_9_FFX_RST,
      O => maccontrol_phydi(9)
    );
  maccontrol_phydi_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_9_FFX_RST
    );
  memtest2_datain_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(17),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_17_FFX_RST,
      O => memtest2_datain(17)
    );
  memtest2_datain_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_17_FFX_RST
    );
  memtest2_datain_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(25),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_25_FFX_RST,
      O => memtest2_datain(25)
    );
  memtest2_datain_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_25_FFX_RST
    );
  memtest2_MD_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(11),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_11_FFX_RST,
      O => d2(11)
    );
  d2_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_11_FFX_RST
    );
  memtest2_datain_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(18),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_19_FFY_RST,
      O => memtest2_datain(18)
    );
  memtest2_datain_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_19_FFY_RST
    );
  memtest2_MD_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(12),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_13_FFY_RST,
      O => d2(12)
    );
  d2_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_13_FFY_RST
    );
  memtest2_datain_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(19),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_19_FFX_RST,
      O => memtest2_datain(19)
    );
  memtest2_datain_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_19_FFX_RST
    );
  memtest2_datain_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(27),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_27_FFY_RST,
      O => memtest2_datain(27)
    );
  memtest2_datain_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_27_FFY_RST
    );
  memtest2_MD_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(21),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_21_FFY_RST,
      O => d2(21)
    );
  d2_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_21_FFY_RST
    );
  memtest2_MD_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(13),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_13_FFX_RST,
      O => d2(13)
    );
  d2_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_13_FFX_RST
    );
  memtest2_datain_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(28),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_29_FFY_RST,
      O => memtest2_datain(28)
    );
  memtest2_datain_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_29_FFY_RST
    );
  memtest2_datain_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(29),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_29_FFX_RST,
      O => memtest2_datain(29)
    );
  memtest2_datain_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_29_FFX_RST
    );
  memtest2_MD_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(30),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_31_FFY_RST,
      O => d2(30)
    );
  d2_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_31_FFY_RST
    );
  memtest_Mshreg_dataw4_15_22_856 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_15_net33,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_15_22_FFY_RST,
      O => memtest_Mshreg_dataw4_15_22
    );
  memtest_Mshreg_dataw4_15_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_15_22_FFY_RST
    );
  memtest_Mshreg_dataw4_23_14_857 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_23_net17,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_23_14_FFY_RST,
      O => memtest_Mshreg_dataw4_23_14
    );
  memtest_Mshreg_dataw4_23_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_23_14_FFY_RST
    );
  memtest2_Mshreg_data4_7_62_858 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_7_net113,
      CE => memtest2_n00511_1,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_7_62_FFY_RST,
      O => memtest2_Mshreg_data4_7_62
    );
  memtest2_Mshreg_data4_7_62_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_7_62_FFY_RST
    );
  memtest_Mshreg_dataw4_16_21_859 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_16_net31,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_16_21_FFY_RST,
      O => memtest_Mshreg_dataw4_16_21
    );
  memtest_Mshreg_dataw4_16_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_16_21_FFY_RST
    );
  memtest_Mshreg_dataw4_24_13_860 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_24_net15,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_24_13_FFY_RST,
      O => memtest_Mshreg_dataw4_24_13
    );
  memtest_Mshreg_dataw4_24_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_24_13_FFY_RST
    );
  memtest2_Mshreg_data4_8_61_861 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_8_net111,
      CE => memtest2_n00511_1,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_8_61_FFY_RST,
      O => memtest2_Mshreg_data4_8_61
    );
  memtest2_Mshreg_data4_8_61_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_8_61_FFY_RST
    );
  memtest_Mshreg_dataw4_17_20_862 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_17_net29,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_17_20_FFY_RST,
      O => memtest_Mshreg_dataw4_17_20
    );
  memtest_Mshreg_dataw4_17_20_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_17_20_FFY_RST
    );
  memtest_Mshreg_dataw4_25_12_863 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_25_net13,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_25_12_FFY_RST,
      O => memtest_Mshreg_dataw4_25_12
    );
  memtest_Mshreg_dataw4_25_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_25_12_FFY_RST
    );
  memtest_Mshreg_dataw4_18_19_864 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_18_net27,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_18_19_FFY_RST,
      O => memtest_Mshreg_dataw4_18_19
    );
  memtest_Mshreg_dataw4_18_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_18_19_FFY_RST
    );
  memtest2_Mshreg_data4_9_60_865 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_Mshreg_data4_9_net109,
      CE => memtest2_n00511_1,
      CLK => clk,
      SET => GND,
      RST => memtest2_Mshreg_data4_9_60_FFY_RST,
      O => memtest2_Mshreg_data4_9_60
    );
  memtest2_Mshreg_data4_9_60_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_Mshreg_data4_9_60_FFY_RST
    );
  memtest_Mshreg_dataw4_26_11_866 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_Mshreg_dataw4_26_net11,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_Mshreg_dataw4_26_11_FFY_RST,
      O => memtest_Mshreg_dataw4_26_11
    );
  memtest_Mshreg_dataw4_26_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_Mshreg_dataw4_26_11_FFY_RST
    );
  memcontroller_Q4_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(1),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_1_FFX_RST,
      O => q4(1)
    );
  q4_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_1_FFX_RST
    );
  memcontroller_Q4_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(2),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_3_FFY_RST,
      O => q4(2)
    );
  q4_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_3_FFY_RST
    );
  memcontroller_Q4_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(3),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_3_FFX_RST,
      O => q4(3)
    );
  q4_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_3_FFX_RST
    );
  memcontroller_Q4_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(4),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_5_FFY_RST,
      O => q4(4)
    );
  q4_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_5_FFY_RST
    );
  memcontroller_Q4_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(5),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_5_FFX_RST,
      O => q4(5)
    );
  q4_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_5_FFX_RST
    );
  memcontroller_Q4_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(6),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_7_FFY_RST,
      O => q4(6)
    );
  q4_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_7_FFY_RST
    );
  memcontroller_Q4_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(7),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_7_FFX_RST,
      O => q4(7)
    );
  q4_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_7_FFX_RST
    );
  memcontroller_Q4_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(8),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_9_FFY_RST,
      O => q4(8)
    );
  q4_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_9_FFY_RST
    );
  memcontroller_Q4_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(9),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_9_FFX_RST,
      O => q4(9)
    );
  q4_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_9_FFX_RST
    );
  maccontrol_phyaddr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(0),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_1_FFY_RST,
      O => maccontrol_phyaddr(0)
    );
  maccontrol_phyaddr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_1_FFY_RST
    );
  memtest2_MD_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(31),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_31_FFX_RST,
      O => d2(31)
    );
  d2_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_31_FFX_RST
    );
  memtest2_MD_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(22),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_22_FFY_RST,
      O => d2(22)
    );
  d2_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_22_FFY_RST
    );
  memtest2_MD_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(14),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_15_FFY_RST,
      O => d2(14)
    );
  d2_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_15_FFY_RST
    );
  memtest2_MD_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(15),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_15_FFX_RST,
      O => d2(15)
    );
  d2_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_15_FFX_RST
    );
  memtest2_MD_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(24),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_25_FFY_RST,
      O => d2(24)
    );
  d2_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_25_FFY_RST
    );
  memtest2_MD_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(25),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_25_FFX_RST,
      O => d2(25)
    );
  d2_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_25_FFX_RST
    );
  memtest2_MD_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(16),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_17_FFY_RST,
      O => d2(16)
    );
  d2_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_17_FFY_RST
    );
  memtest2_MD_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(17),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_17_FFX_RST,
      O => d2(17)
    );
  d2_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_17_FFX_RST
    );
  memtest2_MD_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(26),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_27_FFY_RST,
      O => d2(26)
    );
  d2_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_27_FFY_RST
    );
  memtest2_MD_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(27),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_27_FFX_RST,
      O => d2(27)
    );
  d2_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_27_FFX_RST
    );
  memtest2_MD_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(18),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_19_FFY_RST,
      O => d2(18)
    );
  d2_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_19_FFY_RST
    );
  memtest2_MD_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(19),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_19_FFX_RST,
      O => d2(19)
    );
  d2_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_19_FFX_RST
    );
  memtest2_MD_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(28),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_29_FFY_RST,
      O => d2(28)
    );
  d2_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_29_FFY_RST
    );
  memtest2_MD_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(29),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_29_FFX_RST,
      O => d2(29)
    );
  d2_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_29_FFX_RST
    );
  maccontrol_PHY_status_PHYDOUT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(0),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_1_FFY_RST,
      O => maccontrol_phydo(0)
    );
  maccontrol_phydo_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_1_FFY_RST
    );
  memcontroller_Q4_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(25),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_25_FFX_RST,
      O => q4(25)
    );
  q4_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_25_FFX_RST
    );
  memcontroller_Q4_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(16),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_17_FFY_RST,
      O => q4(16)
    );
  q4_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_17_FFY_RST
    );
  memcontroller_Q4_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(17),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_17_FFX_RST,
      O => q4(17)
    );
  q4_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_17_FFX_RST
    );
  memcontroller_Q4_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(26),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_27_FFY_RST,
      O => q4(26)
    );
  q4_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_27_FFY_RST
    );
  memcontroller_Q4_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(27),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_27_FFX_RST,
      O => q4(27)
    );
  q4_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_27_FFX_RST
    );
  memcontroller_Q4_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(18),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_19_FFY_RST,
      O => q4(18)
    );
  q4_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_19_FFY_RST
    );
  memcontroller_Q4_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(19),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_19_FFX_RST,
      O => q4(19)
    );
  q4_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_19_FFX_RST
    );
  memcontroller_Q4_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(28),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_29_FFY_RST,
      O => q4(28)
    );
  q4_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_29_FFY_RST
    );
  memcontroller_Q4_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(29),
      CE => memcontroller_n0007,
      CLK => clk,
      SET => GND,
      RST => q4_29_FFX_RST,
      O => q4(29)
    );
  q4_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q4_29_FFX_RST
    );
  memtest2_ldata_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(7),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_7_FFX_RST,
      O => memtest2_ldata(7)
    );
  memtest2_ldata_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_7_FFX_RST
    );
  memcontroller_Q2_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(3),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_3_FFX_RST,
      O => q2(3)
    );
  q2_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_3_FFX_RST
    );
  memtest2_ldata_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(9),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_9_FFX_RST,
      O => memtest2_ldata(9)
    );
  memtest2_ldata_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_9_FFX_RST
    );
  memcontroller_Q2_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(5),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_5_FFX_RST,
      O => q2(5)
    );
  q2_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_5_FFX_RST
    );
  memcontroller_Q2_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(6),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_7_FFY_RST,
      O => q2(6)
    );
  q2_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_7_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_cs_FFd2,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_done_FFY_RST,
      O => maccontrol_PHY_status_done
    );
  maccontrol_PHY_status_done_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_done_FFY_RST
    );
  memcontroller_Q2_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(7),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_7_FFX_RST,
      O => q2(7)
    );
  q2_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_7_FFX_RST
    );
  memcontroller_Q2_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(8),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_9_FFY_RST,
      O => q2(8)
    );
  q2_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_9_FFY_RST
    );
  memcontroller_Q2_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(9),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_9_FFX_RST,
      O => q2(9)
    );
  q2_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_9_FFX_RST
    );
  memtest_addrcntll_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(3),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_3_FFX_RST,
      O => addr4(3)
    );
  addr4_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_3_FFX_RST
    );
  memtest_addrcntll_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(5),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_5_FFX_RST,
      O => addr4(5)
    );
  addr4_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_5_FFX_RST
    );
  memtest_addrcntll_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(7),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_7_FFX_RST,
      O => addr4(7)
    );
  addr4_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_7_FFX_RST
    );
  memtest_addrcntll_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(9),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_9_FFX_RST,
      O => addr4(9)
    );
  addr4_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_9_FFX_RST
    );
  memtest2_ldata_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(1),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_1_FFX_RST,
      O => memtest2_ldata(1)
    );
  memtest2_ldata_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_1_FFX_RST
    );
  memtest2_ldata_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(2),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_3_FFY_RST,
      O => memtest2_ldata(2)
    );
  memtest2_ldata_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_3_FFY_RST
    );
  memtest2_ldata_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(3),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_3_FFX_RST,
      O => memtest2_ldata(3)
    );
  memtest2_ldata_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_3_FFX_RST
    );
  memtest2_ldata_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(5),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_5_FFX_RST,
      O => memtest2_ldata(5)
    );
  memtest2_ldata_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_5_FFX_RST
    );
  memcontroller_Q2_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(0),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_1_FFY_RST,
      O => q2(0)
    );
  q2_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_1_FFY_RST
    );
  memcontroller_Q2_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(1),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_1_FFX_RST,
      O => q2(1)
    );
  q2_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_1_FFX_RST
    );
  maccontrol_phyaddr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(13),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_13_FFX_RST,
      O => maccontrol_phyaddr(13)
    );
  maccontrol_phyaddr_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_13_FFX_RST
    );
  maccontrol_phyaddr_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(20),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_21_FFY_RST,
      O => maccontrol_phyaddr(20)
    );
  maccontrol_phyaddr_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_21_FFY_RST
    );
  maccontrol_phyaddr_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(21),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_21_FFX_RST,
      O => maccontrol_phyaddr(21)
    );
  maccontrol_phyaddr_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_21_FFX_RST
    );
  maccontrol_phyaddr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(14),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_15_FFY_RST,
      O => maccontrol_phyaddr(14)
    );
  maccontrol_phyaddr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_15_FFY_RST
    );
  maccontrol_phyaddr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(15),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_15_FFX_RST,
      O => maccontrol_phyaddr(15)
    );
  maccontrol_phyaddr_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_15_FFX_RST
    );
  maccontrol_phyaddr_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(30),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_30_FFY_RST,
      O => maccontrol_phyaddr(30)
    );
  maccontrol_phyaddr_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_30_FFY_RST
    );
  maccontrol_phyaddr_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(22),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_22_FFY_RST,
      O => maccontrol_phyaddr(22)
    );
  maccontrol_phyaddr_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_22_FFY_RST
    );
  maccontrol_phyaddr_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(23),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_23_FFY_RST,
      O => maccontrol_phyaddr(23)
    );
  maccontrol_phyaddr_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_23_FFY_RST
    );
  maccontrol_phyaddr_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(16),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_17_FFY_RST,
      O => maccontrol_phyaddr(16)
    );
  maccontrol_phyaddr_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_17_FFY_RST
    );
  maccontrol_phyaddr_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(17),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_17_FFX_RST,
      O => maccontrol_phyaddr(17)
    );
  maccontrol_phyaddr_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_17_FFX_RST
    );
  maccontrol_phyaddr_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(25),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_25_FFX_RST,
      O => maccontrol_phyaddr(25)
    );
  maccontrol_phyaddr_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_25_FFX_RST
    );
  maccontrol_phyaddr_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(26),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_27_FFY_RST,
      O => maccontrol_phyaddr(26)
    );
  maccontrol_phyaddr_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_27_FFY_RST
    );
  maccontrol_phyaddr_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(19),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_19_FFX_RST,
      O => maccontrol_phyaddr(19)
    );
  maccontrol_phyaddr_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_19_FFX_RST
    );
  testrx_rxdll_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_rxdl(7),
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => testrx_rxdll_7_FFX_RST,
      O => testrx_rxdll(7)
    );
  testrx_rxdll_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => testrx_rxdll_7_FFX_RST
    );
  memcontroller_dnl2_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(10),
      CE => memcontroller_dnl2_11_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_11_FFY_RST,
      O => memcontroller_dnl2(10)
    );
  memcontroller_dnl2_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_11_FFY_RST
    );
  memcontroller_dnl2_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(11),
      CE => memcontroller_dnl2_11_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_11_FFX_RST,
      O => memcontroller_dnl2(11)
    );
  memcontroller_dnl2_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_11_FFX_RST
    );
  memtest_dataw1_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(10),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_11_FFY_RST,
      O => memtest_dataw1(10)
    );
  memtest_dataw1_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_11_FFY_RST
    );
  memtest_dataw1_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(11),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_11_FFX_RST,
      O => memtest_dataw1(11)
    );
  memtest_dataw1_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_11_FFX_RST
    );
  memcontroller_dnl2_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(20),
      CE => memcontroller_dnl2_21_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_21_FFY_RST,
      O => memcontroller_dnl2(20)
    );
  memcontroller_dnl2_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_21_FFY_RST
    );
  memcontroller_dnl2_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(21),
      CE => memcontroller_dnl2_21_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_21_FFX_RST,
      O => memcontroller_dnl2(21)
    );
  memcontroller_dnl2_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_21_FFX_RST
    );
  memcontroller_dnl2_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(12),
      CE => memcontroller_dnl2_13_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_13_FFY_RST,
      O => memcontroller_dnl2(12)
    );
  memcontroller_dnl2_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_13_FFY_RST
    );
  memcontroller_dnl2_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(13),
      CE => memcontroller_dnl2_13_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_13_FFX_RST,
      O => memcontroller_dnl2(13)
    );
  memcontroller_dnl2_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_13_FFX_RST
    );
  memtest_dataw1_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(20),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_21_FFY_RST,
      O => memtest_dataw1(20)
    );
  memtest_dataw1_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_21_FFY_RST
    );
  memtest_dataw1_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(21),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_21_FFX_RST,
      O => memtest_dataw1(21)
    );
  memtest_dataw1_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_21_FFX_RST
    );
  memtest_dataw1_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(12),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_13_FFY_RST,
      O => memtest_dataw1(12)
    );
  memtest_dataw1_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_13_FFY_RST
    );
  memtest_dataw1_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(13),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_13_FFX_RST,
      O => memtest_dataw1(13)
    );
  memtest_dataw1_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_13_FFX_RST
    );
  memcontroller_dnl2_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(30),
      CE => memcontroller_dnl2_31_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_31_FFY_RST,
      O => memcontroller_dnl2(30)
    );
  memcontroller_dnl2_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_31_FFY_RST
    );
  maccontrol_phyaddr_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(27),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_27_FFX_RST,
      O => maccontrol_phyaddr(27)
    );
  maccontrol_phyaddr_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_27_FFX_RST
    );
  maccontrol_phyaddr_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(29),
      CE => maccontrol_n00311_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_29_FFX_RST,
      O => maccontrol_phyaddr(29)
    );
  maccontrol_phyaddr_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_29_FFX_RST
    );
  txsim_llltx_867 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_n0002,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => txsim_llltx_FFY_RST,
      O => txsim_llltx
    );
  txsim_llltx_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txsim_llltx_FFY_RST
    );
  memtest_llerr_868 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_llerr_BXMUXNOT,
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => memtest_llerr_FFX_RST,
      O => memtest_llerr
    );
  memtest_llerr_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_llerr_FFX_RST
    );
  testrx_rxdll_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_rxdl(0),
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => testrx_rxdll_1_FFY_RST,
      O => testrx_rxdll(0)
    );
  testrx_rxdll_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => testrx_rxdll_1_FFY_RST
    );
  testrx_rxdll_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_rxdl(1),
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => testrx_rxdll_1_FFX_RST,
      O => testrx_rxdll(1)
    );
  testrx_rxdll_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => testrx_rxdll_1_FFX_RST
    );
  testrx_rxdll_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_rxdl(2),
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => testrx_rxdll_3_FFY_RST,
      O => testrx_rxdll(2)
    );
  testrx_rxdll_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => testrx_rxdll_3_FFY_RST
    );
  testrx_rxdll_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_rxdl(4),
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => testrx_rxdll_5_FFY_RST,
      O => testrx_rxdll(4)
    );
  testrx_rxdll_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => testrx_rxdll_5_FFY_RST
    );
  testrx_rxdll_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_rxdl(3),
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => testrx_rxdll_3_FFX_RST,
      O => testrx_rxdll(3)
    );
  testrx_rxdll_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => testrx_rxdll_3_FFX_RST
    );
  memtest2_cs_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => memtest2_cs_0_BYMUXNOT,
      CE => memtest2_n0117,
      CLK => clk,
      SET => memtest2_cs_0_FFY_SET,
      RST => GND,
      O => memtest2_cs(0)
    );
  memtest2_cs_0_FFY_SETOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_cs_0_FFY_SET
    );
  testrx_rxdll_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_rxdl(6),
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => testrx_rxdll_7_FFY_RST,
      O => testrx_rxdll(6)
    );
  testrx_rxdll_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => testrx_rxdll_7_FFY_RST
    );
  testrx_rxdll_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_rxdl(5),
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => testrx_rxdll_5_FFX_RST,
      O => testrx_rxdll(5)
    );
  testrx_rxdll_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => testrx_rxdll_5_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(7),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_7_FFX_RST,
      O => maccontrol_PHY_status_dout(7)
    );
  maccontrol_PHY_status_dout_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_7_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(9),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_9_FFX_RST,
      O => maccontrol_PHY_status_dout(9)
    );
  maccontrol_PHY_status_dout_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_9_FFX_RST
    );
  maccontrol_PHY_status_PHYDOUT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(11),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_11_FFX_RST,
      O => maccontrol_phydo(11)
    );
  maccontrol_phydo_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_11_FFX_RST
    );
  maccontrol_PHY_status_PHYDOUT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(13),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_13_FFX_RST,
      O => maccontrol_phydo(13)
    );
  maccontrol_phydo_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_13_FFX_RST
    );
  maccontrol_PHY_status_PHYDOUT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(15),
      CE => maccontrol_PHY_status_n0021,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydo_15_FFX_RST,
      O => maccontrol_phydo(15)
    );
  maccontrol_phydo_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydo_15_FFX_RST
    );
  memtest_addrcntll_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(11),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_11_FFX_RST,
      O => addr4(11)
    );
  addr4_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_11_FFX_RST
    );
  memtest_addrcntll_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(13),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_13_FFX_RST,
      O => addr4(13)
    );
  addr4_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_13_FFX_RST
    );
  memtest2_datalfsr_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(9),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(10)
    );
  memtest_addrcntll_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_addrcntl(15),
      CE => clken4,
      CLK => clk,
      SET => GND,
      RST => addr4_15_FFX_RST,
      O => addr4(15)
    );
  addr4_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr4_15_FFX_RST
    );
  maccontrol_lmacaddr_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(7),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_23_FFX_RST,
      O => maccontrol_lmacaddr(23)
    );
  maccontrol_lmacaddr_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_23_FFX_RST
    );
  maccontrol_lmacaddr_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(15),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_31_FFX_RST,
      O => maccontrol_lmacaddr(31)
    );
  maccontrol_lmacaddr_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_31_FFX_RST
    );
  maccontrol_lmacaddr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(15),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_15_FFX_RST,
      O => maccontrol_lmacaddr(15)
    );
  maccontrol_lmacaddr_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_15_FFX_RST
    );
  memtest2_ldata_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(11),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_11_FFX_RST,
      O => memtest2_ldata(11)
    );
  memtest2_ldata_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_11_FFX_RST
    );
  memcontroller_dnl2_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(6),
      CE => memcontroller_dnl2_7_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_7_FFY_RST,
      O => memcontroller_dnl2(6)
    );
  memcontroller_dnl2_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_7_FFY_RST
    );
  memcontroller_dnl2_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(7),
      CE => memcontroller_dnl2_7_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_7_FFX_RST,
      O => memcontroller_dnl2(7)
    );
  memcontroller_dnl2_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_7_FFX_RST
    );
  maccontrol_lmacaddr_32 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(0),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_33_FFY_RST,
      O => maccontrol_lmacaddr(32)
    );
  maccontrol_lmacaddr_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_33_FFY_RST
    );
  maccontrol_lmacaddr_33 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(1),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_33_FFX_RST,
      O => maccontrol_lmacaddr(33)
    );
  maccontrol_lmacaddr_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_33_FFX_RST
    );
  maccontrol_lmacaddr_41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(9),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_41_FFX_RST,
      O => maccontrol_lmacaddr(41)
    );
  maccontrol_lmacaddr_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_41_FFX_RST
    );
  maccontrol_lmacaddr_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(1),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_17_FFX_RST,
      O => maccontrol_lmacaddr(17)
    );
  maccontrol_lmacaddr_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_17_FFX_RST
    );
  memcontroller_clknum_0_1_869 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_0_2_BYMUXNOT,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memcontroller_clknum_0_2_FFY_RST,
      O => memcontroller_clknum_0_1
    );
  memcontroller_clknum_0_2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_0_2_FFY_RST
    );
  memtest2_datalfsr_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(10),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(11)
    );
  memtest2_datalfsr_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(19),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(20)
    );
  memtest2_datalfsr_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(20),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(21)
    );
  memtest2_datalfsr_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(12),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(13)
    );
  memtest2_datalfsr_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(14),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(15)
    );
  memtest2_datalfsr_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(22),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(23)
    );
  memtest2_datalfsr_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(30),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(31)
    );
  memtest2_datalfsr_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(17),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(18)
    );
  memtest2_datalfsr_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(16),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(17)
    );
  memtest2_datalfsr_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(24),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(25)
    );
  memcontroller_dnl2_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(1),
      CE => memcontroller_dnl2_1_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_1_FFX_RST,
      O => memcontroller_dnl2(1)
    );
  memcontroller_dnl2_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_1_FFX_RST
    );
  memtest2_datalfsr_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(25),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(26)
    );
  memtest2_datalfsr_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(18),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(19)
    );
  memtest2_datalfsr_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(26),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(27)
    );
  maccontrol_lmacaddr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(11),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_11_FFX_RST,
      O => maccontrol_lmacaddr(11)
    );
  maccontrol_lmacaddr_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_11_FFX_RST
    );
  memcontroller_dnl2_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(3),
      CE => memcontroller_dnl2_3_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_3_FFX_RST,
      O => memcontroller_dnl2(3)
    );
  memcontroller_dnl2_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_3_FFX_RST
    );
  memtest2_datalfsr_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(27),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(28)
    );
  maccontrol_lmacaddr_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(4),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_21_FFY_RST,
      O => maccontrol_lmacaddr(20)
    );
  maccontrol_lmacaddr_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_21_FFY_RST
    );
  memtest2_datalfsr_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(28),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(29)
    );
  maccontrol_lmacaddr_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(5),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_21_FFX_RST,
      O => maccontrol_lmacaddr(21)
    );
  maccontrol_lmacaddr_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_21_FFX_RST
    );
  maccontrol_lmacaddr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(13),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_13_FFX_RST,
      O => maccontrol_lmacaddr(13)
    );
  maccontrol_lmacaddr_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_13_FFX_RST
    );
  memcontroller_dnl2_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(5),
      CE => memcontroller_dnl2_5_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_5_FFX_RST,
      O => memcontroller_dnl2(5)
    );
  memcontroller_dnl2_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_5_FFX_RST
    );
  maccontrol_lmacaddr_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(6),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_23_FFY_RST,
      O => maccontrol_lmacaddr(22)
    );
  maccontrol_lmacaddr_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_23_FFY_RST
    );
  maccontrol_lmacaddr_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(14),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_31_FFY_RST,
      O => maccontrol_lmacaddr(30)
    );
  maccontrol_lmacaddr_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_31_FFY_RST
    );
  maccontrol_lmacaddr_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(9),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_25_FFX_RST,
      O => maccontrol_lmacaddr(25)
    );
  maccontrol_lmacaddr_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_25_FFX_RST
    );
  memcontroller_clknum_0_2_870 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_0_2_BXMUXNOT,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memcontroller_clknum_0_2_FFX_RST,
      O => memcontroller_clknum_0_2
    );
  memcontroller_clknum_0_2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_0_2_FFX_RST
    );
  memtest2_ldata_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(20),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_21_FFY_RST,
      O => memtest2_ldata(20)
    );
  memtest2_ldata_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_21_FFY_RST
    );
  memtest2_ldata_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(21),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_21_FFX_RST,
      O => memtest2_ldata(21)
    );
  memtest2_ldata_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_21_FFX_RST
    );
  memtest2_ldata_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(12),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_13_FFY_RST,
      O => memtest2_ldata(12)
    );
  memtest2_ldata_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_13_FFY_RST
    );
  memtest2_ldata_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(13),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_13_FFX_RST,
      O => memtest2_ldata(13)
    );
  memtest2_ldata_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_13_FFX_RST
    );
  memcontroller_dnl2_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(8),
      CE => memcontroller_dnl2_9_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_9_FFY_RST,
      O => memcontroller_dnl2(8)
    );
  memcontroller_dnl2_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_9_FFY_RST
    );
  memcontroller_dnl2_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(9),
      CE => memcontroller_dnl2_9_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_9_FFX_RST,
      O => memcontroller_dnl2(9)
    );
  memcontroller_dnl2_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_9_FFX_RST
    );
  maccontrol_lmacaddr_34 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(2),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_35_FFY_RST,
      O => maccontrol_lmacaddr(34)
    );
  maccontrol_lmacaddr_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_35_FFY_RST
    );
  maccontrol_lmacaddr_35 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(3),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_35_FFX_RST,
      O => maccontrol_lmacaddr(35)
    );
  maccontrol_lmacaddr_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_35_FFX_RST
    );
  maccontrol_lmacaddr_42 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(10),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_43_FFY_RST,
      O => maccontrol_lmacaddr(42)
    );
  maccontrol_lmacaddr_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_43_FFY_RST
    );
  maccontrol_lmacaddr_43 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(11),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_43_FFX_RST,
      O => maccontrol_lmacaddr(43)
    );
  maccontrol_lmacaddr_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_43_FFX_RST
    );
  maccontrol_lmacaddr_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(3),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_19_FFX_RST,
      O => maccontrol_lmacaddr(19)
    );
  maccontrol_lmacaddr_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_19_FFX_RST
    );
  maccontrol_lmacaddr_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(10),
      CE => maccontrol_n0036,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_27_FFY_RST,
      O => maccontrol_lmacaddr(26)
    );
  maccontrol_lmacaddr_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_27_FFY_RST
    );
  memtest2_ldata_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(17),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_17_FFX_RST,
      O => memtest2_ldata(17)
    );
  memtest2_ldata_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_17_FFX_RST
    );
  maccontrol_lmacaddr_39 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(7),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_39_FFX_RST,
      O => maccontrol_lmacaddr(39)
    );
  maccontrol_lmacaddr_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_39_FFX_RST
    );
  maccontrol_lmacaddr_47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(15),
      CE => maccontrol_n0037,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_47_FFX_RST,
      O => maccontrol_lmacaddr(47)
    );
  maccontrol_lmacaddr_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_47_FFX_RST
    );
  memtest2_ldata_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(27),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_27_FFX_RST,
      O => memtest2_ldata(27)
    );
  memtest2_ldata_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_27_FFX_RST
    );
  memtest2_ldata_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(18),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_19_FFY_RST,
      O => memtest2_ldata(18)
    );
  memtest2_ldata_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_19_FFY_RST
    );
  memtest2_ldata_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(19),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_19_FFX_RST,
      O => memtest2_ldata(19)
    );
  memtest2_ldata_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_19_FFX_RST
    );
  memtest2_ldata_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(28),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_29_FFY_RST,
      O => memtest2_ldata(28)
    );
  memtest2_ldata_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_29_FFY_RST
    );
  memtest2_ldata_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(29),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_ldata_29_FFX_RST,
      O => memtest2_ldata(29)
    );
  memtest2_ldata_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_ldata_29_FFX_RST
    );
  memcontroller_Q2_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(10),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_11_FFY_RST,
      O => q2(10)
    );
  q2_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_11_FFY_RST
    );
  memcontroller_Q2_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(11),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_11_FFX_RST,
      O => q2(11)
    );
  q2_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_11_FFX_RST
    );
  memcontroller_Q2_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(20),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_21_FFY_RST,
      O => q2(20)
    );
  q2_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_21_FFY_RST
    );
  memcontroller_Q2_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(21),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_21_FFX_RST,
      O => q2(21)
    );
  q2_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_21_FFX_RST
    );
  memcontroller_Q2_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(12),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_13_FFY_RST,
      O => q2(12)
    );
  q2_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_13_FFY_RST
    );
  memcontroller_Q2_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(30),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_31_FFY_RST,
      O => q2(30)
    );
  q2_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_31_FFY_RST
    );
  maccontrol_phyaddr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(10),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_11_FFY_RST,
      O => maccontrol_phyaddr(10)
    );
  maccontrol_phyaddr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_11_FFY_RST
    );
  maccontrol_phyaddr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(11),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_11_FFX_RST,
      O => maccontrol_phyaddr(11)
    );
  maccontrol_phyaddr_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_11_FFX_RST
    );
  maccontrol_phyaddr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(12),
      CE => maccontrol_n0031,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phyaddr_13_FFY_RST,
      O => maccontrol_phyaddr(12)
    );
  maccontrol_phyaddr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phyaddr_13_FFY_RST
    );
  memtest_dataw1_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(29),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_29_FFX_RST,
      O => memtest_dataw1(29)
    );
  memtest_dataw1_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_29_FFX_RST
    );
  maccontrol_phydi_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(10),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_11_FFY_RST,
      O => maccontrol_phydi(10)
    );
  maccontrol_phydi_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_11_FFY_RST
    );
  maccontrol_phydi_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(11),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_11_FFX_RST,
      O => maccontrol_phydi(11)
    );
  maccontrol_phydi_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_11_FFX_RST
    );
  maccontrol_phydi_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(13),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_13_FFX_RST,
      O => maccontrol_phydi(13)
    );
  maccontrol_phydi_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_13_FFX_RST
    );
  maccontrol_phydi_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(20),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_21_FFY_RST,
      O => maccontrol_phydi(20)
    );
  maccontrol_phydi_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_21_FFY_RST
    );
  maccontrol_phydi_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(21),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_21_FFX_RST,
      O => maccontrol_phydi(21)
    );
  maccontrol_phydi_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_21_FFX_RST
    );
  maccontrol_phydi_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(22),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_22_FFY_RST,
      O => maccontrol_phydi(22)
    );
  maccontrol_phydi_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_22_FFY_RST
    );
  maccontrol_phydi_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(15),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_15_FFX_RST,
      O => maccontrol_phydi(15)
    );
  maccontrol_phydi_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_15_FFX_RST
    );
  memcontroller_Q2_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(13),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_13_FFX_RST,
      O => q2(13)
    );
  q2_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_13_FFX_RST
    );
  memcontroller_Q2_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(31),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_31_FFX_RST,
      O => q2(31)
    );
  q2_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_31_FFX_RST
    );
  memcontroller_Q2_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(22),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_23_FFY_RST,
      O => q2(22)
    );
  q2_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_23_FFY_RST
    );
  memcontroller_Q2_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(23),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_23_FFX_RST,
      O => q2(23)
    );
  q2_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_23_FFX_RST
    );
  memcontroller_Q2_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(14),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_15_FFY_RST,
      O => q2(14)
    );
  q2_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_15_FFY_RST
    );
  memcontroller_Q2_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(15),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_15_FFX_RST,
      O => q2(15)
    );
  q2_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_15_FFX_RST
    );
  memcontroller_Q2_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(24),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_25_FFY_RST,
      O => q2(24)
    );
  q2_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_25_FFY_RST
    );
  memcontroller_Q2_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(25),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_25_FFX_RST,
      O => q2(25)
    );
  q2_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_25_FFX_RST
    );
  memcontroller_Q2_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(16),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_17_FFY_RST,
      O => q2(16)
    );
  q2_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_17_FFY_RST
    );
  memcontroller_Q2_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(17),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_17_FFX_RST,
      O => q2(17)
    );
  q2_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_17_FFX_RST
    );
  memtest2_lfsr_rst_871 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_n0021,
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_lfsr_rst_FFY_RST,
      O => memtest2_lfsr_rst
    );
  memtest2_lfsr_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_lfsr_rst_FFY_RST
    );
  memcontroller_Q2_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(27),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_27_FFX_RST,
      O => q2(27)
    );
  q2_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_27_FFX_RST
    );
  memcontroller_Q2_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(26),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_27_FFY_RST,
      O => q2(26)
    );
  q2_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_27_FFY_RST
    );
  memcontroller_Q2_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(18),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_19_FFY_RST,
      O => q2(18)
    );
  q2_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_19_FFY_RST
    );
  memcontroller_Q2_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(28),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_29_FFY_RST,
      O => q2(28)
    );
  q2_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_29_FFY_RST
    );
  memcontroller_Q2_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(19),
      CE => memcontroller_n0005,
      CLK => clk,
      SET => GND,
      RST => q2_19_FFX_RST,
      O => q2(19)
    );
  q2_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_19_FFX_RST
    );
  memcontroller_dnl2_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(31),
      CE => memcontroller_dnl2_31_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_31_FFX_RST,
      O => memcontroller_dnl2(31)
    );
  memcontroller_dnl2_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_31_FFX_RST
    );
  memcontroller_dnl2_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(22),
      CE => memcontroller_dnl2_23_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_23_FFY_RST,
      O => memcontroller_dnl2(22)
    );
  memcontroller_dnl2_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_23_FFY_RST
    );
  memcontroller_dnl2_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(23),
      CE => memcontroller_dnl2_23_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_23_FFX_RST,
      O => memcontroller_dnl2(23)
    );
  memcontroller_dnl2_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_23_FFX_RST
    );
  memcontroller_dnl2_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(14),
      CE => memcontroller_dnl2_15_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_15_FFY_RST,
      O => memcontroller_dnl2(14)
    );
  memcontroller_dnl2_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_15_FFY_RST
    );
  memcontroller_dnl2_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(15),
      CE => memcontroller_dnl2_15_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_15_FFX_RST,
      O => memcontroller_dnl2(15)
    );
  memcontroller_dnl2_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_15_FFX_RST
    );
  memtest_dataw1_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(30),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_31_FFY_RST,
      O => memtest_dataw1(30)
    );
  memtest_dataw1_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_31_FFY_RST
    );
  memtest_dataw1_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(31),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_31_FFX_RST,
      O => memtest_dataw1(31)
    );
  memtest_dataw1_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_31_FFX_RST
    );
  memtest_dataw1_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(22),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_23_FFY_RST,
      O => memtest_dataw1(22)
    );
  memtest_dataw1_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_23_FFY_RST
    );
  memtest_dataw1_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(23),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_23_FFX_RST,
      O => memtest_dataw1(23)
    );
  memtest_dataw1_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_23_FFX_RST
    );
  memtest_dataw1_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(14),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_15_FFY_RST,
      O => memtest_dataw1(14)
    );
  memtest_dataw1_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_15_FFY_RST
    );
  memtest_dataw1_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(15),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_15_FFX_RST,
      O => memtest_dataw1(15)
    );
  memtest_dataw1_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_15_FFX_RST
    );
  memcontroller_dnl2_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(24),
      CE => memcontroller_dnl2_25_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_25_FFY_RST,
      O => memcontroller_dnl2(24)
    );
  memcontroller_dnl2_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_25_FFY_RST
    );
  memcontroller_dnl2_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(25),
      CE => memcontroller_dnl2_25_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_25_FFX_RST,
      O => memcontroller_dnl2(25)
    );
  memcontroller_dnl2_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_25_FFX_RST
    );
  memcontroller_dnl2_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(16),
      CE => memcontroller_dnl2_17_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_17_FFY_RST,
      O => memcontroller_dnl2(16)
    );
  memcontroller_dnl2_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_17_FFY_RST
    );
  memtest_dataw1_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(24),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_25_FFY_RST,
      O => memtest_dataw1(24)
    );
  memtest_dataw1_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_25_FFY_RST
    );
  memcontroller_dnl2_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(17),
      CE => memcontroller_dnl2_17_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_17_FFX_RST,
      O => memcontroller_dnl2(17)
    );
  memcontroller_dnl2_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_17_FFX_RST
    );
  memtest2_datain_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(8),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_9_FFY_RST,
      O => memtest2_datain(8)
    );
  memtest2_datain_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_9_FFY_RST
    );
  memtest2_datain_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(9),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_9_FFX_RST,
      O => memtest2_datain(9)
    );
  memtest2_datain_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_9_FFX_RST
    );
  maccontrol_sclkdeltall_872 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_sclkdeltal,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => maccontrol_sclkdeltall_FFY_RST,
      O => maccontrol_sclkdeltall
    );
  maccontrol_sclkdeltall_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_sclkdeltall_FFY_RST
    );
  maccontrol_PHY_status_addrl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyaddr(0),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_addrl_1_FFY_RST,
      O => maccontrol_PHY_status_addrl(0)
    );
  maccontrol_PHY_status_addrl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_addrl_1_FFY_RST
    );
  maccontrol_phydi_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(30),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_31_FFY_RST,
      O => maccontrol_phydi(30)
    );
  maccontrol_phydi_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_31_FFY_RST
    );
  maccontrol_phydi_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(31),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_31_FFX_RST,
      O => maccontrol_phydi(31)
    );
  maccontrol_phydi_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_31_FFX_RST
    );
  maccontrol_phydi_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(16),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_17_FFY_RST,
      O => maccontrol_phydi(16)
    );
  maccontrol_phydi_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_17_FFY_RST
    );
  maccontrol_phydi_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(17),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_17_FFX_RST,
      O => maccontrol_phydi(17)
    );
  maccontrol_phydi_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_17_FFX_RST
    );
  maccontrol_phydi_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(25),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_25_FFX_RST,
      O => maccontrol_phydi(25)
    );
  maccontrol_phydi_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_25_FFX_RST
    );
  maccontrol_phydi_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(19),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_19_FFX_RST,
      O => maccontrol_phydi(19)
    );
  maccontrol_phydi_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_19_FFX_RST
    );
  maccontrol_phydi_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(27),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_27_FFX_RST,
      O => maccontrol_phydi(27)
    );
  maccontrol_phydi_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_27_FFX_RST
    );
  maccontrol_phydi_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(29),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_29_FFX_RST,
      O => maccontrol_phydi(29)
    );
  maccontrol_phydi_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_29_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(1),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_1_FFX_RST,
      O => maccontrol_phystat(1)
    );
  maccontrol_phystat_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_1_FFX_RST
    );
  memtest_dataw1_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(25),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_25_FFX_RST,
      O => memtest_dataw1(25)
    );
  memtest_dataw1_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_25_FFX_RST
    );
  memtest_dataw1_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(16),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_17_FFY_RST,
      O => memtest_dataw1(16)
    );
  memtest_dataw1_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_17_FFY_RST
    );
  memtest_dataw1_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(17),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_17_FFX_RST,
      O => memtest_dataw1(17)
    );
  memtest_dataw1_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_17_FFX_RST
    );
  memcontroller_dnl2_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(26),
      CE => memcontroller_dnl2_27_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_27_FFY_RST,
      O => memcontroller_dnl2(26)
    );
  memcontroller_dnl2_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_27_FFY_RST
    );
  memcontroller_dnl2_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(27),
      CE => memcontroller_dnl2_27_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_27_FFX_RST,
      O => memcontroller_dnl2(27)
    );
  memcontroller_dnl2_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_27_FFX_RST
    );
  memcontroller_dnl2_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(18),
      CE => memcontroller_dnl2_19_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_19_FFY_RST,
      O => memcontroller_dnl2(18)
    );
  memcontroller_dnl2_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_19_FFY_RST
    );
  memcontroller_dnl2_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(19),
      CE => memcontroller_dnl2_19_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_19_FFX_RST,
      O => memcontroller_dnl2(19)
    );
  memcontroller_dnl2_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_19_FFX_RST
    );
  memtest_dataw1_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(26),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_27_FFY_RST,
      O => memtest_dataw1(26)
    );
  memtest_dataw1_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_27_FFY_RST
    );
  memtest_dataw1_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(27),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_27_FFX_RST,
      O => memtest_dataw1(27)
    );
  memtest_dataw1_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_27_FFX_RST
    );
  memtest_dataw1_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(18),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_19_FFY_RST,
      O => memtest_dataw1(18)
    );
  memtest_dataw1_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_19_FFY_RST
    );
  memtest_dataw1_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(19),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_19_FFX_RST,
      O => memtest_dataw1(19)
    );
  memtest_dataw1_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_19_FFX_RST
    );
  memcontroller_dnl2_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(28),
      CE => memcontroller_dnl2_29_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_29_FFY_RST,
      O => memcontroller_dnl2(28)
    );
  memcontroller_dnl2_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_29_FFY_RST
    );
  memcontroller_dnl2_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(29),
      CE => memcontroller_dnl2_29_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_dnl2_29_FFX_RST,
      O => memcontroller_dnl2(29)
    );
  memcontroller_dnl2_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_29_FFX_RST
    );
  memtest_dataw1_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(28),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_29_FFY_RST,
      O => memtest_dataw1(28)
    );
  memtest_dataw1_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_29_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(3),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_3_FFX_RST,
      O => maccontrol_phystat(3)
    );
  maccontrol_phystat_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_3_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(4),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_5_FFY_RST,
      O => maccontrol_phystat(4)
    );
  maccontrol_phystat_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_5_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(5),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_5_FFX_RST,
      O => maccontrol_phystat(5)
    );
  maccontrol_phystat_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_5_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(6),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_7_FFY_RST,
      O => maccontrol_phystat(6)
    );
  maccontrol_phystat_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_7_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(7),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_7_FFX_RST,
      O => maccontrol_phystat(7)
    );
  maccontrol_phystat_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_7_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(8),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_9_FFY_RST,
      O => maccontrol_phystat(8)
    );
  maccontrol_phystat_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_9_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(9),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_9_FFX_RST,
      O => maccontrol_phystat(9)
    );
  maccontrol_phystat_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_9_FFX_RST
    );
  testrx_cs_FFd1_873 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => testrx_cs_FFd1_In,
      CE => VCC,
      CLK => rx_clk_int,
      SET => GND,
      RST => testrx_cs_FFd1_FFY_RST,
      O => testrx_cs_FFd1
    );
  testrx_cs_FFd1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => testrx_cs_FFd1_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(10),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_12_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(11)
    );
  maccontrol_PHY_status_MII_Interface_dreg_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_12_FFY_RST
    );
  memtest2_datain_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(0),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_1_FFY_RST,
      O => memtest2_datain(0)
    );
  memtest2_datain_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_1_FFY_RST
    );
  memtest2_datain_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(1),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_1_FFX_RST,
      O => memtest2_datain(1)
    );
  memtest2_datain_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_1_FFX_RST
    );
  memtest2_datain_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(2),
      CE => memtest2_n00511_O,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_2_FFY_RST,
      O => memtest2_datain(2)
    );
  memtest2_datain_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_2_FFY_RST
    );
  memtest2_datain_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(3),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_3_FFY_RST,
      O => memtest2_datain(3)
    );
  memtest2_datain_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_3_FFY_RST
    );
  memtest2_datain_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(4),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_5_FFY_RST,
      O => memtest2_datain(4)
    );
  memtest2_datain_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_5_FFY_RST
    );
  memtest2_datain_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(5),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_5_FFX_RST,
      O => memtest2_datain(5)
    );
  memtest2_datain_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_5_FFX_RST
    );
  memtest2_datain_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(6),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_7_FFY_RST,
      O => memtest2_datain(6)
    );
  memtest2_datain_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_7_FFY_RST
    );
  memtest2_datain_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q2(7),
      CE => memtest2_n00511_4,
      CLK => clk,
      SET => GND,
      RST => memtest2_datain_7_FFX_RST,
      O => memtest2_datain(7)
    );
  memtest2_datain_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_datain_7_FFX_RST
    );
  maccontrol_din_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(16),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_17_FFX_RST,
      O => maccontrol_din(17)
    );
  maccontrol_din_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_17_FFX_RST
    );
  maccontrol_din_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(23),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_25_FFY_RST,
      O => maccontrol_din(24)
    );
  maccontrol_din_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_25_FFY_RST
    );
  maccontrol_din_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(24),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_25_FFX_RST,
      O => maccontrol_din(25)
    );
  maccontrol_din_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_25_FFX_RST
    );
  maccontrol_din_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(17),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_19_FFY_RST,
      O => maccontrol_din(18)
    );
  maccontrol_din_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_19_FFY_RST
    );
  maccontrol_din_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(18),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_19_FFX_RST,
      O => maccontrol_din(19)
    );
  maccontrol_din_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_19_FFX_RST
    );
  maccontrol_din_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(25),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_27_FFY_RST,
      O => maccontrol_din(26)
    );
  maccontrol_din_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_27_FFY_RST
    );
  maccontrol_din_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(26),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_27_FFX_RST,
      O => maccontrol_din(27)
    );
  maccontrol_din_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_27_FFX_RST
    );
  maccontrol_din_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(27),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_29_FFY_RST,
      O => maccontrol_din(28)
    );
  maccontrol_din_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_29_FFY_RST
    );
  maccontrol_din_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(28),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_29_FFX_RST,
      O => maccontrol_din(29)
    );
  maccontrol_din_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_29_FFX_RST
    );
  maccontrol_PHY_status_din_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(0),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_1_FFY_RST,
      O => maccontrol_PHY_status_din(0)
    );
  maccontrol_PHY_status_din_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_1_FFY_RST
    );
  maccontrol_PHY_status_din_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(1),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_1_FFX_RST,
      O => maccontrol_PHY_status_din(1)
    );
  maccontrol_PHY_status_din_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_1_FFX_RST
    );
  maccontrol_PHY_status_din_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(2),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_3_FFY_RST,
      O => maccontrol_PHY_status_din(2)
    );
  maccontrol_PHY_status_din_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_3_FFY_RST
    );
  maccontrol_PHY_status_din_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(3),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_3_FFX_RST,
      O => maccontrol_PHY_status_din(3)
    );
  maccontrol_PHY_status_din_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_3_FFX_RST
    );
  maccontrol_PHY_status_din_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(4),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_5_FFY_RST,
      O => maccontrol_PHY_status_din(4)
    );
  maccontrol_PHY_status_din_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_5_FFY_RST
    );
  maccontrol_PHY_status_din_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(5),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_5_FFX_RST,
      O => maccontrol_PHY_status_din(5)
    );
  maccontrol_PHY_status_din_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_5_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(12),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_14_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(13)
    );
  maccontrol_PHY_status_MII_Interface_dreg_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_14_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(11),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_12_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(12)
    );
  maccontrol_PHY_status_MII_Interface_dreg_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_12_FFX_RST
    );
  maccontrol_PHY_status_din_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(11),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_11_FFX_RST,
      O => maccontrol_PHY_status_din(11)
    );
  maccontrol_PHY_status_din_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_11_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(13),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_14_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(14)
    );
  maccontrol_PHY_status_MII_Interface_dreg_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_14_FFX_RST
    );
  maccontrol_PHY_status_din_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(13),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_13_FFX_RST,
      O => maccontrol_PHY_status_din(13)
    );
  maccontrol_PHY_status_din_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_13_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(14),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_15_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(15)
    );
  maccontrol_PHY_status_MII_Interface_dreg_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_15_FFY_RST
    );
  maccontrol_PHY_status_din_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(14),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_15_FFY_RST,
      O => maccontrol_PHY_status_din(14)
    );
  maccontrol_PHY_status_din_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_15_FFY_RST
    );
  maccontrol_PHY_status_din_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(15),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_15_FFX_RST,
      O => maccontrol_PHY_status_din(15)
    );
  maccontrol_PHY_status_din_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_15_FFX_RST
    );
  maccontrol_PHY_status_addrl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyaddr(1),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_addrl_1_FFX_RST,
      O => maccontrol_PHY_status_addrl(1)
    );
  maccontrol_PHY_status_addrl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_addrl_1_FFX_RST
    );
  memtest2_datalfsr_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(1),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(2)
    );
  memtest2_datalfsr_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(2),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(3)
    );
  maccontrol_PHY_status_addrl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyaddr(3),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_addrl_3_FFX_RST,
      O => maccontrol_PHY_status_addrl(3)
    );
  maccontrol_PHY_status_addrl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_addrl_3_FFX_RST
    );
  maccontrol_PHY_status_addrl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyaddr(2),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_addrl_3_FFY_RST,
      O => maccontrol_PHY_status_addrl(2)
    );
  maccontrol_PHY_status_addrl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_addrl_3_FFY_RST
    );
  memtest2_datalfsr_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(3),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(4)
    );
  memtest2_datalfsr_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(4),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(5)
    );
  maccontrol_lmacaddr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(1),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_1_FFX_RST,
      O => maccontrol_lmacaddr(1)
    );
  maccontrol_lmacaddr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_1_FFX_RST
    );
  maccontrol_lmacaddr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(0),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_1_FFY_RST,
      O => maccontrol_lmacaddr(0)
    );
  maccontrol_lmacaddr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_1_FFY_RST
    );
  maccontrol_PHY_status_addrl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyaddr(4),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_addrl_4_FFY_RST,
      O => maccontrol_PHY_status_addrl(4)
    );
  maccontrol_PHY_status_addrl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_addrl_4_FFY_RST
    );
  memtest2_datalfsr_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(5),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(6)
    );
  memtest2_datalfsr_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(6),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(7)
    );
  maccontrol_lmacaddr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(3),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_3_FFX_RST,
      O => maccontrol_lmacaddr(3)
    );
  maccontrol_lmacaddr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_3_FFX_RST
    );
  maccontrol_lmacaddr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(2),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_3_FFY_RST,
      O => maccontrol_lmacaddr(2)
    );
  maccontrol_lmacaddr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_3_FFY_RST
    );
  clken_clkcnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => clken_clkcnt_n0000(1),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => clken_n0002,
      O => clken_clkcnt(1)
    );
  memtest2_datalfsr_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(7),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(8)
    );
  clken_clkcnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => clken_clkcnt_0_BXMUXNOT,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => clken_n0002,
      O => clken_clkcnt(0)
    );
  memtest2_datalfsr_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_datalfsr(8),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_datalfsr(9)
    );
  maccontrol_lmacaddr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(4),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_5_FFY_RST,
      O => maccontrol_lmacaddr(4)
    );
  maccontrol_lmacaddr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_5_FFY_RST
    );
  maccontrol_lmacaddr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(5),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_5_FFX_RST,
      O => maccontrol_lmacaddr(5)
    );
  maccontrol_lmacaddr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_5_FFX_RST
    );
  maccontrol_lmacaddr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(6),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_7_FFY_RST,
      O => maccontrol_lmacaddr(6)
    );
  maccontrol_lmacaddr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_7_FFY_RST
    );
  maccontrol_lmacaddr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(7),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_7_FFX_RST,
      O => maccontrol_lmacaddr(7)
    );
  maccontrol_lmacaddr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_7_FFX_RST
    );
  maccontrol_lmacaddr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(8),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_9_FFY_RST,
      O => maccontrol_lmacaddr(8)
    );
  maccontrol_lmacaddr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_9_FFY_RST
    );
  maccontrol_lmacaddr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(9),
      CE => maccontrol_n0035,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lmacaddr_9_FFX_RST,
      O => maccontrol_lmacaddr(9)
    );
  maccontrol_lmacaddr_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lmacaddr_9_FFX_RST
    );
  maccontrol_addr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mshreg_sinlll_83,
      CE => maccontrol_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_addr_1_FFY_RST,
      O => maccontrol_addr(0)
    );
  maccontrol_addr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_addr_1_FFY_RST
    );
  maccontrol_addr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_addr_1_1,
      CE => maccontrol_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_addr_3_FFY_RST,
      O => maccontrol_addr(2)
    );
  maccontrol_addr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_addr_3_FFY_RST
    );
  maccontrol_addr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_addr_0_1,
      CE => maccontrol_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_addr_1_FFX_RST,
      O => maccontrol_addr(1)
    );
  maccontrol_addr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_addr_1_FFX_RST
    );
  maccontrol_addr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_addr(3),
      CE => maccontrol_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_addr_5_FFY_RST,
      O => maccontrol_addr(4)
    );
  maccontrol_addr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_addr_5_FFY_RST
    );
  maccontrol_addr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_addr(2),
      CE => maccontrol_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_addr_3_FFX_RST,
      O => maccontrol_addr(3)
    );
  maccontrol_addr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_addr_3_FFX_RST
    );
  maccontrol_addr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_addr(4),
      CE => maccontrol_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_addr_5_FFX_RST,
      O => maccontrol_addr(5)
    );
  maccontrol_addr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_addr_5_FFX_RST
    );
  memtest_lerr_874 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest_llerr,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest_lerr_FFY_RST,
      O => memtest_lerr
    );
  memtest_lerr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_lerr_FFY_RST
    );
  maccontrol_addr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_addr(5),
      CE => maccontrol_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_addr_7_FFY_RST,
      O => maccontrol_addr(6)
    );
  maccontrol_addr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_addr_7_FFY_RST
    );
  maccontrol_addr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_addr(6),
      CE => maccontrol_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_addr_7_FFX_RST,
      O => maccontrol_addr(7)
    );
  maccontrol_addr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_addr_7_FFX_RST
    );
  maccontrol_lrxbcast_875 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(0),
      CE => maccontrol_n0032,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lrxbcast_FFY_RST,
      O => maccontrol_lrxbcast
    );
  maccontrol_lrxbcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lrxbcast_FFY_RST
    );
  maccontrol_addr_0_1_876 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_Mshreg_sinlll_83,
      CE => maccontrol_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_addr_0_1_FFY_RST,
      O => maccontrol_addr_0_1
    );
  maccontrol_addr_0_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_addr_0_1_FFY_RST
    );
  maccontrol_addr_1_1_877 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_addr_0_1,
      CE => maccontrol_n0010,
      CLK => clk,
      SET => GND,
      RST => maccontrol_addr_1_1_FFY_RST,
      O => maccontrol_addr_1_1
    );
  maccontrol_addr_1_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_addr_1_1_FFY_RST
    );
  memtest_dataw1_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(0),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_1_FFY_RST,
      O => memtest_dataw1(0)
    );
  memtest_dataw1_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_1_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(11),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_11_FFX_RST,
      O => maccontrol_PHY_status_dout(11)
    );
  maccontrol_PHY_status_dout_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_11_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(12),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_13_FFY_RST,
      O => maccontrol_PHY_status_dout(12)
    );
  maccontrol_PHY_status_dout_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_13_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(13),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_13_FFX_RST,
      O => maccontrol_PHY_status_dout(13)
    );
  maccontrol_PHY_status_dout_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_13_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(14),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_15_FFY_RST,
      O => maccontrol_PHY_status_dout(14)
    );
  maccontrol_PHY_status_dout_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_15_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_DOUT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(15),
      CE => maccontrol_PHY_status_MII_Interface_n0016,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_dout_15_FFX_RST,
      O => maccontrol_PHY_status_dout(15)
    );
  maccontrol_PHY_status_dout_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_dout_15_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(10),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_11_FFY_RST,
      O => maccontrol_phystat(10)
    );
  maccontrol_phystat_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_11_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(11),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_11_FFX_RST,
      O => maccontrol_phystat(11)
    );
  maccontrol_phystat_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_11_FFX_RST
    );
  memtest_dataw1_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(1),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_1_FFX_RST,
      O => memtest_dataw1(1)
    );
  memtest_dataw1_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_1_FFX_RST
    );
  memtest_dataw1_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(2),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_3_FFY_RST,
      O => memtest_dataw1(2)
    );
  memtest_dataw1_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_3_FFY_RST
    );
  memtest_dataw1_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(3),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_3_FFX_RST,
      O => memtest_dataw1(3)
    );
  memtest_dataw1_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_3_FFX_RST
    );
  memtest_dataw1_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(4),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_5_FFY_RST,
      O => memtest_dataw1(4)
    );
  memtest_dataw1_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_5_FFY_RST
    );
  memtest_dataw1_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(5),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_5_FFX_RST,
      O => memtest_dataw1(5)
    );
  memtest_dataw1_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_5_FFX_RST
    );
  memtest_dataw1_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(6),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_7_FFY_RST,
      O => memtest_dataw1(6)
    );
  memtest_dataw1_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_7_FFY_RST
    );
  memtest_dataw1_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(7),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_7_FFX_RST,
      O => memtest_dataw1(7)
    );
  memtest_dataw1_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_7_FFX_RST
    );
  memtest_dataw1_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(8),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_9_FFY_RST,
      O => memtest_dataw1(8)
    );
  memtest_dataw1_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_9_FFY_RST
    );
  memtest_dataw1_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => d1(9),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_dataw1_9_FFX_RST,
      O => memtest_dataw1(9)
    );
  memtest_dataw1_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_dataw1_9_FFX_RST
    );
  maccontrol_phydi_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(0),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_1_FFY_RST,
      O => maccontrol_phydi(0)
    );
  maccontrol_phydi_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_1_FFY_RST
    );
  maccontrol_phydi_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(1),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_1_FFX_RST,
      O => maccontrol_phydi(1)
    );
  maccontrol_phydi_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_1_FFX_RST
    );
  maccontrol_phydi_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(2),
      CE => maccontrol_n0013,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_2_FFY_RST,
      O => maccontrol_phydi(2)
    );
  maccontrol_phydi_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_2_FFY_RST
    );
  maccontrol_phydi_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(3),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_3_FFY_RST,
      O => maccontrol_phydi(3)
    );
  maccontrol_phydi_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_3_FFY_RST
    );
  maccontrol_din_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(9),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_11_FFY_RST,
      O => maccontrol_din(10)
    );
  maccontrol_din_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_11_FFY_RST
    );
  maccontrol_phydi_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(4),
      CE => maccontrol_n00131_1,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phydi_5_FFY_RST,
      O => maccontrol_phydi(4)
    );
  maccontrol_phydi_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phydi_5_FFY_RST
    );
  maccontrol_din_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(4),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_5_FFX_RST,
      O => maccontrol_din(5)
    );
  maccontrol_din_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_5_FFX_RST
    );
  maccontrol_din_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(6),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_7_FFX_RST,
      O => maccontrol_din(7)
    );
  maccontrol_din_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_7_FFX_RST
    );
  maccontrol_din_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(7),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_9_FFY_RST,
      O => maccontrol_din(8)
    );
  maccontrol_din_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_9_FFY_RST
    );
  maccontrol_din_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(8),
      CE => maccontrol_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_din_9_FFX_RST,
      O => maccontrol_din(9)
    );
  maccontrol_din_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_din_9_FFX_RST
    );
  memtest2_addrlfsr_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(1),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(2)
    );
  memtest2_addrlfsr_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(3),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(4)
    );
  memtest2_addrlfsr_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(2),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(3)
    );
  memtest2_addrlfsr_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(4),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(5)
    );
  memtest2_addrlfsr_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(6),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(7)
    );
  clken_clken : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => clken_lclken,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => clkslen_FFY_RST,
      O => clkslen
    );
  clkslen_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => clkslen_FFY_RST
    );
  memtest2_addrlfsr_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(8),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(9)
    );
  maccontrol_PHY_status_din_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(6),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_7_FFY_RST,
      O => maccontrol_PHY_status_din(6)
    );
  maccontrol_PHY_status_din_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_7_FFY_RST
    );
  maccontrol_PHY_status_din_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(7),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_7_FFX_RST,
      O => maccontrol_PHY_status_din(7)
    );
  maccontrol_PHY_status_din_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_7_FFX_RST
    );
  maccontrol_PHY_status_din_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(8),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_9_FFY_RST,
      O => maccontrol_PHY_status_din(8)
    );
  maccontrol_PHY_status_din_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_9_FFY_RST
    );
  maccontrol_PHY_status_din_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phydi(9),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_din_9_FFX_RST,
      O => maccontrol_PHY_status_din(9)
    );
  maccontrol_PHY_status_din_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_din_9_FFX_RST
    );
  maccontrol_sclkdeltal_878 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_sclkdelta,
      CE => maccontrol_N30273,
      CLK => clk,
      SET => GND,
      RST => maccontrol_sclkdeltal_FFY_RST,
      O => maccontrol_sclkdeltal
    );
  maccontrol_sclkdeltal_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_sclkdeltal_FFY_RST
    );
  memtest2_addrlfsr_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(9),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(10)
    );
  memtest2_addrlfsr_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(10),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(11)
    );
  memtest2_addrlfsr_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(12),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(13)
    );
  memtest2_addrlfsr_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(13),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(14)
    );
  memtest2_addrlfsr_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(14),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => memtest2_lfsr_rst,
      O => memtest2_addrlfsr(15)
    );
  memcontroller_oel_879 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel_BYMUXNOT,
      CE => memcontroller_oel_CEMUXNOT,
      CLK => clk,
      SET => GND,
      RST => memcontroller_oel_FFY_RST,
      O => memcontroller_oel
    );
  memcontroller_oel_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_oel_FFY_RST
    );
  maccontrol_lrxallf_880 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => maccontrol_din(0),
      CE => maccontrol_n0234,
      CLK => clk,
      SET => maccontrol_lrxallf_FFY_SET,
      RST => GND,
      O => maccontrol_lrxallf
    );
  maccontrol_lrxallf_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => maccontrol_lrxallf_FFY_SET
    );
  memtest2_deql_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_deq(1),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_deql_0_FFY_RST,
      O => memtest2_deql(1)
    );
  memtest2_deql_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_deql_0_FFY_RST
    );
  memtest2_deql_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_deq_0_rt,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_deql_0_FFX_RST,
      O => memtest2_deql(0)
    );
  memtest2_deql_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_deql_0_FFX_RST
    );
  txsim_ltxd_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_ramout(0),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => txsim_ltxd_1_FFY_RST,
      O => txsim_ltxd(0)
    );
  txsim_ltxd_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txsim_ltxd_1_FFY_RST
    );
  txsim_ltxd_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_ramout(1),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => txsim_ltxd_1_FFX_RST,
      O => txsim_ltxd(1)
    );
  txsim_ltxd_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txsim_ltxd_1_FFX_RST
    );
  txsim_ltxd_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_ramout(2),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => txsim_ltxd_3_FFY_RST,
      O => txsim_ltxd(2)
    );
  txsim_ltxd_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txsim_ltxd_3_FFY_RST
    );
  txsim_ltxd_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_ramout(3),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => txsim_ltxd_3_FFX_RST,
      O => txsim_ltxd(3)
    );
  txsim_ltxd_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txsim_ltxd_3_FFX_RST
    );
  txsim_ltxd_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_ramout(4),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => txsim_ltxd_5_FFY_RST,
      O => txsim_ltxd(4)
    );
  txsim_ltxd_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txsim_ltxd_5_FFY_RST
    );
  txsim_ltxd_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_ramout(5),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => txsim_ltxd_5_FFX_RST,
      O => txsim_ltxd(5)
    );
  txsim_ltxd_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txsim_ltxd_5_FFX_RST
    );
  txsim_ltxd_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_ramout(6),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => txsim_ltxd_7_FFY_RST,
      O => txsim_ltxd(6)
    );
  txsim_ltxd_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txsim_ltxd_7_FFY_RST
    );
  txsim_ltxd_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txsim_ramout(7),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => txsim_ltxd_7_FFX_RST,
      O => txsim_ltxd(7)
    );
  txsim_ltxd_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txsim_ltxd_7_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(0),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_2_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(1)
    );
  maccontrol_PHY_status_MII_Interface_dreg_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_2_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(1),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_2_FFX_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(2)
    );
  maccontrol_PHY_status_MII_Interface_dreg_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_2_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(2),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_4_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(3)
    );
  maccontrol_PHY_status_MII_Interface_dreg_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_4_FFY_RST
    );
  maccontrol_PHY_status_MII_Interface_dreg_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_dreg(4),
      CE => maccontrol_PHY_status_MII_Interface_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_dreg_6_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_dreg(5)
    );
  maccontrol_PHY_status_MII_Interface_dreg_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_MII_Interface_dreg_6_FFY_RST
    );
  memtest2_MA_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(0),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_1_FFY_RST,
      O => addr2(0)
    );
  addr2_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_1_FFY_RST
    );
  memtest2_MA_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(1),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_1_FFX_RST,
      O => addr2(1)
    );
  addr2_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_1_FFX_RST
    );
  memtest2_MA_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(2),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_3_FFY_RST,
      O => addr2(2)
    );
  addr2_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_3_FFY_RST
    );
  memtest2_MA_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(3),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_3_FFX_RST,
      O => addr2(3)
    );
  addr2_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_3_FFX_RST
    );
  memtest2_MA_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(4),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_5_FFY_RST,
      O => addr2(4)
    );
  addr2_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_5_FFY_RST
    );
  memtest2_MA_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(5),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_5_FFX_RST,
      O => addr2(5)
    );
  addr2_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_5_FFX_RST
    );
  memtest2_MA_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(6),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_7_FFY_RST,
      O => addr2(6)
    );
  addr2_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_7_FFY_RST
    );
  memtest2_MA_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(7),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_7_FFX_RST,
      O => addr2(7)
    );
  addr2_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_7_FFX_RST
    );
  memtest2_MWE : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_cs(0),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => mwe2_FFY_RST,
      O => mwe2
    );
  mwe2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mwe2_FFY_RST
    );
  memtest2_MA_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(8),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_9_FFY_RST,
      O => addr2(8)
    );
  addr2_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_9_FFY_RST
    );
  maccontrol_PHY_status_rwl_881 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_phyaddr(5),
      CE => maccontrol_PHY_status_n0011,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_rwl_FFY_RST,
      O => maccontrol_PHY_status_rwl
    );
  maccontrol_PHY_status_rwl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_PHY_status_rwl_FFY_RST
    );
  memtest2_MA_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(9),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_9_FFX_RST,
      O => addr2(9)
    );
  addr2_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_9_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(13),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_29_FFX_RST,
      O => maccontrol_phystat(29)
    );
  maccontrol_phystat_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_29_FFX_RST
    );
  memtest_addrcntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(9),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_9_FFX_RST,
      O => memtest_addrcntl(9)
    );
  memtest_addrcntl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_9_FFX_RST
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd2_882 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_MII_Interface_cs_FFd2_In,
      CE => clkslen,
      CLK => clk,
      SET => GND,
      RST => maccontrol_PHY_status_MII_Interface_cs_FFd2_FFY_RST,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd2
    );
  maccontrol_PHY_status_MII_Interface_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => maccontrol_PHY_status_MII_Interface_cs_FFd2_FFY_RST
    );
  maccontrol_lrxucast_883 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_din(0),
      CE => maccontrol_n0034,
      CLK => clk,
      SET => GND,
      RST => maccontrol_lrxucast_FFY_RST,
      O => maccontrol_lrxucast
    );
  maccontrol_lrxucast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_lrxucast_FFY_RST
    );
  memtest2_laddr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(0),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_1_FFY_RST,
      O => memtest2_laddr(0)
    );
  memtest2_laddr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_1_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(12),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_13_FFY_RST,
      O => maccontrol_phystat(12)
    );
  maccontrol_phystat_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_13_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(4),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_21_FFY_RST,
      O => maccontrol_phystat(20)
    );
  maccontrol_phystat_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_21_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(5),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_21_FFX_RST,
      O => maccontrol_phystat(21)
    );
  maccontrol_phystat_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_21_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(13),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_13_FFX_RST,
      O => maccontrol_phystat(13)
    );
  maccontrol_phystat_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_13_FFX_RST
    );
  memtest_addrcntl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(0),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_1_FFY_RST,
      O => memtest_addrcntl(0)
    );
  memtest_addrcntl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_1_FFY_RST
    );
  memtest_addrcntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(1),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_1_FFX_RST,
      O => memtest_addrcntl(1)
    );
  memtest_addrcntl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_1_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(6),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_23_FFY_RST,
      O => maccontrol_phystat(22)
    );
  maccontrol_phystat_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_23_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(7),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_23_FFX_RST,
      O => maccontrol_phystat(23)
    );
  maccontrol_phystat_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_23_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(14),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_31_FFY_RST,
      O => maccontrol_phystat(30)
    );
  maccontrol_phystat_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_31_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(15),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_31_FFX_RST,
      O => maccontrol_phystat(31)
    );
  maccontrol_phystat_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_31_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(14),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_15_FFY_RST,
      O => maccontrol_phystat(14)
    );
  maccontrol_phystat_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_15_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(15),
      CE => maccontrol_PHY_status_n0019,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_15_FFX_RST,
      O => maccontrol_phystat(15)
    );
  maccontrol_phystat_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_15_FFX_RST
    );
  memtest_addrcntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(2),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_3_FFY_RST,
      O => memtest_addrcntl(2)
    );
  memtest_addrcntl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_3_FFY_RST
    );
  memtest_addrcntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(3),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_3_FFX_RST,
      O => memtest_addrcntl(3)
    );
  memtest_addrcntl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_3_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(8),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_25_FFY_RST,
      O => maccontrol_phystat(24)
    );
  maccontrol_phystat_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_25_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(0),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_17_FFY_RST,
      O => maccontrol_phystat(16)
    );
  maccontrol_phystat_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_17_FFY_RST
    );
  memtest2_laddr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(1),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_1_FFX_RST,
      O => memtest2_laddr(1)
    );
  memtest2_laddr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_1_FFX_RST
    );
  memtest2_laddr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(3),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_3_FFX_RST,
      O => memtest2_laddr(3)
    );
  memtest2_laddr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_3_FFX_RST
    );
  memtest2_laddr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(10),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_11_FFY_RST,
      O => memtest2_laddr(10)
    );
  memtest2_laddr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_11_FFY_RST
    );
  memtest2_laddr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(11),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_11_FFX_RST,
      O => memtest2_laddr(11)
    );
  memtest2_laddr_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_11_FFX_RST
    );
  memtest2_laddr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(5),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_5_FFX_RST,
      O => memtest2_laddr(5)
    );
  memtest2_laddr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_5_FFX_RST
    );
  memtest2_laddr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(13),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_13_FFX_RST,
      O => memtest2_laddr(13)
    );
  memtest2_laddr_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_13_FFX_RST
    );
  memtest2_laddr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(6),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_7_FFY_RST,
      O => memtest2_laddr(6)
    );
  memtest2_laddr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_7_FFY_RST
    );
  memtest2_laddr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(7),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_7_FFX_RST,
      O => memtest2_laddr(7)
    );
  memtest2_laddr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_7_FFX_RST
    );
  memtest2_laddr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(15),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_15_FFX_RST,
      O => memtest2_laddr(15)
    );
  memtest2_laddr_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_15_FFX_RST
    );
  memtest2_laddr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(8),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_9_FFY_RST,
      O => memtest2_laddr(8)
    );
  memtest2_laddr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_9_FFY_RST
    );
  memtest2_laddr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_addrlfsr(9),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memtest2_laddr_9_FFX_RST,
      O => memtest2_laddr(9)
    );
  memtest2_laddr_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest2_laddr_9_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(9),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_25_FFX_RST,
      O => maccontrol_phystat(25)
    );
  maccontrol_phystat_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_25_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(1),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_17_FFX_RST,
      O => maccontrol_phystat(17)
    );
  maccontrol_phystat_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_17_FFX_RST
    );
  memtest_addrcntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(4),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_5_FFY_RST,
      O => memtest_addrcntl(4)
    );
  memtest_addrcntl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_5_FFY_RST
    );
  memtest_addrcntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(5),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_5_FFX_RST,
      O => memtest_addrcntl(5)
    );
  memtest_addrcntl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_5_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(10),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_27_FFY_RST,
      O => maccontrol_phystat(26)
    );
  maccontrol_phystat_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_27_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(11),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_27_FFX_RST,
      O => maccontrol_phystat(27)
    );
  maccontrol_phystat_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_27_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(2),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_19_FFY_RST,
      O => maccontrol_phystat(18)
    );
  maccontrol_phystat_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_19_FFY_RST
    );
  maccontrol_PHY_status_PHYSTAT_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(3),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_19_FFX_RST,
      O => maccontrol_phystat(19)
    );
  maccontrol_phystat_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_19_FFX_RST
    );
  memtest_addrcntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(6),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_7_FFY_RST,
      O => memtest_addrcntl(6)
    );
  memtest_addrcntl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_7_FFY_RST
    );
  memtest_addrcntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(7),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_7_FFX_RST,
      O => memtest_addrcntl(7)
    );
  memtest_addrcntl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_7_FFX_RST
    );
  maccontrol_PHY_status_PHYSTAT_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => maccontrol_PHY_status_dout(12),
      CE => maccontrol_PHY_status_n0020,
      CLK => clk,
      SET => GND,
      RST => maccontrol_phystat_29_FFY_RST,
      O => maccontrol_phystat(28)
    );
  maccontrol_phystat_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => maccontrol_phystat_29_FFY_RST
    );
  memtest_addrcntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr1(8),
      CE => clken1,
      CLK => clk,
      SET => GND,
      RST => memtest_addrcntl_9_FFY_RST,
      O => memtest_addrcntl(8)
    );
  memtest_addrcntl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memtest_addrcntl_9_FFY_RST
    );
  memcontroller_clknum_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_1_BYMUXNOT,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memcontroller_clknum_1_FFY_RST,
      O => memcontroller_clknum(0)
    );
  memcontroller_clknum_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_1_FFY_RST
    );
  memcontroller_clknum_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_n0001(1),
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => memcontroller_clknum_1_FFX_RST,
      O => memcontroller_clknum(1)
    );
  memcontroller_clknum_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_1_FFX_RST
    );
  memtest2_MD_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(1),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_1_FFY_RST,
      O => d2(1)
    );
  d2_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_1_FFY_RST
    );
  memtest2_MD_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(2),
      CE => memtest2_n0116,
      CLK => clk,
      SET => GND,
      RST => d2_2_FFY_RST,
      O => d2(2)
    );
  d2_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_2_FFY_RST
    );
  memtest2_MD_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(4),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_5_FFY_RST,
      O => d2(4)
    );
  d2_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_5_FFY_RST
    );
  memtest2_MD_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(5),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_5_FFX_RST,
      O => d2(5)
    );
  d2_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_5_FFX_RST
    );
  clken_lclken_884 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => clken_lclken_LOGIC_ONE,
      CE => VCC,
      CLK => clk,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => clken_n0005,
      O => clken_lclken
    );
  memtest2_MD_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(6),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_7_FFY_RST,
      O => d2(6)
    );
  d2_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_7_FFY_RST
    );
  memtest2_MD_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(7),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_7_FFX_RST,
      O => d2(7)
    );
  d2_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_7_FFX_RST
    );
  memtest2_MD_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(8),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_9_FFY_RST,
      O => d2(8)
    );
  d2_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_9_FFY_RST
    );
  memtest2_MD_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_ldata(9),
      CE => memtest2_n01161_1,
      CLK => clk,
      SET => GND,
      RST => d2_9_FFX_RST,
      O => d2(9)
    );
  d2_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => d2_9_FFX_RST
    );
  memtest2_MA_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(10),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_11_FFY_RST,
      O => addr2(10)
    );
  addr2_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_11_FFY_RST
    );
  memtest2_MA_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memtest2_laddr(11),
      CE => memcontroller_Ker256691_O,
      CLK => clk,
      SET => GND,
      RST => addr2_11_FFX_RST,
      O => addr2(11)
    );
  addr2_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr2_11_FFX_RST
    );
  CLKFB_BUF : X_CKBUF
    port map (
      I => CLKFB,
      O => CLKFB_IBUFG
    );
  CLKIN_BUF : X_CKBUF
    port map (
      I => CLKIN,
      O => CLKIN_IBUFG
    );
  IFCLK_BUF : X_CKBUF
    port map (
      I => IFCLK,
      O => IFCLK_IBUFG
    );
  RX_CLK_BUF : X_CKBUF
    port map (
      I => RX_CLK,
      O => RX_CLK_IBUFG
    );
  ifclk_bufg_BUF : X_CKBUF
    port map (
      I => ifclk_to_bufg,
      O => ifclk_int
    );
  rx_clk_bufg_BUF : X_CKBUF
    port map (
      I => rx_clk_to_bufg,
      O => rx_clk_int
    );
  clk_bufg_BUF : X_CKBUF
    port map (
      I => clk_to_bufg,
      O => clk
    );
  PWR_VCC_0_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_0_FROM
    );
  PWR_VCC_0_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_0_GROM
    );
  PWR_VCC_0_XUSED : X_BUF
    port map (
      I => PWR_VCC_0_FROM,
      O => GLOBAL_LOGIC1
    );
  PWR_VCC_0_YUSED : X_BUF
    port map (
      I => PWR_VCC_0_GROM,
      O => GLOBAL_LOGIC0_67
    );
  PWR_VCC_1_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_1_FROM
    );
  PWR_VCC_1_XUSED : X_BUF
    port map (
      I => PWR_VCC_1_FROM,
      O => GLOBAL_LOGIC1_0
    );
  PWR_VCC_2_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_2_FROM
    );
  PWR_VCC_2_XUSED : X_BUF
    port map (
      I => PWR_VCC_2_FROM,
      O => GLOBAL_LOGIC1_1
    );
  PWR_VCC_3_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_3_FROM
    );
  PWR_VCC_3_XUSED : X_BUF
    port map (
      I => PWR_VCC_3_FROM,
      O => GLOBAL_LOGIC1_2
    );
  PWR_VCC_4_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_4_FROM
    );
  PWR_VCC_4_XUSED : X_BUF
    port map (
      I => PWR_VCC_4_FROM,
      O => GLOBAL_LOGIC1_3
    );
  PWR_VCC_5_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_5_FROM
    );
  PWR_VCC_5_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_5_GROM
    );
  PWR_VCC_5_XUSED : X_BUF
    port map (
      I => PWR_VCC_5_FROM,
      O => GLOBAL_LOGIC1_4
    );
  PWR_VCC_5_YUSED : X_BUF
    port map (
      I => PWR_VCC_5_GROM,
      O => GLOBAL_LOGIC0_58
    );
  PWR_VCC_6_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_6_FROM
    );
  PWR_VCC_6_XUSED : X_BUF
    port map (
      I => PWR_VCC_6_FROM,
      O => GLOBAL_LOGIC1_5
    );
  PWR_VCC_7_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_7_FROM
    );
  PWR_VCC_7_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_7_GROM
    );
  PWR_VCC_7_XUSED : X_BUF
    port map (
      I => PWR_VCC_7_FROM,
      O => GLOBAL_LOGIC1_6
    );
  PWR_VCC_7_YUSED : X_BUF
    port map (
      I => PWR_VCC_7_GROM,
      O => GLOBAL_LOGIC0_57
    );
  PWR_VCC_8_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_8_FROM
    );
  PWR_VCC_8_XUSED : X_BUF
    port map (
      I => PWR_VCC_8_FROM,
      O => GLOBAL_LOGIC1_7
    );
  PWR_VCC_9_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_9_FROM
    );
  PWR_VCC_9_XUSED : X_BUF
    port map (
      I => PWR_VCC_9_FROM,
      O => GLOBAL_LOGIC1_8
    );
  PWR_VCC_10_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_10_FROM
    );
  PWR_VCC_10_XUSED : X_BUF
    port map (
      I => PWR_VCC_10_FROM,
      O => GLOBAL_LOGIC1_9
    );
  PWR_VCC_11_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_11_FROM
    );
  PWR_VCC_11_XUSED : X_BUF
    port map (
      I => PWR_VCC_11_FROM,
      O => GLOBAL_LOGIC1_10
    );
  PWR_VCC_12_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_12_FROM
    );
  PWR_VCC_12_XUSED : X_BUF
    port map (
      I => PWR_VCC_12_FROM,
      O => GLOBAL_LOGIC1_11
    );
  PWR_VCC_13_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_13_FROM
    );
  PWR_VCC_13_XUSED : X_BUF
    port map (
      I => PWR_VCC_13_FROM,
      O => GLOBAL_LOGIC1_12
    );
  PWR_VCC_14_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_14_FROM
    );
  PWR_VCC_14_XUSED : X_BUF
    port map (
      I => PWR_VCC_14_FROM,
      O => GLOBAL_LOGIC1_13
    );
  PWR_VCC_15_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_15_FROM
    );
  PWR_VCC_15_XUSED : X_BUF
    port map (
      I => PWR_VCC_15_FROM,
      O => GLOBAL_LOGIC1_14
    );
  PWR_VCC_16_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_16_FROM
    );
  PWR_VCC_16_XUSED : X_BUF
    port map (
      I => PWR_VCC_16_FROM,
      O => GLOBAL_LOGIC1_15
    );
  PWR_VCC_17_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_17_FROM
    );
  PWR_VCC_17_XUSED : X_BUF
    port map (
      I => PWR_VCC_17_FROM,
      O => GLOBAL_LOGIC1_16
    );
  PWR_VCC_18_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_18_FROM
    );
  PWR_VCC_18_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_18_GROM
    );
  PWR_VCC_18_XUSED : X_BUF
    port map (
      I => PWR_VCC_18_FROM,
      O => GLOBAL_LOGIC1_17
    );
  PWR_VCC_18_YUSED : X_BUF
    port map (
      I => PWR_VCC_18_GROM,
      O => GLOBAL_LOGIC0_51
    );
  PWR_VCC_19_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_19_FROM
    );
  PWR_VCC_19_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_19_GROM
    );
  PWR_VCC_19_XUSED : X_BUF
    port map (
      I => PWR_VCC_19_FROM,
      O => GLOBAL_LOGIC1_18
    );
  PWR_VCC_19_YUSED : X_BUF
    port map (
      I => PWR_VCC_19_GROM,
      O => GLOBAL_LOGIC0_50
    );
  PWR_VCC_20_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_20_FROM
    );
  PWR_VCC_20_XUSED : X_BUF
    port map (
      I => PWR_VCC_20_FROM,
      O => GLOBAL_LOGIC1_19
    );
  PWR_VCC_21_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_21_FROM
    );
  PWR_VCC_21_XUSED : X_BUF
    port map (
      I => PWR_VCC_21_FROM,
      O => GLOBAL_LOGIC1_20
    );
  PWR_VCC_22_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_22_FROM
    );
  PWR_VCC_22_XUSED : X_BUF
    port map (
      I => PWR_VCC_22_FROM,
      O => GLOBAL_LOGIC1_21
    );
  PWR_VCC_23_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_23_FROM
    );
  PWR_VCC_23_XUSED : X_BUF
    port map (
      I => PWR_VCC_23_FROM,
      O => GLOBAL_LOGIC1_22
    );
  PWR_VCC_24_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_24_FROM
    );
  PWR_VCC_24_XUSED : X_BUF
    port map (
      I => PWR_VCC_24_FROM,
      O => GLOBAL_LOGIC1_23
    );
  PWR_VCC_25_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_25_FROM
    );
  PWR_VCC_25_XUSED : X_BUF
    port map (
      I => PWR_VCC_25_FROM,
      O => GLOBAL_LOGIC1_24
    );
  PWR_VCC_26_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_26_FROM
    );
  PWR_VCC_26_XUSED : X_BUF
    port map (
      I => PWR_VCC_26_FROM,
      O => GLOBAL_LOGIC1_25
    );
  PWR_VCC_27_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_27_FROM
    );
  PWR_VCC_27_XUSED : X_BUF
    port map (
      I => PWR_VCC_27_FROM,
      O => GLOBAL_LOGIC1_26
    );
  PWR_VCC_28_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_28_FROM
    );
  PWR_VCC_28_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_28_GROM
    );
  PWR_VCC_28_XUSED : X_BUF
    port map (
      I => PWR_VCC_28_FROM,
      O => GLOBAL_LOGIC1_27
    );
  PWR_VCC_28_YUSED : X_BUF
    port map (
      I => PWR_VCC_28_GROM,
      O => GLOBAL_LOGIC0_47
    );
  PWR_VCC_29_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_29_FROM
    );
  PWR_VCC_29_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_29_GROM
    );
  PWR_VCC_29_XUSED : X_BUF
    port map (
      I => PWR_VCC_29_FROM,
      O => GLOBAL_LOGIC1_28
    );
  PWR_VCC_29_YUSED : X_BUF
    port map (
      I => PWR_VCC_29_GROM,
      O => GLOBAL_LOGIC0_45
    );
  PWR_VCC_30_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_30_FROM
    );
  PWR_VCC_30_XUSED : X_BUF
    port map (
      I => PWR_VCC_30_FROM,
      O => GLOBAL_LOGIC1_29
    );
  PWR_VCC_31_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_31_FROM
    );
  PWR_VCC_31_XUSED : X_BUF
    port map (
      I => PWR_VCC_31_FROM,
      O => GLOBAL_LOGIC1_30
    );
  PWR_VCC_32_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_32_FROM
    );
  PWR_VCC_32_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_32_GROM
    );
  PWR_VCC_32_XUSED : X_BUF
    port map (
      I => PWR_VCC_32_FROM,
      O => GLOBAL_LOGIC1_31
    );
  PWR_VCC_32_YUSED : X_BUF
    port map (
      I => PWR_VCC_32_GROM,
      O => GLOBAL_LOGIC0_41
    );
  PWR_VCC_33_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_33_FROM
    );
  PWR_VCC_33_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_33_GROM
    );
  PWR_VCC_33_XUSED : X_BUF
    port map (
      I => PWR_VCC_33_FROM,
      O => GLOBAL_LOGIC1_32
    );
  PWR_VCC_33_YUSED : X_BUF
    port map (
      I => PWR_VCC_33_GROM,
      O => GLOBAL_LOGIC0_40
    );
  PWR_VCC_34_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_34_FROM
    );
  PWR_VCC_34_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_34_GROM
    );
  PWR_VCC_34_XUSED : X_BUF
    port map (
      I => PWR_VCC_34_FROM,
      O => GLOBAL_LOGIC1_33
    );
  PWR_VCC_34_YUSED : X_BUF
    port map (
      I => PWR_VCC_34_GROM,
      O => GLOBAL_LOGIC0_39
    );
  PWR_VCC_35_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_35_FROM
    );
  PWR_VCC_35_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_35_GROM
    );
  PWR_VCC_35_XUSED : X_BUF
    port map (
      I => PWR_VCC_35_FROM,
      O => GLOBAL_LOGIC1_34
    );
  PWR_VCC_35_YUSED : X_BUF
    port map (
      I => PWR_VCC_35_GROM,
      O => GLOBAL_LOGIC0_36
    );
  PWR_VCC_36_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_36_FROM
    );
  PWR_VCC_36_XUSED : X_BUF
    port map (
      I => PWR_VCC_36_FROM,
      O => GLOBAL_LOGIC1_35
    );
  PWR_VCC_37_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_37_FROM
    );
  PWR_VCC_37_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_37_GROM
    );
  PWR_VCC_37_XUSED : X_BUF
    port map (
      I => PWR_VCC_37_FROM,
      O => GLOBAL_LOGIC1_36
    );
  PWR_VCC_37_YUSED : X_BUF
    port map (
      I => PWR_VCC_37_GROM,
      O => GLOBAL_LOGIC0_34
    );
  PWR_VCC_38_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_38_FROM
    );
  PWR_VCC_38_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_38_GROM
    );
  PWR_VCC_38_XUSED : X_BUF
    port map (
      I => PWR_VCC_38_FROM,
      O => GLOBAL_LOGIC1_37
    );
  PWR_VCC_38_YUSED : X_BUF
    port map (
      I => PWR_VCC_38_GROM,
      O => GLOBAL_LOGIC0_32
    );
  PWR_VCC_39_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_39_FROM
    );
  PWR_VCC_39_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_39_GROM
    );
  PWR_VCC_39_XUSED : X_BUF
    port map (
      I => PWR_VCC_39_FROM,
      O => GLOBAL_LOGIC1_38
    );
  PWR_VCC_39_YUSED : X_BUF
    port map (
      I => PWR_VCC_39_GROM,
      O => GLOBAL_LOGIC0_30
    );
  PWR_VCC_40_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_40_FROM
    );
  PWR_VCC_40_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_40_GROM
    );
  PWR_VCC_40_XUSED : X_BUF
    port map (
      I => PWR_VCC_40_FROM,
      O => GLOBAL_LOGIC1_39
    );
  PWR_VCC_40_YUSED : X_BUF
    port map (
      I => PWR_VCC_40_GROM,
      O => GLOBAL_LOGIC0_29
    );
  PWR_VCC_41_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_41_FROM
    );
  PWR_VCC_41_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_41_GROM
    );
  PWR_VCC_41_XUSED : X_BUF
    port map (
      I => PWR_VCC_41_FROM,
      O => GLOBAL_LOGIC1_40
    );
  PWR_VCC_41_YUSED : X_BUF
    port map (
      I => PWR_VCC_41_GROM,
      O => GLOBAL_LOGIC0_28
    );
  PWR_VCC_42_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_42_FROM
    );
  PWR_VCC_42_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_42_GROM
    );
  PWR_VCC_42_XUSED : X_BUF
    port map (
      I => PWR_VCC_42_FROM,
      O => GLOBAL_LOGIC1_41
    );
  PWR_VCC_42_YUSED : X_BUF
    port map (
      I => PWR_VCC_42_GROM,
      O => GLOBAL_LOGIC0_23
    );
  PWR_VCC_43_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_43_FROM
    );
  PWR_VCC_43_XUSED : X_BUF
    port map (
      I => PWR_VCC_43_FROM,
      O => GLOBAL_LOGIC1_42
    );
  PWR_VCC_44_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_44_FROM
    );
  PWR_VCC_44_XUSED : X_BUF
    port map (
      I => PWR_VCC_44_FROM,
      O => GLOBAL_LOGIC1_43
    );
  PWR_VCC_45_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_45_FROM
    );
  PWR_VCC_45_XUSED : X_BUF
    port map (
      I => PWR_VCC_45_FROM,
      O => GLOBAL_LOGIC1_44
    );
  PWR_VCC_46_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_46_FROM
    );
  PWR_VCC_46_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_46_GROM
    );
  PWR_VCC_46_XUSED : X_BUF
    port map (
      I => PWR_VCC_46_FROM,
      O => GLOBAL_LOGIC1_45
    );
  PWR_VCC_46_YUSED : X_BUF
    port map (
      I => PWR_VCC_46_GROM,
      O => GLOBAL_LOGIC0_16
    );
  PWR_VCC_47_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_47_FROM
    );
  PWR_VCC_47_XUSED : X_BUF
    port map (
      I => PWR_VCC_47_FROM,
      O => GLOBAL_LOGIC1_46
    );
  PWR_GND_0_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_0_GROM
    );
  PWR_GND_0_YUSED : X_BUF
    port map (
      I => PWR_GND_0_GROM,
      O => GLOBAL_LOGIC0
    );
  PWR_GND_1_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_1_GROM
    );
  PWR_GND_1_YUSED : X_BUF
    port map (
      I => PWR_GND_1_GROM,
      O => GLOBAL_LOGIC0_0
    );
  PWR_GND_2_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_2_GROM
    );
  PWR_GND_2_YUSED : X_BUF
    port map (
      I => PWR_GND_2_GROM,
      O => GLOBAL_LOGIC0_1
    );
  PWR_GND_3_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_3_GROM
    );
  PWR_GND_3_YUSED : X_BUF
    port map (
      I => PWR_GND_3_GROM,
      O => GLOBAL_LOGIC0_2
    );
  PWR_GND_4_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_4_GROM
    );
  PWR_GND_4_YUSED : X_BUF
    port map (
      I => PWR_GND_4_GROM,
      O => GLOBAL_LOGIC0_3
    );
  PWR_GND_5_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_5_GROM
    );
  PWR_GND_5_YUSED : X_BUF
    port map (
      I => PWR_GND_5_GROM,
      O => GLOBAL_LOGIC0_4
    );
  PWR_GND_6_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_6_GROM
    );
  PWR_GND_6_YUSED : X_BUF
    port map (
      I => PWR_GND_6_GROM,
      O => GLOBAL_LOGIC0_5
    );
  PWR_GND_7_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_7_GROM
    );
  PWR_GND_7_YUSED : X_BUF
    port map (
      I => PWR_GND_7_GROM,
      O => GLOBAL_LOGIC0_6
    );
  PWR_GND_8_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_8_GROM
    );
  PWR_GND_8_YUSED : X_BUF
    port map (
      I => PWR_GND_8_GROM,
      O => GLOBAL_LOGIC0_7
    );
  PWR_GND_9_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_9_GROM
    );
  PWR_GND_9_YUSED : X_BUF
    port map (
      I => PWR_GND_9_GROM,
      O => GLOBAL_LOGIC0_8
    );
  PWR_GND_10_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_10_GROM
    );
  PWR_GND_10_YUSED : X_BUF
    port map (
      I => PWR_GND_10_GROM,
      O => GLOBAL_LOGIC0_9
    );
  PWR_GND_11_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_11_GROM
    );
  PWR_GND_11_YUSED : X_BUF
    port map (
      I => PWR_GND_11_GROM,
      O => GLOBAL_LOGIC0_10
    );
  PWR_GND_12_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_12_GROM
    );
  PWR_GND_12_YUSED : X_BUF
    port map (
      I => PWR_GND_12_GROM,
      O => GLOBAL_LOGIC0_11
    );
  PWR_GND_13_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_13_GROM
    );
  PWR_GND_13_YUSED : X_BUF
    port map (
      I => PWR_GND_13_GROM,
      O => GLOBAL_LOGIC0_12
    );
  PWR_GND_14_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_14_GROM
    );
  PWR_GND_14_YUSED : X_BUF
    port map (
      I => PWR_GND_14_GROM,
      O => GLOBAL_LOGIC0_13
    );
  PWR_GND_15_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_15_GROM
    );
  PWR_GND_15_YUSED : X_BUF
    port map (
      I => PWR_GND_15_GROM,
      O => GLOBAL_LOGIC0_14
    );
  PWR_GND_16_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_16_GROM
    );
  PWR_GND_16_YUSED : X_BUF
    port map (
      I => PWR_GND_16_GROM,
      O => GLOBAL_LOGIC0_15
    );
  PWR_GND_17_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_17_GROM
    );
  PWR_GND_17_YUSED : X_BUF
    port map (
      I => PWR_GND_17_GROM,
      O => GLOBAL_LOGIC0_17
    );
  PWR_GND_18_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_18_GROM
    );
  PWR_GND_18_YUSED : X_BUF
    port map (
      I => PWR_GND_18_GROM,
      O => GLOBAL_LOGIC0_18
    );
  PWR_GND_19_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_19_GROM
    );
  PWR_GND_19_YUSED : X_BUF
    port map (
      I => PWR_GND_19_GROM,
      O => GLOBAL_LOGIC0_19
    );
  PWR_GND_20_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_20_GROM
    );
  PWR_GND_20_YUSED : X_BUF
    port map (
      I => PWR_GND_20_GROM,
      O => GLOBAL_LOGIC0_20
    );
  PWR_GND_21_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_21_GROM
    );
  PWR_GND_21_YUSED : X_BUF
    port map (
      I => PWR_GND_21_GROM,
      O => GLOBAL_LOGIC0_21
    );
  PWR_GND_22_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_22_GROM
    );
  PWR_GND_22_YUSED : X_BUF
    port map (
      I => PWR_GND_22_GROM,
      O => GLOBAL_LOGIC0_22
    );
  PWR_GND_23_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_23_GROM
    );
  PWR_GND_23_YUSED : X_BUF
    port map (
      I => PWR_GND_23_GROM,
      O => GLOBAL_LOGIC0_24
    );
  PWR_GND_24_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_24_GROM
    );
  PWR_GND_24_YUSED : X_BUF
    port map (
      I => PWR_GND_24_GROM,
      O => GLOBAL_LOGIC0_25
    );
  PWR_GND_25_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_25_GROM
    );
  PWR_GND_25_YUSED : X_BUF
    port map (
      I => PWR_GND_25_GROM,
      O => GLOBAL_LOGIC0_26
    );
  PWR_GND_26_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_26_GROM
    );
  PWR_GND_26_YUSED : X_BUF
    port map (
      I => PWR_GND_26_GROM,
      O => GLOBAL_LOGIC0_27
    );
  PWR_GND_27_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_27_GROM
    );
  PWR_GND_27_YUSED : X_BUF
    port map (
      I => PWR_GND_27_GROM,
      O => GLOBAL_LOGIC0_31
    );
  PWR_GND_28_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_28_GROM
    );
  PWR_GND_28_YUSED : X_BUF
    port map (
      I => PWR_GND_28_GROM,
      O => GLOBAL_LOGIC0_33
    );
  PWR_GND_29_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_29_GROM
    );
  PWR_GND_29_YUSED : X_BUF
    port map (
      I => PWR_GND_29_GROM,
      O => GLOBAL_LOGIC0_35
    );
  PWR_GND_30_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_30_GROM
    );
  PWR_GND_30_YUSED : X_BUF
    port map (
      I => PWR_GND_30_GROM,
      O => GLOBAL_LOGIC0_37
    );
  PWR_GND_31_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_31_GROM
    );
  PWR_GND_31_YUSED : X_BUF
    port map (
      I => PWR_GND_31_GROM,
      O => GLOBAL_LOGIC0_38
    );
  PWR_GND_32_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_32_GROM
    );
  PWR_GND_32_YUSED : X_BUF
    port map (
      I => PWR_GND_32_GROM,
      O => GLOBAL_LOGIC0_42
    );
  PWR_GND_33_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_33_GROM
    );
  PWR_GND_33_YUSED : X_BUF
    port map (
      I => PWR_GND_33_GROM,
      O => GLOBAL_LOGIC0_43
    );
  PWR_GND_34_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_34_GROM
    );
  PWR_GND_34_YUSED : X_BUF
    port map (
      I => PWR_GND_34_GROM,
      O => GLOBAL_LOGIC0_44
    );
  PWR_GND_35_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_35_GROM
    );
  PWR_GND_35_YUSED : X_BUF
    port map (
      I => PWR_GND_35_GROM,
      O => GLOBAL_LOGIC0_46
    );
  PWR_GND_36_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_36_GROM
    );
  PWR_GND_36_YUSED : X_BUF
    port map (
      I => PWR_GND_36_GROM,
      O => GLOBAL_LOGIC0_48
    );
  PWR_GND_37_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_37_GROM
    );
  PWR_GND_37_YUSED : X_BUF
    port map (
      I => PWR_GND_37_GROM,
      O => GLOBAL_LOGIC0_49
    );
  PWR_GND_38_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_38_GROM
    );
  PWR_GND_38_YUSED : X_BUF
    port map (
      I => PWR_GND_38_GROM,
      O => GLOBAL_LOGIC0_52
    );
  PWR_GND_39_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_39_GROM
    );
  PWR_GND_39_YUSED : X_BUF
    port map (
      I => PWR_GND_39_GROM,
      O => GLOBAL_LOGIC0_53
    );
  PWR_GND_40_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_40_GROM
    );
  PWR_GND_40_YUSED : X_BUF
    port map (
      I => PWR_GND_40_GROM,
      O => GLOBAL_LOGIC0_54
    );
  PWR_GND_41_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_41_GROM
    );
  PWR_GND_41_YUSED : X_BUF
    port map (
      I => PWR_GND_41_GROM,
      O => GLOBAL_LOGIC0_55
    );
  PWR_GND_42_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_42_GROM
    );
  PWR_GND_42_YUSED : X_BUF
    port map (
      I => PWR_GND_42_GROM,
      O => GLOBAL_LOGIC0_56
    );
  PWR_GND_43_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_43_GROM
    );
  PWR_GND_43_YUSED : X_BUF
    port map (
      I => PWR_GND_43_GROM,
      O => GLOBAL_LOGIC0_59
    );
  PWR_GND_44_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_44_GROM
    );
  PWR_GND_44_YUSED : X_BUF
    port map (
      I => PWR_GND_44_GROM,
      O => GLOBAL_LOGIC0_60
    );
  PWR_GND_45_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_45_GROM
    );
  PWR_GND_45_YUSED : X_BUF
    port map (
      I => PWR_GND_45_GROM,
      O => GLOBAL_LOGIC0_61
    );
  PWR_GND_46_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_46_GROM
    );
  PWR_GND_46_YUSED : X_BUF
    port map (
      I => PWR_GND_46_GROM,
      O => GLOBAL_LOGIC0_62
    );
  PWR_GND_47_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_47_GROM
    );
  PWR_GND_47_YUSED : X_BUF
    port map (
      I => PWR_GND_47_GROM,
      O => GLOBAL_LOGIC0_63
    );
  PWR_GND_48_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_48_GROM
    );
  PWR_GND_48_YUSED : X_BUF
    port map (
      I => PWR_GND_48_GROM,
      O => GLOBAL_LOGIC0_64
    );
  PWR_GND_49_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_49_GROM
    );
  PWR_GND_49_YUSED : X_BUF
    port map (
      I => PWR_GND_49_GROM,
      O => GLOBAL_LOGIC0_65
    );
  PWR_GND_50_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_50_GROM
    );
  PWR_GND_50_YUSED : X_BUF
    port map (
      I => PWR_GND_50_GROM,
      O => GLOBAL_LOGIC0_66
    );
  PWR_GND_51_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_51_GROM
    );
  PWR_GND_51_YUSED : X_BUF
    port map (
      I => PWR_GND_51_GROM,
      O => GLOBAL_LOGIC0_68
    );
  PWR_GND_52_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_52_GROM
    );
  PWR_GND_52_YUSED : X_BUF
    port map (
      I => PWR_GND_52_GROM,
      O => GLOBAL_LOGIC0_69
    );
  PWR_GND_53_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_53_GROM
    );
  PWR_GND_53_YUSED : X_BUF
    port map (
      I => PWR_GND_53_GROM,
      O => GLOBAL_LOGIC0_70
    );
  NlwBlock_testsuite_GND : X_ZERO
    port map (
      O => GND
    );
  NlwBlock_testsuite_VCC : X_ONE
    port map (
      O => VCC
    );
  NlwBlockROC : X_ROC
    generic map (ROC_WIDTH => 100 ns)
    port map (O => GSR);
  NlwBlockTOC : X_TOC
    port map (O => GTS);

end Structure;

