-- Xilinx Vhdl netlist produced by netgen application (version G.24)
-- Command       : -intstyle ise -s 6 -pcf network.pcf -ngm network.ngm -rpw 100 -tpw 0 -ar Structure -xon false -w -ofmt vhdl -sim network.ncd network_PR.vhd 
-- Input file    : network.ncd
-- Output file   : network_PR.vhd
-- Design name   : network
-- # of Entities : 1
-- Xilinx        : C:/Xilinx
-- Device        : 2s300epq208-6 (PRODUCTION 1.17 2003-06-19)

-- This vhdl netlist is a simulation model and uses simulation 
-- primitives which may not represent the true implementation of the 
-- device, however the netlist is functionally correct and should not 
-- be modified. This file cannot be synthesized and should only be used 
-- with supported simulation tools.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library SIMPRIM;
use SIMPRIM.VCOMPONENTS.ALL;
use SIMPRIM.VPACKAGE.ALL;

entity network is
  port (
    DOUTEN : out STD_LOGIC; 
    MCLK : out STD_LOGIC; 
    LED100 : out STD_LOGIC; 
    LED1000 : out STD_LOGIC; 
    PHYRESET : out STD_LOGIC; 
    GTX_CLK : out STD_LOGIC; 
    LEDACT : out STD_LOGIC; 
    SOUT : out STD_LOGIC; 
    MWE : out STD_LOGIC; 
    TX_EN : out STD_LOGIC; 
    LEDDPX : out STD_LOGIC; 
    LEDTX : out STD_LOGIC; 
    LEDRX : out STD_LOGIC; 
    MDC : out STD_LOGIC; 
    MDIO : inout STD_LOGIC; 
    SCS : in STD_LOGIC := 'X'; 
    NEXTFRAME : in STD_LOGIC := 'X'; 
    SCLK : in STD_LOGIC := 'X'; 
    DINEN : in STD_LOGIC := 'X'; 
    CLKIOIN : in STD_LOGIC := 'X'; 
    RX_CLK : in STD_LOGIC := 'X'; 
    NEWFRAME : in STD_LOGIC := 'X'; 
    RESET : in STD_LOGIC := 'X'; 
    CLKIN : in STD_LOGIC := 'X'; 
    RX_ER : in STD_LOGIC := 'X'; 
    RX_DV : in STD_LOGIC := 'X'; 
    SIN : in STD_LOGIC := 'X'; 
    DOUT : out STD_LOGIC_VECTOR ( 15 downto 0 ); 
    TXD : out STD_LOGIC_VECTOR ( 7 downto 0 ); 
    MA : out STD_LOGIC_VECTOR ( 16 downto 0 ); 
    MD : inout STD_LOGIC_VECTOR ( 31 downto 0 ); 
    RXD : in STD_LOGIC_VECTOR ( 7 downto 0 ); 
    DIN : in STD_LOGIC_VECTOR ( 15 downto 0 ) 
  );
end network;

architecture Structure of network is
  signal rx_input_fifo_fifo_N1552 : STD_LOGIC; 
  signal clkrx : STD_LOGIC; 
  signal rx_input_fifo_RESET_1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1559 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1524 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1497 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1573 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1495 : STD_LOGIC; 
  signal GTX_CLK_OBUF : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1538 : STD_LOGIC; 
  signal rx_input_ince : STD_LOGIC; 
  signal rx_input_fifo_fifo_full : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3373 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3366 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1580 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1545 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2718 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1539 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3368 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1582 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1540 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1547 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1581 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1546 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4321 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2708 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1525 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1526 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1541 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3370 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1584 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1542 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1549 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1583 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1548 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1553 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1554 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1574 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1575 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4313 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1561 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1560 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2698 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1527 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1528 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1586 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1544 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1551 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1585 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1543 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1550 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1555 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1556 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1576 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1577 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4305 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1563 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1562 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3676 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1529 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1530 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1557 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1558 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1578 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1579 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1565 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1564 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N17 : STD_LOGIC; 
  signal rx_input_rx_nearf : STD_LOGIC; 
  signal rx_input_fifo_rd_en : STD_LOGIC; 
  signal rx_input_fifo_fifo_empty : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2449 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2442 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1594 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1891 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2444 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1596 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1595 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1881 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2446 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1598 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1597 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1871 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1600 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1599 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N16 : STD_LOGIC; 
  signal mac_control_n0024 : STD_LOGIC; 
  signal mac_control_CLKSL_4 : STD_LOGIC; 
  signal rx_input_memio_N80955 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_1 : STD_LOGIC; 
  signal rx_input_memio_RESET_1 : STD_LOGIC; 
  signal rx_input_memio_crcrst : STD_LOGIC; 
  signal mac_control_sclkl : STD_LOGIC; 
  signal RESET_IBUF : STD_LOGIC; 
  signal mac_control_CLKSL_1 : STD_LOGIC; 
  signal mac_control_sclkll : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE1101 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N70497 : STD_LOGIC; 
  signal rx_input_memio_n0044 : STD_LOGIC; 
  signal RESET_IBUF_2 : STD_LOGIC; 
  signal rx_input_memio_n0045 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N38617 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE951 : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd2 : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd1 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1623 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1588 : STD_LOGIC; 
  signal rx_output_cs_FFd7 : STD_LOGIC; 
  signal rx_output_nf : STD_LOGIC; 
  signal rx_output_fifo_full : STD_LOGIC; 
  signal rx_output_cs_FFd5 : STD_LOGIC; 
  signal rx_output_CHOICE1106 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1602 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1581 : STD_LOGIC; 
  signal rx_input_fifo_control_n0008 : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4 : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd3 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1591 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1630 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1644 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1584 : STD_LOGIC; 
  signal tx_output_bcnt_42 : STD_LOGIC; 
  signal tx_output_bcnt_43 : STD_LOGIC; 
  signal tx_output_bcnt_44 : STD_LOGIC; 
  signal tx_output_bcnt_45 : STD_LOGIC; 
  signal tx_output_CHOICE1871 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1595 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1637 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1647 : STD_LOGIC; 
  signal tx_output_n0033 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_219 : STD_LOGIC; 
  signal tx_output_cs_FFd12 : STD_LOGIC; 
  signal tx_output_bcnt_53 : STD_LOGIC; 
  signal tx_output_bcnt_50 : STD_LOGIC; 
  signal tx_output_bcnt_51 : STD_LOGIC; 
  signal tx_output_bcnt_52 : STD_LOGIC; 
  signal tx_output_CHOICE1886 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1640 : STD_LOGIC; 
  signal tx_output_bcnt_46 : STD_LOGIC; 
  signal tx_output_bcnt_47 : STD_LOGIC; 
  signal tx_output_bcnt_48 : STD_LOGIC; 
  signal tx_output_bcnt_49 : STD_LOGIC; 
  signal tx_output_CHOICE1879 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1609 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1616 : STD_LOGIC; 
  signal tx_output_cs_FFd4_In : STD_LOGIC; 
  signal tx_output_N80951 : STD_LOGIC; 
  signal tx_output_cs_FFd5_1 : STD_LOGIC; 
  signal tx_output_n0007 : STD_LOGIC; 
  signal tx_output_cs_FFd4 : STD_LOGIC; 
  signal tx_output_cs_FFd4_1 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1633 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1619 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1626 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1612 : STD_LOGIC; 
  signal rx_input_ce : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1605 : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1598 : STD_LOGIC; 
  signal rx_output_cs_FFd1 : STD_LOGIC; 
  signal rx_output_cs_FFd11 : STD_LOGIC; 
  signal rx_output_N34486 : STD_LOGIC; 
  signal rx_output_n0018 : STD_LOGIC; 
  signal rx_output_cs_FFd9 : STD_LOGIC; 
  signal tx_output_n0025 : STD_LOGIC; 
  signal tx_output_cs_FFd16_1 : STD_LOGIC; 
  signal tx_output_crc_6_Q : STD_LOGIC; 
  signal mac_control_N69572 : STD_LOGIC; 
  signal mac_control_sclkdeltal : STD_LOGIC; 
  signal mac_control_addr_0_1 : STD_LOGIC; 
  signal mac_control_N53109 : STD_LOGIC; 
  signal mac_control_n0028 : STD_LOGIC; 
  signal mac_control_N69759 : STD_LOGIC; 
  signal mac_control_N53132 : STD_LOGIC; 
  signal mac_control_N53144 : STD_LOGIC; 
  signal mac_control_n0033 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0004 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd3 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd2 : STD_LOGIC; 
  signal tx_output_crc_7_Q : STD_LOGIC; 
  signal tx_input_N80947 : STD_LOGIC; 
  signal tx_input_CHOICE1988 : STD_LOGIC; 
  signal tx_input_CHOICE2014 : STD_LOGIC; 
  signal tx_input_CHOICE1991 : STD_LOGIC; 
  signal mac_control_n0012 : STD_LOGIC; 
  signal clksl : STD_LOGIC; 
  signal mac_control_n0060 : STD_LOGIC; 
  signal mac_control_CHOICE2625 : STD_LOGIC; 
  signal mac_control_n0086 : STD_LOGIC; 
  signal mac_control_sclkdeltall : STD_LOGIC; 
  signal mac_control_N81427 : STD_LOGIC; 
  signal mac_control_PHY_status_n0011 : STD_LOGIC; 
  signal mac_control_CLKSL_3 : STD_LOGIC; 
  signal mac_control_CLKSL_2 : STD_LOGIC; 
  signal mac_control_CHOICE2651 : STD_LOGIC; 
  signal mac_control_N81431 : STD_LOGIC; 
  signal txfifofull : STD_LOGIC; 
  signal RESET_IBUF_1 : STD_LOGIC; 
  signal tx_input_fifofulll : STD_LOGIC; 
  signal mac_control_CHOICE2449 : STD_LOGIC; 
  signal mac_control_N81435 : STD_LOGIC; 
  signal tx_output_crc_8_Q : STD_LOGIC; 
  signal mac_control_CLKSL_5 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1839 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1846 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1832 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1808 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1812 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1822 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1848 : STD_LOGIC; 
  signal rx_input_memio_crcequal : STD_LOGIC; 
  signal rx_input_memio_menl : STD_LOGIC; 
  signal rx_input_memio_men : STD_LOGIC; 
  signal rx_input_RESET_1 : STD_LOGIC; 
  signal rx_input_memio_n0033 : STD_LOGIC; 
  signal rx_input_memio_n00331_1 : STD_LOGIC; 
  signal mac_control_CHOICE2424 : STD_LOGIC; 
  signal mac_control_N81439 : STD_LOGIC; 
  signal rx_output_fifo_nearfull : STD_LOGIC; 
  signal tx_output_crc_9_Q : STD_LOGIC; 
  signal mac_control_CHOICE2677 : STD_LOGIC; 
  signal mac_control_N81443 : STD_LOGIC; 
  signal tx_input_addr_17 : STD_LOGIC; 
  signal tx_input_addr_16 : STD_LOGIC; 
  signal tx_input_mrw : STD_LOGIC; 
  signal tx_input_addr_19 : STD_LOGIC; 
  signal tx_input_addr_18 : STD_LOGIC; 
  signal tx_input_addr_21 : STD_LOGIC; 
  signal tx_input_addr_20 : STD_LOGIC; 
  signal tx_input_addr_23 : STD_LOGIC; 
  signal tx_input_addr_22 : STD_LOGIC; 
  signal tx_input_addr_25 : STD_LOGIC; 
  signal tx_input_addr_24 : STD_LOGIC; 
  signal rx_output_cs_FFd13 : STD_LOGIC; 
  signal rx_output_cs_FFd12 : STD_LOGIC; 
  signal rx_output_cs_FFd15 : STD_LOGIC; 
  signal rx_output_cs_FFd14 : STD_LOGIC; 
  signal rx_output_cs_FFd17 : STD_LOGIC; 
  signal rx_output_cs_FFd16 : STD_LOGIC; 
  signal rx_output_cs_FFd8 : STD_LOGIC; 
  signal rx_output_ceinl : STD_LOGIC; 
  signal rx_output_n0033 : STD_LOGIC; 
  signal rx_output_cs_FFd19 : STD_LOGIC; 
  signal rx_output_cs_FFd10 : STD_LOGIC; 
  signal rx_output_fifo_reset : STD_LOGIC; 
  signal rx_output_n0034 : STD_LOGIC; 
  signal mac_control_CHOICE2703 : STD_LOGIC; 
  signal mac_control_N81447 : STD_LOGIC; 
  signal rxf : STD_LOGIC; 
  signal mac_control_rxf_cross : STD_LOGIC; 
  signal tx_input_cs_FFd2 : STD_LOGIC; 
  signal tx_input_den : STD_LOGIC; 
  signal tx_input_cs_FFd6 : STD_LOGIC; 
  signal tx_input_cs_FFd7 : STD_LOGIC; 
  signal tx_input_n0023 : STD_LOGIC; 
  signal tx_input_n0021 : STD_LOGIC; 
  signal mac_control_CHOICE2474 : STD_LOGIC; 
  signal mac_control_N81451 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_156 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_158 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159 : STD_LOGIC; 
  signal mac_control_CHOICE1266 : STD_LOGIC; 
  signal mac_control_CHOICE1269 : STD_LOGIC; 
  signal mac_control_CHOICE1272 : STD_LOGIC; 
  signal mac_control_n0040 : STD_LOGIC; 
  signal mac_control_phyrstcnt_128 : STD_LOGIC; 
  signal mac_control_phyrstcnt_129 : STD_LOGIC; 
  signal mac_control_phyrstcnt_111 : STD_LOGIC; 
  signal mac_control_phyrstcnt_130 : STD_LOGIC; 
  signal mac_control_CHOICE1384 : STD_LOGIC; 
  signal mac_control_CHOICE1387 : STD_LOGIC; 
  signal mac_control_CHOICE1388 : STD_LOGIC; 
  signal mac_control_phyrstcnt_117 : STD_LOGIC; 
  signal mac_control_phyrstcnt_118 : STD_LOGIC; 
  signal mac_control_phyrstcnt_125 : STD_LOGIC; 
  signal mac_control_phyrstcnt_126 : STD_LOGIC; 
  signal mac_control_phyrstcnt_124 : STD_LOGIC; 
  signal mac_control_phyrstcnt_127 : STD_LOGIC; 
  signal mac_control_N80971 : STD_LOGIC; 
  signal mac_control_phyrstcnt_138 : STD_LOGIC; 
  signal mac_control_phyrstcnt_139 : STD_LOGIC; 
  signal mac_control_phyrstcnt_112 : STD_LOGIC; 
  signal mac_control_phyrstcnt_140 : STD_LOGIC; 
  signal mac_control_phyrstcnt_135 : STD_LOGIC; 
  signal mac_control_phyrstcnt_136 : STD_LOGIC; 
  signal mac_control_phyrstcnt_137 : STD_LOGIC; 
  signal mac_control_CHOICE1333 : STD_LOGIC; 
  signal mac_control_CHOICE1395 : STD_LOGIC; 
  signal mac_control_phyrstcnt_134 : STD_LOGIC; 
  signal mac_control_CHOICE1325 : STD_LOGIC; 
  signal mac_control_phyrstcnt_120 : STD_LOGIC; 
  signal mac_control_phyrstcnt_132 : STD_LOGIC; 
  signal mac_control_phyrstcnt_133 : STD_LOGIC; 
  signal mac_control_CHOICE1326 : STD_LOGIC; 
  signal mac_control_phyrstcnt_113 : STD_LOGIC; 
  signal mac_control_CHOICE1399 : STD_LOGIC; 
  signal mac_control_phyrstcnt_114 : STD_LOGIC; 
  signal mac_control_phyrstcnt_115 : STD_LOGIC; 
  signal mac_control_phyrstcnt_116 : STD_LOGIC; 
  signal mac_control_CHOICE1402 : STD_LOGIC; 
  signal mac_control_CHOICE1340 : STD_LOGIC; 
  signal mac_control_CHOICE1341 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0011 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_152 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_153 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_142 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143 : STD_LOGIC; 
  signal mac_control_CHOICE1280 : STD_LOGIC; 
  signal mac_control_CHOICE1308 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_144 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_146 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147 : STD_LOGIC; 
  signal mac_control_CHOICE1277 : STD_LOGIC; 
  signal mac_control_CHOICE1283 : STD_LOGIC; 
  signal mac_control_n0038 : STD_LOGIC; 
  signal mac_control_ledtx_rst : STD_LOGIC; 
  signal mac_control_CHOICE1302 : STD_LOGIC; 
  signal mac_control_CHOICE1305 : STD_LOGIC; 
  signal mac_control_CHOICE1311 : STD_LOGIC; 
  signal mac_control_n0037 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_164 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_165 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_154 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155 : STD_LOGIC; 
  signal mac_control_CHOICE1294 : STD_LOGIC; 
  signal mac_control_ledrx_rst : STD_LOGIC; 
  signal mac_control_CHOICE1288 : STD_LOGIC; 
  signal mac_control_CHOICE1291 : STD_LOGIC; 
  signal mac_control_CHOICE1297 : STD_LOGIC; 
  signal mac_control_n0039 : STD_LOGIC; 
  signal mac_control_CHOICE2729 : STD_LOGIC; 
  signal mac_control_N81455 : STD_LOGIC; 
  signal rx_input_memio_crccomb_N81261 : STD_LOGIC; 
  signal tx_input_n0020 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_37 : STD_LOGIC; 
  signal MDC_OBUF : STD_LOGIC; 
  signal mac_control_CHOICE2524 : STD_LOGIC; 
  signal mac_control_N81459 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_1_68 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_0_69 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_3_66 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_2_67 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_5_64 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_4_65 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_7_62 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_6_63 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_9_60 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_8_61 : STD_LOGIC; 
  signal memcontroller_n00061_1 : STD_LOGIC; 
  signal memcontroller_n00051_1 : STD_LOGIC; 
  signal mac_control_n0064 : STD_LOGIC; 
  signal mac_control_n0065 : STD_LOGIC; 
  signal mac_control_CHOICE2634 : STD_LOGIC; 
  signal mac_control_CHOICE2738 : STD_LOGIC; 
  signal mac_control_n0067 : STD_LOGIC; 
  signal mac_control_n0062 : STD_LOGIC; 
  signal mac_control_CHOICE2508 : STD_LOGIC; 
  signal mac_control_CHOICE2483 : STD_LOGIC; 
  signal mac_control_CHOICE2105 : STD_LOGIC; 
  signal mac_control_CHOICE2128 : STD_LOGIC; 
  signal mac_control_CHOICE2243 : STD_LOGIC; 
  signal mac_control_CHOICE2533 : STD_LOGIC; 
  signal mac_control_CHOICE2583 : STD_LOGIC; 
  signal mac_control_CHOICE2558 : STD_LOGIC; 
  signal mac_control_CHOICE2712 : STD_LOGIC; 
  signal mac_control_CHOICE2360 : STD_LOGIC; 
  signal mac_control_CHOICE2174 : STD_LOGIC; 
  signal mac_control_CHOICE2289 : STD_LOGIC; 
  signal mac_control_CHOICE2384 : STD_LOGIC; 
  signal mac_control_CHOICE2764 : STD_LOGIC; 
  signal mac_control_n0066 : STD_LOGIC; 
  signal mac_control_n0059 : STD_LOGIC; 
  signal mac_control_CHOICE2387 : STD_LOGIC; 
  signal mac_control_CHOICE1895 : STD_LOGIC; 
  signal mac_control_CHOICE2082 : STD_LOGIC; 
  signal mac_control_CHOICE2151 : STD_LOGIC; 
  signal mac_control_n00851_1 : STD_LOGIC; 
  signal mac_control_n0063 : STD_LOGIC; 
  signal mac_control_CHOICE2698 : STD_LOGIC; 
  signal mac_control_CHOICE1904 : STD_LOGIC; 
  signal mac_control_n0061 : STD_LOGIC; 
  signal mac_control_n0056 : STD_LOGIC; 
  signal mac_control_CHOICE1899 : STD_LOGIC; 
  signal mac_control_N81050 : STD_LOGIC; 
  signal mac_control_CHOICE2660 : STD_LOGIC; 
  signal mac_control_CHOICE2312 : STD_LOGIC; 
  signal mac_control_CHOICE2637 : STD_LOGIC; 
  signal mac_control_CHOICE2611 : STD_LOGIC; 
  signal mac_control_CHOICE2043 : STD_LOGIC; 
  signal mac_control_CHOICE2336 : STD_LOGIC; 
  signal mac_control_CHOICE2408 : STD_LOGIC; 
  signal mac_control_CHOICE2197 : STD_LOGIC; 
  signal mac_control_CHOICE2615 : STD_LOGIC; 
  signal mac_control_N81034 : STD_LOGIC; 
  signal mac_control_CHOICE1892 : STD_LOGIC; 
  signal mac_control_CHOICE1907 : STD_LOGIC; 
  signal mac_control_N81030 : STD_LOGIC; 
  signal mac_control_n0044 : STD_LOGIC; 
  signal mac_control_CHOICE2220 : STD_LOGIC; 
  signal mac_control_CHOICE2059 : STD_LOGIC; 
  signal mac_control_CHOICE2641 : STD_LOGIC; 
  signal mac_control_N81062 : STD_LOGIC; 
  signal mac_control_CHOICE2372 : STD_LOGIC; 
  signal mac_control_CHOICE2646 : STD_LOGIC; 
  signal mac_control_CHOICE2608 : STD_LOGIC; 
  signal mac_control_CHOICE2620 : STD_LOGIC; 
  signal mac_control_CHOICE2623 : STD_LOGIC; 
  signal mac_control_n0057 : STD_LOGIC; 
  signal mac_control_CHOICE2108 : STD_LOGIC; 
  signal mac_control_CHOICE2436 : STD_LOGIC; 
  signal mac_control_CHOICE2433 : STD_LOGIC; 
  signal mac_control_CHOICE2266 : STD_LOGIC; 
  signal mac_control_CHOICE2296 : STD_LOGIC; 
  signal mac_control_CHOICE2440 : STD_LOGIC; 
  signal mac_control_CHOICE2649 : STD_LOGIC; 
  signal mac_control_CHOICE2246 : STD_LOGIC; 
  signal mac_control_CHOICE2411 : STD_LOGIC; 
  signal mac_control_CHOICE2444 : STD_LOGIC; 
  signal mac_control_N81106 : STD_LOGIC; 
  signal mac_control_CHOICE2447 : STD_LOGIC; 
  signal mac_control_CHOICE2715 : STD_LOGIC; 
  signal mac_control_CHOICE2663 : STD_LOGIC; 
  signal mac_control_CHOICE2419 : STD_LOGIC; 
  signal mac_control_N81122 : STD_LOGIC; 
  signal mac_control_CHOICE2415 : STD_LOGIC; 
  signal mac_control_CHOICE2422 : STD_LOGIC; 
  signal mac_control_CHOICE2667 : STD_LOGIC; 
  signal mac_control_N81054 : STD_LOGIC; 
  signal mac_control_CHOICE2324 : STD_LOGIC; 
  signal mac_control_CHOICE2672 : STD_LOGIC; 
  signal mac_control_CHOICE2741 : STD_LOGIC; 
  signal mac_control_CHOICE2689 : STD_LOGIC; 
  signal mac_control_CHOICE2693 : STD_LOGIC; 
  signal mac_control_N81078 : STD_LOGIC; 
  signal mac_control_CHOICE2675 : STD_LOGIC; 
  signal mac_control_CHOICE2292 : STD_LOGIC; 
  signal mac_control_CHOICE2461 : STD_LOGIC; 
  signal mac_control_CHOICE2250 : STD_LOGIC; 
  signal mac_control_CHOICE2465 : STD_LOGIC; 
  signal mac_control_CHOICE2686 : STD_LOGIC; 
  signal mac_control_CHOICE2701 : STD_LOGIC; 
  signal tx_output_crc_loigc_N81257 : STD_LOGIC; 
  signal tx_output_CHOICE1439 : STD_LOGIC; 
  signal mac_control_CHOICE2469 : STD_LOGIC; 
  signal mac_control_N81150 : STD_LOGIC; 
  signal mac_control_CHOICE2458 : STD_LOGIC; 
  signal mac_control_CHOICE2472 : STD_LOGIC; 
  signal mac_control_CHOICE2719 : STD_LOGIC; 
  signal mac_control_N81066 : STD_LOGIC; 
  signal mac_control_CHOICE2396 : STD_LOGIC; 
  signal mac_control_CHOICE2724 : STD_LOGIC; 
  signal mac_control_CHOICE2177 : STD_LOGIC; 
  signal mac_control_CHOICE2511 : STD_LOGIC; 
  signal mac_control_CHOICE2540 : STD_LOGIC; 
  signal mac_control_CHOICE2515 : STD_LOGIC; 
  signal mac_control_CHOICE2727 : STD_LOGIC; 
  signal mac_control_CHOICE2519 : STD_LOGIC; 
  signal mac_control_N81114 : STD_LOGIC; 
  signal mac_control_CHOICE2522 : STD_LOGIC; 
  signal rx_output_cs_FFd6 : STD_LOGIC; 
  signal rx_output_cs_FFd3 : STD_LOGIC; 
  signal rx_output_cs_FFd2 : STD_LOGIC; 
  signal rx_output_CHOICE1800 : STD_LOGIC; 
  signal rx_output_CHOICE876 : STD_LOGIC; 
  signal clkio : STD_LOGIC; 
  signal rx_output_cs_FFd4 : STD_LOGIC; 
  signal rx_output_CHOICE879 : STD_LOGIC; 
  signal rx_output_denl : STD_LOGIC; 
  signal mac_control_lrxbcast : STD_LOGIC; 
  signal rxbcast : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81159 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE886 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE901 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE892 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE902 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE900 : STD_LOGIC; 
  signal tx_input_cs_FFd4 : STD_LOGIC; 
  signal tx_input_cs_FFd11 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1525 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1535 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1542 : STD_LOGIC; 
  signal tx_output_CHOICE1505 : STD_LOGIC; 
  signal tx_output_CHOICE1516 : STD_LOGIC; 
  signal tx_output_CHOICE1521 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0015 : STD_LOGIC; 
  signal tx_output_CHOICE1483 : STD_LOGIC; 
  signal tx_output_CHOICE1494 : STD_LOGIC; 
  signal tx_output_CHOICE1499 : STD_LOGIC; 
  signal tx_output_CHOICE1510 : STD_LOGIC; 
  signal tx_output_CHOICE1488 : STD_LOGIC; 
  signal tx_output_CHOICE1450 : STD_LOGIC; 
  signal tx_output_CHOICE1461 : STD_LOGIC; 
  signal tx_output_CHOICE1466 : STD_LOGIC; 
  signal tx_output_CHOICE1472 : STD_LOGIC; 
  signal tx_output_CHOICE1477 : STD_LOGIC; 
  signal tx_output_CHOICE1455 : STD_LOGIC; 
  signal tx_output_CHOICE1444 : STD_LOGIC; 
  signal mac_control_lrxmcast : STD_LOGIC; 
  signal rxmcast : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1950 : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1957 : STD_LOGIC; 
  signal mac_control_CHOICE2755 : STD_LOGIC; 
  signal mac_control_N81463 : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1972 : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1965 : STD_LOGIC; 
  signal rx_fifocheck_n0003 : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1973 : STD_LOGIC; 
  signal rx_fifocheck_n0002 : STD_LOGIC; 
  signal mac_control_lrxucast : STD_LOGIC; 
  signal rxucast : STD_LOGIC; 
  signal mac_control_CHOICE2139 : STD_LOGIC; 
  signal mac_control_CHOICE2131 : STD_LOGIC; 
  signal mac_control_CHOICE2135 : STD_LOGIC; 
  signal mac_control_N81102 : STD_LOGIC; 
  signal mac_control_CHOICE2142 : STD_LOGIC; 
  signal mac_control_CHOICE2499 : STD_LOGIC; 
  signal mac_control_N81467 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd1 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0032 : STD_LOGIC; 
  signal tx_output_cs_FFd16 : STD_LOGIC; 
  signal tx_output_crc_12_Q : STD_LOGIC; 
  signal tx_output_crcenl : STD_LOGIC; 
  signal tx_output_cs_FFd10 : STD_LOGIC; 
  signal tx_output_cs_FFd9 : STD_LOGIC; 
  signal tx_output_cs_FFd8 : STD_LOGIC; 
  signal tx_output_cs_FFd6_1 : STD_LOGIC; 
  signal tx_output_cs_FFd11 : STD_LOGIC; 
  signal tx_output_cs_FFd13 : STD_LOGIC; 
  signal tx_output_CHOICE1775 : STD_LOGIC; 
  signal tx_output_CHOICE1760 : STD_LOGIC; 
  signal tx_output_cs_FFd7 : STD_LOGIC; 
  signal tx_output_cs_FFd3 : STD_LOGIC; 
  signal tx_output_CHOICE1682 : STD_LOGIC; 
  signal tx_output_CHOICE1779 : STD_LOGIC; 
  signal tx_output_cs_FFd2 : STD_LOGIC; 
  signal tx_output_cs_FFd1 : STD_LOGIC; 
  signal tx_output_cs_FFd15 : STD_LOGIC; 
  signal tx_output_CHOICE1782 : STD_LOGIC; 
  signal mac_control_CHOICE2549 : STD_LOGIC; 
  signal mac_control_N81471 : STD_LOGIC; 
  signal mac_control_CHOICE2367 : STD_LOGIC; 
  signal mac_control_CHOICE2363 : STD_LOGIC; 
  signal mac_control_N81038 : STD_LOGIC; 
  signal mac_control_CHOICE2375 : STD_LOGIC; 
  signal mac_control_PHY_status_rwl : STD_LOGIC; 
  signal tx_output_crc_0_Q : STD_LOGIC; 
  signal tx_output_crc_2_Q : STD_LOGIC; 
  signal mac_control_CHOICE2116 : STD_LOGIC; 
  signal mac_control_CHOICE2112 : STD_LOGIC; 
  signal mac_control_N81090 : STD_LOGIC; 
  signal mac_control_CHOICE2119 : STD_LOGIC; 
  signal mac_control_CHOICE2300 : STD_LOGIC; 
  signal mac_control_N81094 : STD_LOGIC; 
  signal mac_control_CHOICE2303 : STD_LOGIC; 
  signal mac_control_CHOICE2574 : STD_LOGIC; 
  signal mac_control_N81475 : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_net187 : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_103 : STD_LOGIC; 
  signal rx_input_GMII_rx_of : STD_LOGIC; 
  signal mac_control_CHOICE2185 : STD_LOGIC; 
  signal mac_control_N80963 : STD_LOGIC; 
  signal mac_control_CHOICE2162 : STD_LOGIC; 
  signal mac_control_CHOICE2154 : STD_LOGIC; 
  signal mac_control_CHOICE2158 : STD_LOGIC; 
  signal mac_control_N81134 : STD_LOGIC; 
  signal mac_control_CHOICE2165 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1817 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1821 : STD_LOGIC; 
  signal mac_control_CHOICE2781 : STD_LOGIC; 
  signal mac_control_N81479 : STD_LOGIC; 
  signal mac_control_CHOICE2599 : STD_LOGIC; 
  signal mac_control_N81483 : STD_LOGIC; 
  signal tx_output_CHOICE1670 : STD_LOGIC; 
  signal tx_output_N81401 : STD_LOGIC; 
  signal mac_control_CHOICE2391 : STD_LOGIC; 
  signal mac_control_N81046 : STD_LOGIC; 
  signal mac_control_CHOICE2399 : STD_LOGIC; 
  signal mac_control_CHOICE2319 : STD_LOGIC; 
  signal mac_control_CHOICE2315 : STD_LOGIC; 
  signal mac_control_N81074 : STD_LOGIC; 
  signal mac_control_CHOICE2327 : STD_LOGIC; 
  signal mac_control_sclkdelta : STD_LOGIC; 
  signal mac_control_N53154 : STD_LOGIC; 
  signal mac_control_n0015 : STD_LOGIC; 
  signal mac_control_n0010 : STD_LOGIC; 
  signal tx_output_ltxen2 : STD_LOGIC; 
  signal tx_output_cs_FFd14 : STD_LOGIC; 
  signal tx_output_N80959 : STD_LOGIC; 
  signal tx_output_ltxen3 : STD_LOGIC; 
  signal mac_control_n0013 : STD_LOGIC; 
  signal mac_control_n0025 : STD_LOGIC; 
  signal mac_control_n0030 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_160 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_162 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163 : STD_LOGIC; 
  signal mac_control_n0029 : STD_LOGIC; 
  signal mac_control_n0026 : STD_LOGIC; 
  signal mac_control_phyrstcnt_121 : STD_LOGIC; 
  signal mac_control_phyrstcnt_122 : STD_LOGIC; 
  signal mac_control_phyrstcnt_123 : STD_LOGIC; 
  signal mac_control_phyrstcnt_119 : STD_LOGIC; 
  signal mac_control_phyrstcnt_110 : STD_LOGIC; 
  signal mac_control_CHOICE1380 : STD_LOGIC; 
  signal mac_control_CHOICE1381 : STD_LOGIC; 
  signal mac_control_N53204 : STD_LOGIC; 
  signal mac_control_n0027 : STD_LOGIC; 
  signal mac_control_n0036 : STD_LOGIC; 
  signal mac_control_n0035 : STD_LOGIC; 
  signal mac_control_CHOICE2208 : STD_LOGIC; 
  signal mac_control_CHOICE2200 : STD_LOGIC; 
  signal mac_control_CHOICE2204 : STD_LOGIC; 
  signal mac_control_N81098 : STD_LOGIC; 
  signal mac_control_CHOICE2211 : STD_LOGIC; 
  signal tx_input_DONE : STD_LOGIC; 
  signal mac_control_N53125 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_148 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_150 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151 : STD_LOGIC; 
  signal mac_control_N81417 : STD_LOGIC; 
  signal mac_control_N53118 : STD_LOGIC; 
  signal mac_control_CHOICE2536 : STD_LOGIC; 
  signal mac_control_CHOICE2343 : STD_LOGIC; 
  signal mac_control_CHOICE2339 : STD_LOGIC; 
  signal mac_control_CHOICE2348 : STD_LOGIC; 
  signal mac_control_N81070 : STD_LOGIC; 
  signal mac_control_CHOICE2351 : STD_LOGIC; 
  signal mac_control_CHOICE2181 : STD_LOGIC; 
  signal mac_control_N81154 : STD_LOGIC; 
  signal mac_control_CHOICE2188 : STD_LOGIC; 
  signal mac_control_CHOICE2070 : STD_LOGIC; 
  signal mac_control_CHOICE2062 : STD_LOGIC; 
  signal mac_control_CHOICE2066 : STD_LOGIC; 
  signal mac_control_N81130 : STD_LOGIC; 
  signal mac_control_CHOICE2073 : STD_LOGIC; 
  signal tx_output_CHOICE1742 : STD_LOGIC; 
  signal tx_output_N80998 : STD_LOGIC; 
  signal mac_control_PHY_status_miirw : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE872 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_sts : STD_LOGIC; 
  signal mac_control_CHOICE2093 : STD_LOGIC; 
  signal mac_control_CHOICE2085 : STD_LOGIC; 
  signal mac_control_CHOICE2089 : STD_LOGIC; 
  signal mac_control_N81146 : STD_LOGIC; 
  signal mac_control_CHOICE2096 : STD_LOGIC; 
  signal mac_control_CHOICE2231 : STD_LOGIC; 
  signal mac_control_CHOICE2223 : STD_LOGIC; 
  signal mac_control_CHOICE2227 : STD_LOGIC; 
  signal mac_control_N81142 : STD_LOGIC; 
  signal mac_control_CHOICE2234 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd6 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd5 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd4 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd3 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1789 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0030 : STD_LOGIC; 
  signal rx_input_memio_brdy : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd2 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0031 : STD_LOGIC; 
  signal tx_output_CHOICE1718 : STD_LOGIC; 
  signal tx_output_N81010 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1560 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0027 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0028 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1567 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1563 : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0029 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1546 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1528 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1570 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1574 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1549 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1553 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1577 : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1556 : STD_LOGIC; 
  signal mac_control_N69607 : STD_LOGIC; 
  signal mac_control_N72031 : STD_LOGIC; 
  signal mac_control_n0014 : STD_LOGIC; 
  signal rx_output_denll : STD_LOGIC; 
  signal rx_output_invalid : STD_LOGIC; 
  signal rx_output_ldouten2 : STD_LOGIC; 
  signal mac_control_CHOICE2254 : STD_LOGIC; 
  signal mac_control_N81086 : STD_LOGIC; 
  signal mac_control_CHOICE2257 : STD_LOGIC; 
  signal tx_output_CHOICE1730 : STD_LOGIC; 
  signal tx_output_N81022 : STD_LOGIC; 
  signal mac_control_CHOICE2277 : STD_LOGIC; 
  signal mac_control_CHOICE2269 : STD_LOGIC; 
  signal mac_control_CHOICE2273 : STD_LOGIC; 
  signal mac_control_N81126 : STD_LOGIC; 
  signal mac_control_CHOICE2280 : STD_LOGIC; 
  signal tx_output_CHOICE1706 : STD_LOGIC; 
  signal tx_output_N81002 : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd7 : STD_LOGIC; 
  signal rx_input_memio_n0101 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd5 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd2 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd3 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd1 : STD_LOGIC; 
  signal rx_input_memio_N80990 : STD_LOGIC; 
  signal rx_input_memio_n0030 : STD_LOGIC; 
  signal rx_input_memio_bpen : STD_LOGIC; 
  signal rx_input_memio_n0031 : STD_LOGIC; 
  signal rx_input_endf : STD_LOGIC; 
  signal rx_input_invalid : STD_LOGIC; 
  signal rx_input_memio_CHOICE1113 : STD_LOGIC; 
  signal rx_input_memio_n0032 : STD_LOGIC; 
  signal rx_input_memio_CHOICE1979 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd10 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd15 : STD_LOGIC; 
  signal rx_input_memio_N70855 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd14 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd12 : STD_LOGIC; 
  signal rx_input_memio_n0046 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd13 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd9 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd8 : STD_LOGIC; 
  signal rx_input_memio_n0047 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd7 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_292 : STD_LOGIC; 
  signal mac_control_bitcnt_109 : STD_LOGIC; 
  signal mac_control_bitcnt_105 : STD_LOGIC; 
  signal mac_control_bitcnt_108 : STD_LOGIC; 
  signal mac_control_N69675 : STD_LOGIC; 
  signal tx_output_N81026 : STD_LOGIC; 
  signal SCS_IBUF : STD_LOGIC; 
  signal GLOBAL_LOGIC1 : STD_LOGIC; 
  signal GLOBAL_LOGIC0 : STD_LOGIC; 
  signal rx_output_fifo_N10 : STD_LOGIC; 
  signal rx_output_fifo_N1515 : STD_LOGIC; 
  signal rx_output_fifo_N11 : STD_LOGIC; 
  signal rx_output_fifo_N1546 : STD_LOGIC; 
  signal rx_output_fifo_N1547 : STD_LOGIC; 
  signal rx_output_fifo_N2 : STD_LOGIC; 
  signal rx_output_fifo_N1517 : STD_LOGIC; 
  signal rx_output_fifo_N3 : STD_LOGIC; 
  signal rx_output_fifo_N1610 : STD_LOGIC; 
  signal rx_output_fifo_N1611 : STD_LOGIC; 
  signal rx_output_fifo_N1563 : STD_LOGIC; 
  signal rx_output_fifo_N1562 : STD_LOGIC; 
  signal rx_output_fifo_N1551 : STD_LOGIC; 
  signal rx_output_fifo_N1550 : STD_LOGIC; 
  signal rx_output_fifo_N1567 : STD_LOGIC; 
  signal rx_output_fifo_N1566 : STD_LOGIC; 
  signal rx_output_fifo_empty : STD_LOGIC; 
  signal rx_output_fifo_N18 : STD_LOGIC; 
  signal rx_output_fifo_N2579 : STD_LOGIC; 
  signal rx_output_fifo_N1627 : STD_LOGIC; 
  signal rx_output_fifo_N1626 : STD_LOGIC; 
  signal rx_output_ceinll : STD_LOGIC; 
  signal rx_output_fifo_full_0 : STD_LOGIC; 
  signal rx_output_fifo_N19 : STD_LOGIC; 
  signal rx_output_fifo_N3617 : STD_LOGIC; 
  signal memcontroller_n0005 : STD_LOGIC; 
  signal rx_output_fifo_N1549 : STD_LOGIC; 
  signal rx_output_fifo_N1548 : STD_LOGIC; 
  signal rx_output_fifo_N1565 : STD_LOGIC; 
  signal rx_output_fifo_N1564 : STD_LOGIC; 
  signal rx_output_fifo_N1553 : STD_LOGIC; 
  signal rx_output_fifo_N1552 : STD_LOGIC; 
  signal rx_output_fifo_N1569 : STD_LOGIC; 
  signal rx_output_fifo_N1568 : STD_LOGIC; 
  signal rx_output_fifo_N1613 : STD_LOGIC; 
  signal rx_output_fifo_N1612 : STD_LOGIC; 
  signal rx_output_fifo_N1629 : STD_LOGIC; 
  signal rx_output_fifo_N1628 : STD_LOGIC; 
  signal rx_output_fifo_N1617 : STD_LOGIC; 
  signal rx_output_fifo_N1616 : STD_LOGIC; 
  signal rx_output_fifo_N1633 : STD_LOGIC; 
  signal rx_output_fifo_N1632 : STD_LOGIC; 
  signal rx_output_fifo_N1615 : STD_LOGIC; 
  signal rx_output_fifo_N1614 : STD_LOGIC; 
  signal rx_output_fifo_N1631 : STD_LOGIC; 
  signal rx_output_fifo_N1630 : STD_LOGIC; 
  signal rx_output_fifo_N1573 : STD_LOGIC; 
  signal rx_output_fifo_N1572 : STD_LOGIC; 
  signal rx_output_fifo_N1577 : STD_LOGIC; 
  signal rx_output_fifo_N1576 : STD_LOGIC; 
  signal mac_control_PHY_status_n0019 : STD_LOGIC; 
  signal rx_output_fifo_N1575 : STD_LOGIC; 
  signal rx_output_fifo_N1574 : STD_LOGIC; 
  signal clken3 : STD_LOGIC; 
  signal rx_output_fifo_N5 : STD_LOGIC; 
  signal rx_output_fifo_N4 : STD_LOGIC; 
  signal rx_output_fifo_N1605 : STD_LOGIC; 
  signal rx_output_fifo_N1604 : STD_LOGIC; 
  signal rx_output_fifo_N9 : STD_LOGIC; 
  signal rx_output_fifo_N8 : STD_LOGIC; 
  signal rx_output_fifo_N1609 : STD_LOGIC; 
  signal rx_output_fifo_N1608 : STD_LOGIC; 
  signal mac_control_PHY_status_n0020 : STD_LOGIC; 
  signal memcontroller_n0006 : STD_LOGIC; 
  signal rx_output_fifo_N1585 : STD_LOGIC; 
  signal rx_output_fifo_N1584 : STD_LOGIC; 
  signal rx_output_fifo_N1571 : STD_LOGIC; 
  signal rx_output_fifo_N1570 : STD_LOGIC; 
  signal rx_output_fifo_N1578 : STD_LOGIC; 
  signal rx_output_fifo_N1579 : STD_LOGIC; 
  signal rx_output_fifo_N1586 : STD_LOGIC; 
  signal rx_output_fifo_N1587 : STD_LOGIC; 
  signal rx_output_fifo_N1582 : STD_LOGIC; 
  signal rx_output_fifo_N1583 : STD_LOGIC; 
  signal rx_output_fifo_N3959 : STD_LOGIC; 
  signal rx_output_fifo_N1591 : STD_LOGIC; 
  signal rx_output_fifo_N3958 : STD_LOGIC; 
  signal rx_output_fifo_N1603 : STD_LOGIC; 
  signal rx_output_fifo_N1602 : STD_LOGIC; 
  signal rx_output_fifo_N7 : STD_LOGIC; 
  signal rx_output_fifo_N6 : STD_LOGIC; 
  signal rx_output_fifo_N1607 : STD_LOGIC; 
  signal rx_output_fifo_N1606 : STD_LOGIC; 
  signal rx_output_fifo_N1581 : STD_LOGIC; 
  signal rx_output_fifo_N1580 : STD_LOGIC; 
  signal memcontroller_clknum_0_1 : STD_LOGIC; 
  signal memcontroller_clknum_1_1 : STD_LOGIC; 
  signal tx_output_cs_FFd17 : STD_LOGIC; 
  signal clken2 : STD_LOGIC; 
  signal tx_output_n0006 : STD_LOGIC; 
  signal tx_output_CHOICE1694 : STD_LOGIC; 
  signal tx_output_N81006 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd4 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N70564 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0013 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_192 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd5 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0010 : STD_LOGIC; 
  signal tx_output_crc_10_Q : STD_LOGIC; 
  signal rx_output_lmasell : STD_LOGIC; 
  signal tx_input_enable : STD_LOGIC; 
  signal rx_input_memio_n0034 : STD_LOGIC; 
  signal rx_input_memio_crc_0_Q : STD_LOGIC; 
  signal rx_input_memio_crc_2_Q : STD_LOGIC; 
  signal rx_input_memio_crc_3_Q : STD_LOGIC; 
  signal tx_output_N81018 : STD_LOGIC; 
  signal tx_fifocheck_n0002 : STD_LOGIC; 
  signal tx_output_CHOICE1658 : STD_LOGIC; 
  signal tx_output_N81014 : STD_LOGIC; 
  signal tx_output_bcnt_40 : STD_LOGIC; 
  signal tx_output_bcnt_39 : STD_LOGIC; 
  signal tx_output_bcnt_41 : STD_LOGIC; 
  signal tx_output_crc_11_Q : STD_LOGIC; 
  signal tx_output_N70308 : STD_LOGIC; 
  signal rx_input_GMII_dvdelta : STD_LOGIC; 
  signal rx_input_GMII_endf : STD_LOGIC; 
  signal rx_input_GMII_ro : STD_LOGIC; 
  signal rx_input_memio_crc_4_Q : STD_LOGIC; 
  signal tx_output_N70281 : STD_LOGIC; 
  signal tx_output_N70254 : STD_LOGIC; 
  signal mac_control_Mshreg_sinlll_102 : STD_LOGIC; 
  signal tx_output_N70227 : STD_LOGIC; 
  signal tx_output_N70079 : STD_LOGIC; 
  signal tx_input_cs_FFd9 : STD_LOGIC; 
  signal tx_input_cs_FFd12 : STD_LOGIC; 
  signal tx_input_cs_FFd5 : STD_LOGIC; 
  signal tx_input_n0033 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_sout : STD_LOGIC; 
  signal SIN_IBUF : STD_LOGIC; 
  signal tx_input_newframel : STD_LOGIC; 
  signal CLKIN_IBUFG : STD_LOGIC; 
  signal memcontroller_n0149 : STD_LOGIC; 
  signal RX_CLK_IBUFG : STD_LOGIC; 
  signal rx_input_GMII_rx_erl : STD_LOGIC; 
  signal rx_input_GMII_rx_dvl : STD_LOGIC; 
  signal CLKIOIN_IBUFG : STD_LOGIC; 
  signal mac_control_n0034 : STD_LOGIC; 
  signal clkio_to_bufg : STD_LOGIC; 
  signal clk_to_bufg : STD_LOGIC; 
  signal clkrx_to_bufg : STD_LOGIC; 
  signal rx_input_endfin : STD_LOGIC; 
  signal rx_output_fifo_N12 : STD_LOGIC; 
  signal rx_output_fifo_N13 : STD_LOGIC; 
  signal rx_output_fifo_N14 : STD_LOGIC; 
  signal rx_output_fifo_N15 : STD_LOGIC; 
  signal rx_output_fifo_N16 : STD_LOGIC; 
  signal rx_output_fifo_N17 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE977 : STD_LOGIC; 
  signal memcontroller_clknum_1_3 : STD_LOGIC; 
  signal memcontroller_clknum_1_2 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_182 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_184 : STD_LOGIC; 
  signal tx_output_addrinc : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_1 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_3 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_5 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_7 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_9 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_11 : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_13 : STD_LOGIC; 
  signal rx_input_memio_n0102 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_271 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_2 : STD_LOGIC; 
  signal rx_input_memio_bcnt_86 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_273 : STD_LOGIC; 
  signal rx_input_memio_bcnt_87 : STD_LOGIC; 
  signal rx_input_memio_bcnt_88 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_237 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_275 : STD_LOGIC; 
  signal rx_input_memio_bcnt_89 : STD_LOGIC; 
  signal rx_input_memio_bcnt_90 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_277 : STD_LOGIC; 
  signal rx_input_memio_bcnt_91 : STD_LOGIC; 
  signal rx_input_memio_bcnt_92 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_279 : STD_LOGIC; 
  signal rx_input_memio_bcnt_93 : STD_LOGIC; 
  signal rx_input_memio_bcnt_94 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_281 : STD_LOGIC; 
  signal rx_input_memio_bcnt_95 : STD_LOGIC; 
  signal rx_input_memio_bcnt_96 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_283 : STD_LOGIC; 
  signal rx_input_memio_bcnt_97 : STD_LOGIC; 
  signal rx_input_memio_bcnt_98 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_285 : STD_LOGIC; 
  signal rx_input_memio_bcnt_99 : STD_LOGIC; 
  signal rx_input_memio_bcnt_100 : STD_LOGIC; 
  signal rx_input_memio_bcnt_101 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_49 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_51 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_53 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_55 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_57 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_59 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_61 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178 : STD_LOGIC; 
  signal rxcrcerr : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_rxcrcerr_rst : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_222 : STD_LOGIC; 
  signal rx_input_memio_macnt_70 : STD_LOGIC; 
  signal rx_input_memio_macnt_71 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_224 : STD_LOGIC; 
  signal rx_input_memio_macnt_72 : STD_LOGIC; 
  signal rx_input_memio_macnt_73 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_226 : STD_LOGIC; 
  signal rx_input_memio_macnt_74 : STD_LOGIC; 
  signal rx_input_memio_macnt_75 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_228 : STD_LOGIC; 
  signal rx_input_memio_macnt_76 : STD_LOGIC; 
  signal rx_input_memio_macnt_77 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_230 : STD_LOGIC; 
  signal rx_input_memio_macnt_78 : STD_LOGIC; 
  signal rx_input_memio_macnt_79 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_232 : STD_LOGIC; 
  signal rx_input_memio_macnt_80 : STD_LOGIC; 
  signal rx_input_memio_macnt_81 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_234 : STD_LOGIC; 
  signal rx_input_memio_macnt_82 : STD_LOGIC; 
  signal rx_input_memio_macnt_83 : STD_LOGIC; 
  signal rx_input_memio_macnt_84 : STD_LOGIC; 
  signal rx_input_memio_macnt_85 : STD_LOGIC; 
  signal rxoferr : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_rxoferr_rst : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_341 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_343 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_345 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_347 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_349 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_351 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_195 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_197 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_199 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_201 : STD_LOGIC; 
  signal tx_output_n0035 : STD_LOGIC; 
  signal rxphyerr : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_rxphyerr_rst : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal rxfifowerr : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_rxfifowerr_rst : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal txfifowerr : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_txfifowerr_rst : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_87 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_89 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_91 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_93 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_95 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_97 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_99 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_205 : STD_LOGIC; 
  signal tx_output_bcnt_38 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_207 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_209 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_211 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_213 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_215 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_217 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_79 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_81 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_83 : STD_LOGIC; 
  signal rx_output_n0017 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_162 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_164 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_166 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_168 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_170 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_172 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_174 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_162 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_164 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_166 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_168 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_170 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_172 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_174 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_328 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_330 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_332 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_334 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_336 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_338 : STD_LOGIC; 
  signal rx_output_fifo_N1919 : STD_LOGIC; 
  signal rx_output_fifo_N1929 : STD_LOGIC; 
  signal rx_output_fifo_N1939 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_119 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_121 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_123 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_125 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_127 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_129 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_131 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_188 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_32 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_190 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_34 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_36 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_79 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_81 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_83 : STD_LOGIC; 
  signal txf : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_txf_rst : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal rx_output_n0043 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_102 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_104 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_106 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_108 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_110 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_112 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_114 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_116 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_152 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_154 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_156 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_158 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_152 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_154 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_156 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_158 : STD_LOGIC; 
  signal tx_fifocheck_n0003 : STD_LOGIC; 
  signal mac_control_n0032 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_295 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_297 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_299 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_301 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_303 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_305 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_307 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_309 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_311 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_313 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_315 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_317 : STD_LOGIC; 
  signal mac_control_phyrstcnt_131 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_319 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_321 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_323 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_325 : STD_LOGIC; 
  signal mac_control_phyrstcnt_141 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_254 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_256 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_221 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_258 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_260 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_262 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_264 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_266 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_268 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_64 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_66 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_68 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_70 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_72 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_74 : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_76 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_79 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_81 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_83 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_238 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_240 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_242 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_244 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_246 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_248 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_250 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_135 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_137 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_139 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_141 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_143 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_145 : STD_LOGIC; 
  signal tx_input_addr_26 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_147 : STD_LOGIC; 
  signal tx_input_addr_27 : STD_LOGIC; 
  signal tx_input_addr_28 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_149 : STD_LOGIC; 
  signal tx_input_addr_29 : STD_LOGIC; 
  signal tx_input_addr_30 : STD_LOGIC; 
  signal tx_input_addr_31 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_17 : STD_LOGIC; 
  signal mac_control_rxf_rst : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_19 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_21 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_23 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_25 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_27 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_29 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_31 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_33 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_35 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_37 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_39 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_41 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_43 : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_45 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178 : STD_LOGIC; 
  signal rx_output_fifo_N2847 : STD_LOGIC; 
  signal rx_output_fifo_N2857 : STD_LOGIC; 
  signal rx_output_fifo_N2867 : STD_LOGIC; 
  signal rx_output_fifo_N2576 : STD_LOGIC; 
  signal rx_output_fifo_N2574 : STD_LOGIC; 
  signal rx_output_fifo_N2572 : STD_LOGIC; 
  signal rx_output_fifo_BU172_O : STD_LOGIC; 
  signal rx_output_fifo_N3614 : STD_LOGIC; 
  signal rx_output_fifo_N3612 : STD_LOGIC; 
  signal rx_output_fifo_N3610 : STD_LOGIC; 
  signal rx_output_fifo_BU351_O : STD_LOGIC; 
  signal rx_output_fifo_N4763 : STD_LOGIC; 
  signal rx_output_fifo_N1593 : STD_LOGIC; 
  signal rx_output_fifo_N1592 : STD_LOGIC; 
  signal rx_output_fifo_N4771 : STD_LOGIC; 
  signal rx_output_fifo_N1590 : STD_LOGIC; 
  signal rx_output_fifo_N4779 : STD_LOGIC; 
  signal rx_output_fifo_N1589 : STD_LOGIC; 
  signal rx_output_fifo_N1588 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_288 : STD_LOGIC; 
  signal mac_control_bitcnt_104 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_290 : STD_LOGIC; 
  signal mac_control_bitcnt_106 : STD_LOGIC; 
  signal mac_control_bitcnt_107 : STD_LOGIC; 
  signal tx_output_crc_15_Q : STD_LOGIC; 
  signal rx_input_memio_crc_15_Q : STD_LOGIC; 
  signal rx_input_memio_crc_12_Q : STD_LOGIC; 
  signal rx_input_memio_crcen : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O : STD_LOGIC; 
  signal rx_input_memio_n0016 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd15_In6_O : STD_LOGIC; 
  signal rx_input_memio_cs_Out910_O : STD_LOGIC; 
  signal rx_input_memio_cs_FFd6 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd5 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd2 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd4 : STD_LOGIC; 
  signal mac_control_PHY_status_done : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd3 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd6 : STD_LOGIC; 
  signal mac_control_PHY_status_n0019_SW0_O : STD_LOGIC; 
  signal tx_input_Ker3585921_O : STD_LOGIC; 
  signal tx_input_CHOICE1998 : STD_LOGIC; 
  signal tx_input_CHOICE1999 : STD_LOGIC; 
  signal tx_output_crc_5_Q : STD_LOGIC; 
  signal tx_input_CHOICE2029 : STD_LOGIC; 
  signal tx_input_CHOICE2022 : STD_LOGIC; 
  signal tx_input_Ker35859120_O : STD_LOGIC; 
  signal tx_input_N35861 : STD_LOGIC; 
  signal rx_input_memio_crc_5_Q : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_n0005_Result1_O : STD_LOGIC; 
  signal rx_output_n0046_10_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_11_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_12_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_13_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_14_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_15_SW0_O : STD_LOGIC; 
  signal tx_input_N35872 : STD_LOGIC; 
  signal tx_input_cs_FFd10 : STD_LOGIC; 
  signal tx_output_crc_1_Q : STD_LOGIC; 
  signal rx_output_n0046_2_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_3_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_4_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_5_SW0_O : STD_LOGIC; 
  signal tx_output_cs_FFd5 : STD_LOGIC; 
  signal tx_output_cs_FFd6 : STD_LOGIC; 
  signal tx_output_decbcnt : STD_LOGIC; 
  signal rx_output_n0046_6_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_7_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_8_SW0_O : STD_LOGIC; 
  signal rx_output_n0046_9_SW0_O : STD_LOGIC; 
  signal rx_input_memio_n001618_O : STD_LOGIC; 
  signal rx_output_n0043_SW1_O : STD_LOGIC; 
  signal mac_control_n0085 : STD_LOGIC; 
  signal mac_control_PHY_status_n00181_O : STD_LOGIC; 
  signal tx_input_cs_FFd8 : STD_LOGIC; 
  signal rx_input_memio_crc_1_Q : STD_LOGIC; 
  signal mac_control_PHY_status_n00171_O : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd1 : STD_LOGIC; 
  signal tx_output_addrinc_SW0_O : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_n0005_Result1_O : STD_LOGIC; 
  signal mac_control_N53194 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd11 : STD_LOGIC; 
  signal rx_input_memio_wbpl : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd6 : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd8 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_In : STD_LOGIC; 
  signal rx_input_memio_CHOICE1112 : STD_LOGIC; 
  signal tx_input_enableint : STD_LOGIC; 
  signal tx_input_enableintl : STD_LOGIC; 
  signal mac_control_PHY_status_phyaddrws : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd7 : STD_LOGIC; 
  signal rx_input_GMII_rx_dvll : STD_LOGIC; 
  signal tx_output_cs_FFd16_In : STD_LOGIC; 
  signal memcontroller_oe : STD_LOGIC; 
  signal rxfifofull : STD_LOGIC; 
  signal rx_output_cs_FFd18 : STD_LOGIC; 
  signal rx_output_nfl : STD_LOGIC; 
  signal tx_input_newfint : STD_LOGIC; 
  signal tx_input_N70883 : STD_LOGIC; 
  signal mac_control_txf_cross : STD_LOGIC; 
  signal tx_output_cs_FFd5_In : STD_LOGIC; 
  signal tx_output_cs_FFd6_In : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_10_59 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_11_58 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_12_57 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_13_56 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_14_55 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_15_54 : STD_LOGIC; 
  signal tx_output_crc_13_Q : STD_LOGIC; 
  signal rx_input_memio_crc_6_Q : STD_LOGIC; 
  signal tx_output_crc_30_Q : STD_LOGIC; 
  signal tx_output_crc_14_Q : STD_LOGIC; 
  signal rx_input_memio_crc_7_Q : STD_LOGIC; 
  signal rx_input_fifo_control_N70466 : STD_LOGIC; 
  signal rx_input_memio_cs_FFd4 : STD_LOGIC; 
  signal tx_output_crc_23_Q : STD_LOGIC; 
  signal rx_input_memio_crc_10_Q : STD_LOGIC; 
  signal rx_input_memio_crc_8_Q : STD_LOGIC; 
  signal tx_output_crc_24_Q : STD_LOGIC; 
  signal tx_output_crc_16_Q : STD_LOGIC; 
  signal rx_input_memio_crc_11_Q : STD_LOGIC; 
  signal mac_control_PHY_status_N43105 : STD_LOGIC; 
  signal rx_input_memio_crc_9_Q : STD_LOGIC; 
  signal tx_output_crc_25_Q : STD_LOGIC; 
  signal tx_output_crc_17_Q : STD_LOGIC; 
  signal rx_input_memio_addrchk_N70362 : STD_LOGIC; 
  signal rx_input_memio_addrchk_validbcast : STD_LOGIC; 
  signal rx_input_memio_addrchk_N70335 : STD_LOGIC; 
  signal rx_input_memio_addrchk_validucast : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxbcastl : STD_LOGIC; 
  signal rx_input_memio_addrchk_validmcast : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxmcastl : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxallfl : STD_LOGIC; 
  signal rx_input_memio_addrchk_N72932 : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxucastl : STD_LOGIC; 
  signal rx_input_memio_destok : STD_LOGIC; 
  signal rx_output_CHOICE1797 : STD_LOGIC; 
  signal tx_output_crc_18_Q : STD_LOGIC; 
  signal tx_output_crc_26_Q : STD_LOGIC; 
  signal mac_control_lrxallf : STD_LOGIC; 
  signal rx_input_memio_crc_13_Q : STD_LOGIC; 
  signal tx_output_crc_27_Q : STD_LOGIC; 
  signal rx_output_CHOICE1110 : STD_LOGIC; 
  signal rx_input_memio_crc_30_Q : STD_LOGIC; 
  signal rx_input_memio_crc_14_Q : STD_LOGIC; 
  signal tx_input_N70123 : STD_LOGIC; 
  signal mac_control_CHOICE2745 : STD_LOGIC; 
  signal mac_control_N81058 : STD_LOGIC; 
  signal mac_control_CHOICE2750 : STD_LOGIC; 
  signal mac_control_CHOICE2486 : STD_LOGIC; 
  signal mac_control_CHOICE2490 : STD_LOGIC; 
  signal mac_control_CHOICE2753 : STD_LOGIC; 
  signal mac_control_CHOICE2586 : STD_LOGIC; 
  signal mac_control_CHOICE2494 : STD_LOGIC; 
  signal mac_control_N81110 : STD_LOGIC; 
  signal mac_control_CHOICE2497 : STD_LOGIC; 
  signal tx_output_crc_28_Q : STD_LOGIC; 
  signal mac_control_CHOICE2561 : STD_LOGIC; 
  signal mac_control_CHOICE2544 : STD_LOGIC; 
  signal mac_control_N81138 : STD_LOGIC; 
  signal mac_control_CHOICE2547 : STD_LOGIC; 
  signal mac_control_CHOICE2590 : STD_LOGIC; 
  signal mac_control_CHOICE2565 : STD_LOGIC; 
  signal mac_control_CHOICE2767 : STD_LOGIC; 
  signal mac_control_CHOICE2569 : STD_LOGIC; 
  signal mac_control_N81082 : STD_LOGIC; 
  signal mac_control_CHOICE2572 : STD_LOGIC; 
  signal mac_control_CHOICE2771 : STD_LOGIC; 
  signal mac_control_N81042 : STD_LOGIC; 
  signal mac_control_CHOICE2776 : STD_LOGIC; 
  signal mac_control_CHOICE2039 : STD_LOGIC; 
  signal mac_control_CHOICE2779 : STD_LOGIC; 
  signal mac_control_CHOICE2046 : STD_LOGIC; 
  signal mac_control_CHOICE2594 : STD_LOGIC; 
  signal mac_control_N81118 : STD_LOGIC; 
  signal mac_control_CHOICE2048 : STD_LOGIC; 
  signal mac_control_N81176 : STD_LOGIC; 
  signal mac_control_CHOICE2597 : STD_LOGIC; 
  signal rx_input_memio_crc_23_Q : STD_LOGIC; 
  signal rxallf : STD_LOGIC; 
  signal tx_output_crc_29_Q : STD_LOGIC; 
  signal rx_input_memio_crc_24_Q : STD_LOGIC; 
  signal rx_input_memio_crc_16_Q : STD_LOGIC; 
  signal mac_control_n0011 : STD_LOGIC; 
  signal mac_control_PHY_status_n00151_O : STD_LOGIC; 
  signal mac_control_phyaddrw : STD_LOGIC; 
  signal mac_control_N53159 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE963 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE964 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE980 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81411 : STD_LOGIC; 
  signal rx_input_memio_crc_25_Q : STD_LOGIC; 
  signal tx_output_N72900 : STD_LOGIC; 
  signal rx_input_memio_crc_17_Q : STD_LOGIC; 
  signal tx_output_N70101 : STD_LOGIC; 
  signal memcontroller_oel : STD_LOGIC; 
  signal rx_output_N71130 : STD_LOGIC; 
  signal mac_control_PHY_status_start : STD_LOGIC; 
  signal rx_input_memio_addrchk_N80994 : STD_LOGIC; 
  signal rx_input_memio_crc_18_Q : STD_LOGIC; 
  signal rx_input_memio_crc_26_Q : STD_LOGIC; 
  signal rx_input_fifo_control_celll : STD_LOGIC; 
  signal rx_input_memio_crc_27_Q : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81407 : STD_LOGIC; 
  signal rx_input_fifo_control_cell : STD_LOGIC; 
  signal rx_input_memio_crc_28_Q : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE921 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE935 : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1918 : STD_LOGIC; 
  signal rx_input_memio_crc_29_Q : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1925 : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1940 : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1933 : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1941 : STD_LOGIC; 
  signal rx_input_memio_fifofulll : STD_LOGIC; 
  signal rx_input_memio_N70157 : STD_LOGIC; 
  signal rx_input_memio_N70191 : STD_LOGIC; 
  signal mac_control_CHOICE1404 : STD_LOGIC; 
  signal mac_control_CHOICE1407 : STD_LOGIC; 
  signal mac_control_CHOICE1356 : STD_LOGIC; 
  signal mac_control_CHOICE1364 : STD_LOGIC; 
  signal mac_control_CHOICE1371 : STD_LOGIC; 
  signal mac_control_CHOICE1373 : STD_LOGIC; 
  signal mac_control_N80967 : STD_LOGIC; 
  signal tx_output_CHOICE1767 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81171 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE915 : STD_LOGIC; 
  signal tx_output_crc_3_Q : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81405 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE944 : STD_LOGIC; 
  signal tx_output_crc_4_Q : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81167 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_0 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_1 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_2 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_3 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_4 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_5 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_6 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_7 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_8 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_9 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_10 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_11 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_12 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_13 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_14 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_15 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_16 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_17 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_18 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_19 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_20 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_21 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_22 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_23 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_24 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_25 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_26 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_27 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_28 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_29 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_30 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_31 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_32 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_33 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_34 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_35 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_36 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_37 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_38 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_39 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_40 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_41 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_42 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_43 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_44 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_45 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_46 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_47 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_48 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_49 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_0 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_1 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_2 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_3 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_4 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_5 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_6 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_7 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_8 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_9 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_10 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_11 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_12 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_13 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_14 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_15 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_16 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_17 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_18 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_19 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_20 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_21 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_22 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_23 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_24 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_25 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_26 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_27 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_28 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_29 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_30 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_31 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_32 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_33 : STD_LOGIC; 
  signal GSR : STD_LOGIC; 
  signal GTS : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1559_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1552_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1573_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1538_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1497_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1497_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_full_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_full_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3358 : STD_LOGIC; 
  signal rx_input_fifo_fifo_full_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_BU317_O : STD_LOGIC; 
  signal rx_input_fifo_fifo_full_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3374 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1580_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3239 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2721 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2690 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1545_FFX_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1545_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3360 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1545_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3359 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3367 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1545_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1545_CYINIT : STD_LOGIC; 
  signal rx_input_rx_nearf_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4324 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4297 : STD_LOGIC; 
  signal rx_input_rx_nearf_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1582_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3159 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3199 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2711 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2688 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2716 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2713 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2689 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1547_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3362 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1547_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3361 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3369 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1547_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1547_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1574_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4314 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4321_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4318 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4317 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4321_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3689 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3688 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3079 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3119 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2701 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2686 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2706 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2703 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2687 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1582_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3364 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1549_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3363 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3371 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1549_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1549_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1555_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1576_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4306 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4313_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4310 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4309 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4313_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1562_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3686 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1539_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2999 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3039 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2691 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2684 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N8_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2696 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2693 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N8_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N8_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2685 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1550_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1578_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4298 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4305_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4302 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4301 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4305_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3684 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N3685 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1495_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1495_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1794 : STD_LOGIC; 
  signal rx_input_fifo_fifo_empty_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2434 : STD_LOGIC; 
  signal rx_input_fifo_fifo_empty_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_BU156_O : STD_LOGIC; 
  signal rx_input_fifo_fifo_empty_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2450 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2412 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1894 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1863 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N9_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2436 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1594_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2435 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2443 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1594_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1594_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2372 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2332 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1884 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1861 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1889 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1886 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1862 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2438 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1596_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2437 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2445 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1596_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1596_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2292 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2252 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1874 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1859 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N13_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1879 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1876 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N13_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1860 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2440 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1598_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2439 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2447 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1598_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1598_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2172 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N2212 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1864 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1857 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15_CYMUXG : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1869 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1866 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1858 : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1599_GROM : STD_LOGIC; 
  signal rx_input_memio_N80955_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1553_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcrst_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcrst_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N4_FFX_RST : STD_LOGIC; 
  signal mac_control_sclkll_FFY_RST : STD_LOGIC; 
  signal mac_control_sclkll_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE1101_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE1101_GROM : STD_LOGIC; 
  signal txfbbp_11_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_dout_3_FFY_RST : STD_LOGIC; 
  signal txfbbp_13_FFY_RST : STD_LOGIC; 
  signal txfbbp_13_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_15_FFY_RST : STD_LOGIC; 
  signal txfbbp_15_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_dout_7_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N38617_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N38617_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1623_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1623_GROM : STD_LOGIC; 
  signal rx_output_cs_FFd5_In : STD_LOGIC; 
  signal rx_output_cs_FFd5_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1602_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1602_GROM : STD_LOGIC; 
  signal rx_input_data_0_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1630_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1630_GROM : STD_LOGIC; 
  signal rx_input_data_1_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1871_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1595_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1595_GROM : STD_LOGIC; 
  signal rx_input_data_2_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1539_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_55 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_186 : STD_LOGIC; 
  signal tx_output_bcnt_53_GROM : STD_LOGIC; 
  signal tx_output_bcnt_53_CYINIT : STD_LOGIC; 
  signal rx_input_data_3_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1879_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1609_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1609_GROM : STD_LOGIC; 
  signal tx_output_cs_FFd4_FROM : STD_LOGIC; 
  signal tx_output_cs_FFd4_GROM : STD_LOGIC; 
  signal rx_input_data_4_FROM : STD_LOGIC; 
  signal rx_input_data_5_FROM : STD_LOGIC; 
  signal rx_input_data_6_FROM : STD_LOGIC; 
  signal rx_input_data_7_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd3_In : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd3_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1598_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_CHOICE1598_GROM : STD_LOGIC; 
  signal rx_output_cs_FFd9_FROM : STD_LOGIC; 
  signal rx_output_cs_FFd9_In : STD_LOGIC; 
  signal tx_output_crcl_6_FROM : STD_LOGIC; 
  signal tx_output_n0034_6_1_O : STD_LOGIC; 
  signal mac_control_N53109_FROM : STD_LOGIC; 
  signal mac_control_N53109_GROM : STD_LOGIC; 
  signal mac_control_N53144_FROM : STD_LOGIC; 
  signal mac_control_N53144_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd2_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd2_In : STD_LOGIC; 
  signal macaddr_3_FFY_RST : STD_LOGIC; 
  signal macaddr_5_FFY_RST : STD_LOGIC; 
  signal macaddr_9_FFY_RST : STD_LOGIC; 
  signal tx_output_crc_loigc_n0122_1_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0122_1_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1547_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_7_FROM : STD_LOGIC; 
  signal tx_output_n0034_7_Q : STD_LOGIC; 
  signal tx_input_N80947_FROM : STD_LOGIC; 
  signal tx_input_N80947_GROM : STD_LOGIC; 
  signal tx_input_CHOICE2014_FROM : STD_LOGIC; 
  signal tx_input_CHOICE2014_GROM : STD_LOGIC; 
  signal mac_control_dout_1_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_din_1_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1553_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_7_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_10_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_10_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_11_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_11_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_21_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_21_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_13_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_13_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_31_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_31_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_23_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_23_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_15_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_15_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_25_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_17_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_17_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_27_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_27_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_19_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_29_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_29_CEMUXNOT : STD_LOGIC; 
  signal mac_control_dout_2_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_2_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_18_Xo_0_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_18_Xo_0_GROM : STD_LOGIC; 
  signal tx_input_fifofulll_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1574_FFX_SET : STD_LOGIC; 
  signal mac_control_dout_3_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_3_FROM : STD_LOGIC; 
  signal tx_output_crcl_8_FROM : STD_LOGIC; 
  signal tx_output_n0034_8_1_O : STD_LOGIC; 
  signal mac_control_CLKSL_5_FROM : STD_LOGIC; 
  signal mac_control_CLKSL_5_GROM : STD_LOGIC; 
  signal mac_control_CLKSL_4_FROM : STD_LOGIC; 
  signal mac_control_CLKSL_4_GROM : STD_LOGIC; 
  signal mac_control_CLKSL_3_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1839_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1846_GROM : STD_LOGIC; 
  signal rx_input_memio_crcequal_FROM : STD_LOGIC; 
  signal rx_input_memio_n0059 : STD_LOGIC; 
  signal rx_input_memio_crcequal_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1560_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_n0033_FROM : STD_LOGIC; 
  signal rx_input_memio_n0033_GROM : STD_LOGIC; 
  signal mac_control_dout_4_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_23_Xo_0_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_23_Xo_0_GROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_18_Xo_0_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_18_Xo_0_GROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0122_0_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0122_0_GROM : STD_LOGIC; 
  signal rx_output_fifo_nearfull_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_9_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_9_FROM : STD_LOGIC; 
  signal tx_output_n0034_9_Q : STD_LOGIC; 
  signal mac_control_dout_5_FROM : STD_LOGIC; 
  signal addr4ext_5_FFY_RST : STD_LOGIC; 
  signal addr4ext_7_FFY_RST : STD_LOGIC; 
  signal addr4ext_9_FFY_RST : STD_LOGIC; 
  signal d4_3_FFY_RST : STD_LOGIC; 
  signal d4_5_FFY_RST : STD_LOGIC; 
  signal d4_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1560_FFX_SET : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_11_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1541_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_13_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_15_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd12_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd14_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1584_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd16_FFY_RST : STD_LOGIC; 
  signal rx_output_cein : STD_LOGIC; 
  signal rx_output_ceinl_CEMUXNOT : STD_LOGIC; 
  signal rx_output_ceinl_GROM : STD_LOGIC; 
  signal rx_output_fifo_reset_FROM : STD_LOGIC; 
  signal rx_output_fifo_reset_GROM : STD_LOGIC; 
  signal mac_control_dout_6_FROM : STD_LOGIC; 
  signal tx_input_n0023_FROM : STD_LOGIC; 
  signal tx_input_n0023_GROM : STD_LOGIC; 
  signal mac_control_dout_7_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_2_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_2_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_3_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_5_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_7_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_9_CEMUXNOT : STD_LOGIC; 
  signal mac_control_CHOICE1272_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1272_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1584_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE1387_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1387_GROM : STD_LOGIC; 
  signal mac_control_N80971_FROM : STD_LOGIC; 
  signal mac_control_N80971_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1333_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1333_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1325_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1325_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6_FFY_RST : STD_LOGIC; 
  signal mac_control_CHOICE1399_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1402_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1340_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1340_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1280_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1280_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_7_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_7_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1541_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_9_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_n00061_1_FROM : STD_LOGIC; 
  signal memcontroller_n00061_1_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2634_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2634_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2508_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2508_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2105_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2105_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2243_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2243_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2583_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2583_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2712_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2712_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2174_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2174_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2384_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2384_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2387_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2387_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2082_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2082_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2698_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2698_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1899_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1899_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2660_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2660_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2637_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2637_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2043_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2043_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2408_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2408_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2615_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2615_GROM : STD_LOGIC; 
  signal mac_control_dout_0_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2220_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2220_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1562_FFY_SET : STD_LOGIC; 
  signal mac_control_CHOICE2641_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2641_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2372_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2372_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2623_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2623_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2108_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2108_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2433_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2433_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2296_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2296_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2649_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2649_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1555_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE2246_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2246_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2444_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2444_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2447_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2447_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2715_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2715_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2419_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2419_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2422_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2422_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2667_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2667_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2324_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2324_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2741_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2741_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2693_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2693_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2675_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2675_GROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_7_Xo_1_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_7_Xo_1_GROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_9_Xo_0_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_9_Xo_0_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2292_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2292_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_6_FFY_RST : STD_LOGIC; 
  signal mac_control_CHOICE1283_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1283_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1311_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1311_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_10_FFY_RST : STD_LOGIC; 
  signal mac_control_CHOICE1269_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1269_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1297_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1297_GROM : STD_LOGIC; 
  signal mac_control_dout_8_FROM : STD_LOGIC; 
  signal tx_input_dh_3_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crccomb_N81261_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_N81261_GROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_n0124_0_GROM : STD_LOGIC; 
  signal tx_input_dh_9_FFY_RST : STD_LOGIC; 
  signal txbp_1_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_3_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N6_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_7_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_9_FFY_RST : STD_LOGIC; 
  signal MDC_OBUF_FFY_RST : STD_LOGIC; 
  signal MDC_OBUF_CEMUXNOT : STD_LOGIC; 
  signal mac_control_dout_9_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_9_FROM : STD_LOGIC; 
  signal mac_control_lmacaddr_3_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_5_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_7_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_9_FFY_RST : STD_LOGIC; 
  signal rxbp_1_FFX_RST : STD_LOGIC; 
  signal rxbp_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1549_FFY_RST : STD_LOGIC; 
  signal rxbp_3_FFY_RST : STD_LOGIC; 
  signal rxbp_3_FFX_RST : STD_LOGIC; 
  signal rxbp_3_CEMUXNOT : STD_LOGIC; 
  signal rxbp_5_FFY_RST : STD_LOGIC; 
  signal rxbp_5_FFX_RST : STD_LOGIC; 
  signal rxbp_5_CEMUXNOT : STD_LOGIC; 
  signal rxbp_7_FFY_RST : STD_LOGIC; 
  signal rxbp_7_FFX_RST : STD_LOGIC; 
  signal rxbp_7_CEMUXNOT : STD_LOGIC; 
  signal rxbp_9_FFY_RST : STD_LOGIC; 
  signal rxbp_9_FFX_RST : STD_LOGIC; 
  signal rxbp_9_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_3_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_5_CEMUXNOT : STD_LOGIC; 
  signal mac_control_CHOICE2250_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2250_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1576_FFX_SET : STD_LOGIC; 
  signal mac_control_CHOICE2701_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2701_GROM : STD_LOGIC; 
  signal tx_output_crc_loigc_N81257_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_N81257_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1439_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1439_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2469_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2469_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2472_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2472_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2719_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2719_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2396_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2396_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2177_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2177_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2540_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2540_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2727_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2727_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2519_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2519_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2522_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2522_GROM : STD_LOGIC; 
  signal rx_output_CHOICE1800_FROM : STD_LOGIC; 
  signal rx_output_CHOICE1800_GROM : STD_LOGIC; 
  signal rx_output_denl_FROM : STD_LOGIC; 
  signal rx_output_denl_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_CHOICE880 : STD_LOGIC; 
  signal rxbcast_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81159_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81159_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE892_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE892_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE900_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE900_GROM : STD_LOGIC; 
  signal tx_input_mrw_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1525_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1525_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_mcast_0_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_mcast_0_CEMUXNOT : STD_LOGIC; 
  signal tx_output_CHOICE1505_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1505_GROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_0_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_0_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_dout_13_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_15_FFY_RST : STD_LOGIC; 
  signal tx_output_CHOICE1483_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1483_GROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_1_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_ncrcbytel_2_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_2_CEMUXNOT : STD_LOGIC; 
  signal tx_output_ncrcbytel_3_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_3_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1562_FFX_SET : STD_LOGIC; 
  signal tx_output_CHOICE1450_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1450_GROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_n0007_Xo_0_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_n0007_Xo_0_GROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_4_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_4_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crc_loigc_n0118_0_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0118_0_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1586_FFY_RST : STD_LOGIC; 
  signal tx_output_crc_loigc_n0124_1_GROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_5_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_ncrcbytel_6_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_6_CEMUXNOT : STD_LOGIC; 
  signal tx_output_ncrcbytel_7_FROM : STD_LOGIC; 
  signal tx_output_ncrcbytel_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_11_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_11_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N8_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_21_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_21_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_13_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_13_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1586_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_31_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_31_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_23_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_23_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_15_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_15_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_25_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_17_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_17_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_27_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_27_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_19_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_19_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_29_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_29_CEMUXNOT : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1950_GROM : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1957_GROM : STD_LOGIC; 
  signal mac_control_dout_10_FROM : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1972_GROM : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1973_FROM : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1973_GROM : STD_LOGIC; 
  signal rx_fifocheck_CHOICE1965_GROM : STD_LOGIC; 
  signal mac_control_N81102_FROM : STD_LOGIC; 
  signal mac_control_N81102_GROM : STD_LOGIC; 
  signal mac_control_dout_11_FROM : STD_LOGIC; 
  signal rx_input_memio_RESET_1_FROM : STD_LOGIC; 
  signal rx_input_memio_RESET_1_GROM : STD_LOGIC; 
  signal tx_output_n0034_12_1_O : STD_LOGIC; 
  signal tx_output_crcl_12_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1775_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1775_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1682_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1682_GROM : STD_LOGIC; 
  signal tx_output_crcsell_0_GROM : STD_LOGIC; 
  signal tx_output_crcsell_0_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_3_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_5_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_5_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_7_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_9_CEMUXNOT : STD_LOGIC; 
  signal mac_control_dout_12_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_12_FROM : STD_LOGIC; 
  signal mac_control_N81038_FROM : STD_LOGIC; 
  signal mac_control_N81038_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1550_FFY_SET : STD_LOGIC; 
  signal tx_output_crcl_2_FROM : STD_LOGIC; 
  signal tx_output_n0034_2_Q : STD_LOGIC; 
  signal mac_control_N81090_FROM : STD_LOGIC; 
  signal mac_control_N81090_GROM : STD_LOGIC; 
  signal mac_control_N81094_FROM : STD_LOGIC; 
  signal mac_control_N81094_GROM : STD_LOGIC; 
  signal mac_control_dout_13_FROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N8_FFX_RST : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_103_CEMUXNOT : STD_LOGIC; 
  signal rx_input_GMII_rx_of_FFY_RST : STD_LOGIC; 
  signal mac_control_CHOICE2185_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2185_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1543_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_CHOICE1812_GROM : STD_LOGIC; 
  signal mac_control_N81134_FROM : STD_LOGIC; 
  signal mac_control_N81134_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1821_FROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1821_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1817_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1832_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_11_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_21_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_21_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_13_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_13_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_31_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_31_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_23_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_23_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_15_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_15_CEMUXNOT : STD_LOGIC; 
  signal mac_control_dout_14_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_14_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_25_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_17_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_17_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_27_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_27_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_19_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_19_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_29_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_29_CEMUXNOT : STD_LOGIC; 
  signal mac_control_dout_15_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_15_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1670_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1670_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1543_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_3_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_5_FFY_RST : STD_LOGIC; 
  signal mac_control_N81046_FROM : STD_LOGIC; 
  signal mac_control_N81046_GROM : STD_LOGIC; 
  signal mac_control_N81074_FROM : STD_LOGIC; 
  signal mac_control_N81074_GROM : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_11_FFY_RST : STD_LOGIC; 
  signal mac_control_n0015_FROM : STD_LOGIC; 
  signal mac_control_n0015_GROM : STD_LOGIC; 
  signal tx_output_ltxen3_FROM : STD_LOGIC; 
  signal tx_output_ltxen : STD_LOGIC; 
  signal tx_output_ltxen3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_n0024_FROM : STD_LOGIC; 
  signal mac_control_n0024_GROM : STD_LOGIC; 
  signal mac_control_n0025_FROM : STD_LOGIC; 
  signal mac_control_n0025_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1557_FFY_RST : STD_LOGIC; 
  signal mac_control_CHOICE1291_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1291_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1550_FFX_SET : STD_LOGIC; 
  signal mac_control_n0029_FROM : STD_LOGIC; 
  signal mac_control_n0029_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1380_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1380_GROM : STD_LOGIC; 
  signal mac_control_n0060_FROM : STD_LOGIC; 
  signal mac_control_n0060_GROM : STD_LOGIC; 
  signal mac_control_n0036_FROM : STD_LOGIC; 
  signal mac_control_n0036_GROM : STD_LOGIC; 
  signal mac_control_N81098_FROM : STD_LOGIC; 
  signal mac_control_N81098_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1302_GROM : STD_LOGIC; 
  signal mac_control_n0063_FROM : STD_LOGIC; 
  signal mac_control_n0063_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1305_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1305_GROM : STD_LOGIC; 
  signal mac_control_N81417_FROM : STD_LOGIC; 
  signal mac_control_N81417_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1557_FFX_RST : STD_LOGIC; 
  signal mac_control_n0064_FROM : STD_LOGIC; 
  signal mac_control_n0064_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1288_GROM : STD_LOGIC; 
  signal mac_control_n0057_FROM : STD_LOGIC; 
  signal mac_control_n0057_GROM : STD_LOGIC; 
  signal mac_control_n0065_FROM : STD_LOGIC; 
  signal mac_control_n0065_GROM : STD_LOGIC; 
  signal mac_control_n0066_FROM : STD_LOGIC; 
  signal mac_control_n0066_GROM : STD_LOGIC; 
  signal mac_control_N81070_FROM : STD_LOGIC; 
  signal mac_control_N81070_GROM : STD_LOGIC; 
  signal mac_control_N81154_FROM : STD_LOGIC; 
  signal mac_control_N81154_GROM : STD_LOGIC; 
  signal mac_control_N81130_FROM : STD_LOGIC; 
  signal mac_control_N81130_GROM : STD_LOGIC; 
  signal tx_output_data_0_FROM : STD_LOGIC; 
  signal tx_output_data_0_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE872_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE872_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2608_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2608_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2319_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2319_GROM : STD_LOGIC; 
  signal mac_control_N81146_FROM : STD_LOGIC; 
  signal mac_control_N81146_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1578_FFX_SET : STD_LOGIC; 
  signal mac_control_N81142_FROM : STD_LOGIC; 
  signal mac_control_N81142_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1565_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1789_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1789_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd2_In : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd2_GROM : STD_LOGIC; 
  signal tx_output_data_1_FROM : STD_LOGIC; 
  signal tx_output_data_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1560_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd5_In : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd5_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0028_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1567_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_3_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_3_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0029_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1546_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_0_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_0_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_5_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_5_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1574_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_2_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_2_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_CHOICE1553_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_4_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_4_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_1_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_N69607_FROM : STD_LOGIC; 
  signal mac_control_N69607_GROM : STD_LOGIC; 
  signal mac_control_N69759_FROM : STD_LOGIC; 
  signal mac_control_N69759_GROM : STD_LOGIC; 
  signal mac_control_N72031_FROM : STD_LOGIC; 
  signal mac_control_N72031_GROM : STD_LOGIC; 
  signal tx_output_cs_FFd12_FFY_RST : STD_LOGIC; 
  signal mac_control_N81086_FROM : STD_LOGIC; 
  signal mac_control_N81086_GROM : STD_LOGIC; 
  signal tx_output_data_2_FROM : STD_LOGIC; 
  signal tx_output_data_2_CEMUXNOT : STD_LOGIC; 
  signal mac_control_N81126_FROM : STD_LOGIC; 
  signal mac_control_N81126_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1565_FFX_SET : STD_LOGIC; 
  signal tx_output_data_3_FROM : STD_LOGIC; 
  signal tx_output_data_3_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd7_In : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd7_GROM : STD_LOGIC; 
  signal rx_input_memio_N80990_FROM : STD_LOGIC; 
  signal rx_input_memio_N80990_GROM : STD_LOGIC; 
  signal rx_input_memio_n0031_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1113_FROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1113_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1979_GROM : STD_LOGIC; 
  signal rx_input_memio_N70855_FROM : STD_LOGIC; 
  signal rx_input_memio_N70855_GROM : STD_LOGIC; 
  signal rx_input_memio_n0045_GROM : STD_LOGIC; 
  signal rx_input_fifo_dout_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_n0046_GROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd8_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd8_GROM : STD_LOGIC; 
  signal rx_input_memio_CHOICE1808_GROM : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_191 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_256 : STD_LOGIC; 
  signal mac_control_bitcnt_109_GROM : STD_LOGIC; 
  signal mac_control_bitcnt_109_CYINIT : STD_LOGIC; 
  signal tx_output_data_4_FROM : STD_LOGIC; 
  signal tx_output_data_4_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_12_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_14_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_14_FFX_RST : STD_LOGIC; 
  signal tx_output_bcntl_14_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_15_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_15_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_11_FFX_RST : STD_LOGIC; 
  signal rxfbbp_11_FFY_RST : STD_LOGIC; 
  signal rxfbbp_11_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_13_FFY_RST : STD_LOGIC; 
  signal rxfbbp_13_FFX_RST : STD_LOGIC; 
  signal rxfbbp_13_CEMUXNOT : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_net187_GSHIFT : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_net187_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rxfbbp_15_FFX_RST : STD_LOGIC; 
  signal rxfbbp_15_FFY_RST : STD_LOGIC; 
  signal rxfbbp_15_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifo_N1546_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1546_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N2499 : STD_LOGIC; 
  signal rx_input_fifo_fifo_empty_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1610_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N3427 : STD_LOGIC; 
  signal rx_output_fifo_N1563_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1567_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N18_FROM : STD_LOGIC; 
  signal rx_output_fifo_N18_GROM : STD_LOGIC; 
  signal rx_output_fifo_N19_FROM : STD_LOGIC; 
  signal rx_output_fifo_N19_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1565_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1524_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1569_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N1629_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1629_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1633_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1633_FFX_SET : STD_LOGIC; 
  signal q2_21_FFY_RST : STD_LOGIC; 
  signal q2_21_FFX_RST : STD_LOGIC; 
  signal q2_13_FFY_RST : STD_LOGIC; 
  signal q2_13_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1631_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1631_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1573_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1573_FFX_RST : STD_LOGIC; 
  signal q2_31_FFY_RST : STD_LOGIC; 
  signal q2_31_FFX_RST : STD_LOGIC; 
  signal q2_22_FFY_RST : STD_LOGIC; 
  signal q2_15_FFY_RST : STD_LOGIC; 
  signal q2_15_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1577_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1577_FFX_SET : STD_LOGIC; 
  signal q2_23_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_11_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_11_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1575_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1575_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1517_GROM : STD_LOGIC; 
  signal q2_25_FFX_RST : STD_LOGIC; 
  signal q2_25_FFY_RST : STD_LOGIC; 
  signal q2_17_FFY_RST : STD_LOGIC; 
  signal q2_17_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd3_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd3_FROM : STD_LOGIC; 
  signal rx_output_cs_FFd3_In : STD_LOGIC; 
  signal rx_output_fifo_N1605_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1609_FFY_SET : STD_LOGIC; 
  signal mac_control_phystat_21_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_13_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N9_FFX_RST : STD_LOGIC; 
  signal q2_27_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1525_FFY_RST : STD_LOGIC; 
  signal q2_19_FFY_RST : STD_LOGIC; 
  signal q3_11_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1585_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_23_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_31_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_15_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1571_FFY_SET : STD_LOGIC; 
  signal q2_29_FFY_RST : STD_LOGIC; 
  signal q3_21_FFY_RST : STD_LOGIC; 
  signal q3_13_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1586_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N3974 : STD_LOGIC; 
  signal rx_output_fifo_N1591_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N3970 : STD_LOGIC; 
  signal rx_output_fifo_N1591_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1603_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1607_FFY_SET : STD_LOGIC; 
  signal mac_control_phystat_25_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_17_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1594_FFY_RST : STD_LOGIC; 
  signal q3_31_FFY_RST : STD_LOGIC; 
  signal q3_22_FFY_RST : STD_LOGIC; 
  signal memcontroller_n0006_FROM : STD_LOGIC; 
  signal memcontroller_n0006_GROM : STD_LOGIC; 
  signal mac_control_phystat_19_FFY_RST : STD_LOGIC; 
  signal q3_25_FFY_RST : STD_LOGIC; 
  signal q3_17_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_29_FFY_RST : STD_LOGIC; 
  signal q3_27_FFY_RST : STD_LOGIC; 
  signal q3_19_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1581_FFY_RST : STD_LOGIC; 
  signal q3_29_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd17_FFY_SET : STD_LOGIC; 
  signal tx_output_cs_FFd17_FROM : STD_LOGIC; 
  signal tx_output_cs_FFd17_In : STD_LOGIC; 
  signal rx_output_ceinll_CEMUXNOT : STD_LOGIC; 
  signal tx_output_data_5_FROM : STD_LOGIC; 
  signal tx_output_data_5_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd3_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd3_In : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_39 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_170 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_37_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_37_CYINIT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0013_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0013_GROM : STD_LOGIC; 
  signal tx_output_crcl_10_FROM : STD_LOGIC; 
  signal tx_output_n0034_10_Q : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0015_GROM : STD_LOGIC; 
  signal rx_output_mdl_11_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_11_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_21_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_21_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1596_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_13_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_13_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1594_FFX_SET : STD_LOGIC; 
  signal rx_output_mdl_31_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_31_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_23_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_23_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1525_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_15_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_15_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_25_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_17_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_17_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_27_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_27_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_19_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_19_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_29_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_29_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lmasell_FFY_RST : STD_LOGIC; 
  signal rx_output_lmasell_CEMUXNOT : STD_LOGIC; 
  signal tx_input_enable_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_crcl_2_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_2_Q : STD_LOGIC; 
  signal rx_input_memio_crcl_3_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_3_Q : STD_LOGIC; 
  signal tx_output_data_6_FROM : STD_LOGIC; 
  signal tx_output_data_6_CEMUXNOT : STD_LOGIC; 
  signal txfifofull_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_data_7_FROM : STD_LOGIC; 
  signal tx_output_data_7_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_2_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_4_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_4_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_6_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_6_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_1_FFY_RST : STD_LOGIC; 
  signal rxfbbp_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_8_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_8_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_3_FFY_RST : STD_LOGIC; 
  signal rxfbbp_3_CEMUXNOT : STD_LOGIC; 
  signal tx_output_datal_1_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bcntl_10_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_10_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_5_FFY_RST : STD_LOGIC; 
  signal rxfbbp_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_datal_3_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_3_CEMUXNOT : STD_LOGIC; 
  signal rxfbbp_7_FFY_RST : STD_LOGIC; 
  signal rxfbbp_7_CEMUXNOT : STD_LOGIC; 
  signal tx_output_datal_5_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_11_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_11_FROM : STD_LOGIC; 
  signal tx_output_n0034_11_1_O : STD_LOGIC; 
  signal rxfbbp_9_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1527_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_7_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_1_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_3_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_5_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_7_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_9_CEMUXNOT : STD_LOGIC; 
  signal rx_output_denll_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_1_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_fifo_N13_FFY_RST : STD_LOGIC; 
  signal rx_output_len_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_fifo_N11_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_3_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_3_CEMUXNOT : STD_LOGIC; 
  signal rx_output_mdl_5_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_5_CEMUXNOT : STD_LOGIC; 
  signal rx_output_len_7_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_7_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_7_CEMUXNOT : STD_LOGIC; 
  signal rx_output_len_9_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_9_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_9_CEMUXNOT : STD_LOGIC; 
  signal tx_output_N70308_FROM : STD_LOGIC; 
  signal tx_output_N70308_GROM : STD_LOGIC; 
  signal rx_input_GMII_ro_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_crcl_4_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_4_1_O : STD_LOGIC; 
  signal tx_output_outselll_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_outselll_3_FFY_RST : STD_LOGIC; 
  signal tx_output_outselll_3_CEMUXNOT : STD_LOGIC; 
  signal tx_output_N70281_FROM : STD_LOGIC; 
  signal tx_output_N70281_GROM : STD_LOGIC; 
  signal mac_control_txf_cntl_11_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_21_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_21_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_13_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_13_CEMUXNOT : STD_LOGIC; 
  signal tx_output_N70254_FROM : STD_LOGIC; 
  signal tx_output_N70254_GROM : STD_LOGIC; 
  signal mac_control_txf_cntl_31_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_31_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_23_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_23_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_15_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_15_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_25_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_25_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_17_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_17_CEMUXNOT : STD_LOGIC; 
  signal mac_control_addr_0_1_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_27_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_19_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_29_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_29_CEMUXNOT : STD_LOGIC; 
  signal tx_output_CHOICE1730_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1730_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1694_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1694_GROM : STD_LOGIC; 
  signal tx_output_CHOICE1658_FROM : STD_LOGIC; 
  signal tx_output_CHOICE1658_GROM : STD_LOGIC; 
  signal tx_output_N70227_FROM : STD_LOGIC; 
  signal tx_output_N70227_GROM : STD_LOGIC; 
  signal tx_output_N70079_FROM : STD_LOGIC; 
  signal tx_output_N70079_GROM : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1596_FFX_RST : STD_LOGIC; 
  signal RESET_IBUF_1_FROM : STD_LOGIC; 
  signal RESET_IBUF_1_GROM : STD_LOGIC; 
  signal RESET_IBUF_2_FROM : STD_LOGIC; 
  signal RESET_IBUF_2_GROM : STD_LOGIC; 
  signal MDIO_ENABLE : STD_LOGIC; 
  signal MDIO_TORGTS : STD_LOGIC; 
  signal MDIO_OUTMUX : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_sin : STD_LOGIC; 
  signal DOUT_10_ENABLE : STD_LOGIC; 
  signal DOUT_10_TORGTS : STD_LOGIC; 
  signal DOUT_10_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_10_OBUF : STD_LOGIC; 
  signal DOUT_10_OD : STD_LOGIC; 
  signal DOUT_11_ENABLE : STD_LOGIC; 
  signal DOUT_11_TORGTS : STD_LOGIC; 
  signal DOUT_11_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_11_OBUF : STD_LOGIC; 
  signal DOUT_11_OD : STD_LOGIC; 
  signal DOUT_12_ENABLE : STD_LOGIC; 
  signal DOUT_12_TORGTS : STD_LOGIC; 
  signal DOUT_12_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_12_OBUF : STD_LOGIC; 
  signal DOUT_12_OD : STD_LOGIC; 
  signal DOUT_13_ENABLE : STD_LOGIC; 
  signal DOUT_13_TORGTS : STD_LOGIC; 
  signal DOUT_13_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_13_OBUF : STD_LOGIC; 
  signal DOUT_13_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1527_FFX_RST : STD_LOGIC; 
  signal DOUT_14_ENABLE : STD_LOGIC; 
  signal DOUT_14_TORGTS : STD_LOGIC; 
  signal DOUT_14_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_14_OBUF : STD_LOGIC; 
  signal DOUT_14_OD : STD_LOGIC; 
  signal DOUT_15_ENABLE : STD_LOGIC; 
  signal DOUT_15_TORGTS : STD_LOGIC; 
  signal DOUT_15_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_15_OBUF : STD_LOGIC; 
  signal DOUT_15_OD : STD_LOGIC; 
  signal MDC_ENABLE : STD_LOGIC; 
  signal MDC_TORGTS : STD_LOGIC; 
  signal MDC_OUTMUX : STD_LOGIC; 
  signal SCS_IBUF_1 : STD_LOGIC; 
  signal SIN_IBUF_2 : STD_LOGIC; 
  signal LED100_ENABLE : STD_LOGIC; 
  signal LED100_TORGTS : STD_LOGIC; 
  signal LED100_OUTMUX : STD_LOGIC; 
  signal mac_control_LED100_OBUF : STD_LOGIC; 
  signal LED100_OCEMUXNOT : STD_LOGIC; 
  signal LED100_OD : STD_LOGIC; 
  signal MCLK_ENABLE : STD_LOGIC; 
  signal MCLK_TORGTS : STD_LOGIC; 
  signal MCLK_OUTMUX : STD_LOGIC; 
  signal tx_input_NEWFRAME_IBUF : STD_LOGIC; 
  signal LED1000_ENABLE : STD_LOGIC; 
  signal LED1000_TORGTS : STD_LOGIC; 
  signal LED1000_OUTMUX : STD_LOGIC; 
  signal mac_control_LED1000_OBUF : STD_LOGIC; 
  signal LED1000_OCEMUXNOT : STD_LOGIC; 
  signal LED1000_OD : STD_LOGIC; 
  signal TX_EN_ENABLE : STD_LOGIC; 
  signal TX_EN_TORGTS : STD_LOGIC; 
  signal TX_EN_OUTMUX : STD_LOGIC; 
  signal tx_output_TXEN : STD_LOGIC; 
  signal TX_EN_OCEMUXNOT : STD_LOGIC; 
  signal TX_EN_OD : STD_LOGIC; 
  signal DOUTEN_ENABLE : STD_LOGIC; 
  signal DOUTEN_TORGTS : STD_LOGIC; 
  signal DOUTEN_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUTEN_OBUF : STD_LOGIC; 
  signal DOUTEN_OD : STD_LOGIC; 
  signal MWE_ENABLE : STD_LOGIC; 
  signal MWE_TORGTS : STD_LOGIC; 
  signal MWE_OUTMUX : STD_LOGIC; 
  signal memcontroller_we : STD_LOGIC; 
  signal MWE_OD : STD_LOGIC; 
  signal RESET_IBUF_3 : STD_LOGIC; 
  signal rx_output_NEXTFRAME_IBUF : STD_LOGIC; 
  signal LEDACT_ENABLE : STD_LOGIC; 
  signal LEDACT_TORGTS : STD_LOGIC; 
  signal LEDACT_OUTMUX : STD_LOGIC; 
  signal mac_control_LEDACT_OBUF : STD_LOGIC; 
  signal LEDACT_OCEMUXNOT : STD_LOGIC; 
  signal LEDACT_OD : STD_LOGIC; 
  signal TXD_0_ENABLE : STD_LOGIC; 
  signal TXD_0_TORGTS : STD_LOGIC; 
  signal TXD_0_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_0_OBUF : STD_LOGIC; 
  signal TXD_0_OCEMUXNOT : STD_LOGIC; 
  signal TXD_0_OD : STD_LOGIC; 
  signal TXD_1_ENABLE : STD_LOGIC; 
  signal TXD_1_TORGTS : STD_LOGIC; 
  signal TXD_1_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_1_OBUF : STD_LOGIC; 
  signal TXD_1_OCEMUXNOT : STD_LOGIC; 
  signal TXD_1_OD : STD_LOGIC; 
  signal TXD_2_ENABLE : STD_LOGIC; 
  signal TXD_2_TORGTS : STD_LOGIC; 
  signal TXD_2_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_2_OBUF : STD_LOGIC; 
  signal TXD_2_OCEMUXNOT : STD_LOGIC; 
  signal TXD_2_OD : STD_LOGIC; 
  signal TXD_3_ENABLE : STD_LOGIC; 
  signal TXD_3_TORGTS : STD_LOGIC; 
  signal TXD_3_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_3_OBUF : STD_LOGIC; 
  signal TXD_3_OCEMUXNOT : STD_LOGIC; 
  signal TXD_3_OD : STD_LOGIC; 
  signal TXD_4_ENABLE : STD_LOGIC; 
  signal TXD_4_TORGTS : STD_LOGIC; 
  signal TXD_4_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_4_OBUF : STD_LOGIC; 
  signal TXD_4_OCEMUXNOT : STD_LOGIC; 
  signal TXD_4_OD : STD_LOGIC; 
  signal TXD_5_ENABLE : STD_LOGIC; 
  signal TXD_5_TORGTS : STD_LOGIC; 
  signal TXD_5_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_5_OBUF : STD_LOGIC; 
  signal TXD_5_OCEMUXNOT : STD_LOGIC; 
  signal TXD_5_OD : STD_LOGIC; 
  signal TXD_6_ENABLE : STD_LOGIC; 
  signal TXD_6_TORGTS : STD_LOGIC; 
  signal TXD_6_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_6_OBUF : STD_LOGIC; 
  signal TXD_6_OCEMUXNOT : STD_LOGIC; 
  signal TXD_6_OD : STD_LOGIC; 
  signal TXD_7_ENABLE : STD_LOGIC; 
  signal TXD_7_TORGTS : STD_LOGIC; 
  signal TXD_7_OUTMUX : STD_LOGIC; 
  signal tx_output_TXD_7_OBUF : STD_LOGIC; 
  signal TXD_7_OCEMUXNOT : STD_LOGIC; 
  signal TXD_7_OD : STD_LOGIC; 
  signal LEDDPX_ENABLE : STD_LOGIC; 
  signal LEDDPX_TORGTS : STD_LOGIC; 
  signal LEDDPX_OUTMUX : STD_LOGIC; 
  signal mac_control_LEDDPX_OBUF : STD_LOGIC; 
  signal LEDDPX_OCEMUXNOT : STD_LOGIC; 
  signal LEDDPX_OD : STD_LOGIC; 
  signal rx_input_GMII_RXD_0_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_1_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_2_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_3_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_4_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_5_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_6_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RXD_7_IBUF : STD_LOGIC; 
  signal tx_input_DIN_10_IBUF : STD_LOGIC; 
  signal tx_input_DIN_11_IBUF : STD_LOGIC; 
  signal tx_input_DIN_12_IBUF : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1530_FFY_RST : STD_LOGIC; 
  signal tx_input_DIN_13_IBUF : STD_LOGIC; 
  signal rx_input_fifo_fifo_N13_FFX_RST : STD_LOGIC; 
  signal tx_input_DIN_14_IBUF : STD_LOGIC; 
  signal tx_input_DIN_15_IBUF : STD_LOGIC; 
  signal DOUT_0_ENABLE : STD_LOGIC; 
  signal DOUT_0_TORGTS : STD_LOGIC; 
  signal DOUT_0_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_0_OBUF : STD_LOGIC; 
  signal DOUT_0_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1598_FFY_RST : STD_LOGIC; 
  signal DOUT_1_ENABLE : STD_LOGIC; 
  signal DOUT_1_TORGTS : STD_LOGIC; 
  signal DOUT_1_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_1_OBUF : STD_LOGIC; 
  signal DOUT_1_OD : STD_LOGIC; 
  signal DOUT_2_ENABLE : STD_LOGIC; 
  signal DOUT_2_TORGTS : STD_LOGIC; 
  signal DOUT_2_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_2_OBUF : STD_LOGIC; 
  signal DOUT_2_OD : STD_LOGIC; 
  signal DOUT_3_ENABLE : STD_LOGIC; 
  signal DOUT_3_TORGTS : STD_LOGIC; 
  signal DOUT_3_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_3_OBUF : STD_LOGIC; 
  signal DOUT_3_OD : STD_LOGIC; 
  signal DOUT_4_ENABLE : STD_LOGIC; 
  signal DOUT_4_TORGTS : STD_LOGIC; 
  signal DOUT_4_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_4_OBUF : STD_LOGIC; 
  signal DOUT_4_OD : STD_LOGIC; 
  signal DOUT_5_ENABLE : STD_LOGIC; 
  signal DOUT_5_TORGTS : STD_LOGIC; 
  signal DOUT_5_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_5_OBUF : STD_LOGIC; 
  signal DOUT_5_OD : STD_LOGIC; 
  signal DOUT_6_ENABLE : STD_LOGIC; 
  signal DOUT_6_TORGTS : STD_LOGIC; 
  signal DOUT_6_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_6_OBUF : STD_LOGIC; 
  signal DOUT_6_OD : STD_LOGIC; 
  signal DOUT_7_ENABLE : STD_LOGIC; 
  signal DOUT_7_TORGTS : STD_LOGIC; 
  signal DOUT_7_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_7_OBUF : STD_LOGIC; 
  signal DOUT_7_OD : STD_LOGIC; 
  signal DOUT_8_ENABLE : STD_LOGIC; 
  signal DOUT_8_TORGTS : STD_LOGIC; 
  signal DOUT_8_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_8_OBUF : STD_LOGIC; 
  signal DOUT_8_OD : STD_LOGIC; 
  signal DOUT_9_ENABLE : STD_LOGIC; 
  signal DOUT_9_TORGTS : STD_LOGIC; 
  signal DOUT_9_OUTMUX : STD_LOGIC; 
  signal rx_output_DOUT_9_OBUF : STD_LOGIC; 
  signal DOUT_9_OD : STD_LOGIC; 
  signal SOUT_ENABLE : STD_LOGIC; 
  signal SOUT_TORGTS : STD_LOGIC; 
  signal SOUT_OUTMUX : STD_LOGIC; 
  signal mac_control_SOUT_OBUF : STD_LOGIC; 
  signal SOUT_OCEMUXNOT : STD_LOGIC; 
  signal SOUT_OD : STD_LOGIC; 
  signal SCLK_ICEMUXNOT : STD_LOGIC; 
  signal SCLK_IDELAY : STD_LOGIC; 
  signal mac_control_SCLK_IBUF : STD_LOGIC; 
  signal LEDRX_ENABLE : STD_LOGIC; 
  signal LEDRX_TORGTS : STD_LOGIC; 
  signal LEDRX_OUTMUX : STD_LOGIC; 
  signal mac_control_LEDRX_OBUF : STD_LOGIC; 
  signal LEDRX_OCEMUXNOT : STD_LOGIC; 
  signal LEDRX_OD : STD_LOGIC; 
  signal LEDTX_ENABLE : STD_LOGIC; 
  signal LEDTX_TORGTS : STD_LOGIC; 
  signal LEDTX_OUTMUX : STD_LOGIC; 
  signal mac_control_LEDTX_OBUF : STD_LOGIC; 
  signal LEDTX_OCEMUXNOT : STD_LOGIC; 
  signal LEDTX_OD : STD_LOGIC; 
  signal tx_input_DIN_0_IBUF : STD_LOGIC; 
  signal tx_input_DIN_1_IBUF : STD_LOGIC; 
  signal tx_input_DIN_2_IBUF : STD_LOGIC; 
  signal tx_input_DIN_3_IBUF : STD_LOGIC; 
  signal tx_input_DIN_4_IBUF : STD_LOGIC; 
  signal tx_input_DIN_5_IBUF : STD_LOGIC; 
  signal tx_input_DIN_6_IBUF : STD_LOGIC; 
  signal tx_input_DIN_7_IBUF : STD_LOGIC; 
  signal tx_input_DIN_8_IBUF : STD_LOGIC; 
  signal tx_input_DIN_9_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RX_ER_IBUF : STD_LOGIC; 
  signal rx_input_GMII_RX_DV_IBUF : STD_LOGIC; 
  signal MA_10_ENABLE : STD_LOGIC; 
  signal MA_10_TORGTS : STD_LOGIC; 
  signal MA_10_OUTMUX : STD_LOGIC; 
  signal MA_10_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1530_FFX_RST : STD_LOGIC; 
  signal MA_11_ENABLE : STD_LOGIC; 
  signal MA_11_TORGTS : STD_LOGIC; 
  signal MA_11_OUTMUX : STD_LOGIC; 
  signal MA_11_OD : STD_LOGIC; 
  signal MA_12_ENABLE : STD_LOGIC; 
  signal MA_12_TORGTS : STD_LOGIC; 
  signal MA_12_OUTMUX : STD_LOGIC; 
  signal MA_12_OD : STD_LOGIC; 
  signal MA_13_ENABLE : STD_LOGIC; 
  signal MA_13_TORGTS : STD_LOGIC; 
  signal MA_13_OUTMUX : STD_LOGIC; 
  signal MA_13_OD : STD_LOGIC; 
  signal MA_14_ENABLE : STD_LOGIC; 
  signal MA_14_TORGTS : STD_LOGIC; 
  signal MA_14_OUTMUX : STD_LOGIC; 
  signal MA_14_OD : STD_LOGIC; 
  signal MA_15_ENABLE : STD_LOGIC; 
  signal MA_15_TORGTS : STD_LOGIC; 
  signal MA_15_OUTMUX : STD_LOGIC; 
  signal MA_15_OD : STD_LOGIC; 
  signal MA_16_ENABLE : STD_LOGIC; 
  signal MA_16_TORGTS : STD_LOGIC; 
  signal MA_16_OUTMUX : STD_LOGIC; 
  signal MA_16_OD : STD_LOGIC; 
  signal MD_10_ENABLE : STD_LOGIC; 
  signal MD_10_TORGTS : STD_LOGIC; 
  signal MD_10_OUTMUX : STD_LOGIC; 
  signal MD_10_OD : STD_LOGIC; 
  signal MD_11_ENABLE : STD_LOGIC; 
  signal MD_11_TORGTS : STD_LOGIC; 
  signal MD_11_OUTMUX : STD_LOGIC; 
  signal MD_11_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1599_FFY_SET : STD_LOGIC; 
  signal MD_20_ENABLE : STD_LOGIC; 
  signal MD_20_TORGTS : STD_LOGIC; 
  signal MD_20_OUTMUX : STD_LOGIC; 
  signal MD_20_OD : STD_LOGIC; 
  signal MD_12_ENABLE : STD_LOGIC; 
  signal MD_12_TORGTS : STD_LOGIC; 
  signal MD_12_OUTMUX : STD_LOGIC; 
  signal MD_12_OD : STD_LOGIC; 
  signal MD_21_ENABLE : STD_LOGIC; 
  signal MD_21_TORGTS : STD_LOGIC; 
  signal MD_21_OUTMUX : STD_LOGIC; 
  signal MD_21_OD : STD_LOGIC; 
  signal MD_13_ENABLE : STD_LOGIC; 
  signal MD_13_TORGTS : STD_LOGIC; 
  signal MD_13_OUTMUX : STD_LOGIC; 
  signal MD_13_OD : STD_LOGIC; 
  signal MD_22_ENABLE : STD_LOGIC; 
  signal MD_22_TORGTS : STD_LOGIC; 
  signal MD_22_OUTMUX : STD_LOGIC; 
  signal MD_22_OD : STD_LOGIC; 
  signal MD_14_ENABLE : STD_LOGIC; 
  signal MD_14_TORGTS : STD_LOGIC; 
  signal MD_14_OUTMUX : STD_LOGIC; 
  signal MD_14_OD : STD_LOGIC; 
  signal MD_30_ENABLE : STD_LOGIC; 
  signal MD_30_TORGTS : STD_LOGIC; 
  signal MD_30_OUTMUX : STD_LOGIC; 
  signal MD_30_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15_FFY_RST : STD_LOGIC; 
  signal MD_23_ENABLE : STD_LOGIC; 
  signal MD_23_TORGTS : STD_LOGIC; 
  signal MD_23_OUTMUX : STD_LOGIC; 
  signal MD_23_OD : STD_LOGIC; 
  signal MD_15_ENABLE : STD_LOGIC; 
  signal MD_15_TORGTS : STD_LOGIC; 
  signal MD_15_OUTMUX : STD_LOGIC; 
  signal MD_15_OD : STD_LOGIC; 
  signal MD_31_ENABLE : STD_LOGIC; 
  signal MD_31_TORGTS : STD_LOGIC; 
  signal MD_31_OUTMUX : STD_LOGIC; 
  signal MD_31_OD : STD_LOGIC; 
  signal MD_24_ENABLE : STD_LOGIC; 
  signal MD_24_TORGTS : STD_LOGIC; 
  signal MD_24_OUTMUX : STD_LOGIC; 
  signal MD_24_OD : STD_LOGIC; 
  signal MD_16_ENABLE : STD_LOGIC; 
  signal MD_16_TORGTS : STD_LOGIC; 
  signal MD_16_OUTMUX : STD_LOGIC; 
  signal MD_16_OD : STD_LOGIC; 
  signal MD_17_ENABLE : STD_LOGIC; 
  signal MD_17_TORGTS : STD_LOGIC; 
  signal MD_17_OUTMUX : STD_LOGIC; 
  signal MD_17_OD : STD_LOGIC; 
  signal MD_25_ENABLE : STD_LOGIC; 
  signal MD_25_TORGTS : STD_LOGIC; 
  signal MD_25_OUTMUX : STD_LOGIC; 
  signal MD_25_OD : STD_LOGIC; 
  signal MD_18_ENABLE : STD_LOGIC; 
  signal MD_18_TORGTS : STD_LOGIC; 
  signal MD_18_OUTMUX : STD_LOGIC; 
  signal MD_18_OD : STD_LOGIC; 
  signal MD_26_ENABLE : STD_LOGIC; 
  signal MD_26_TORGTS : STD_LOGIC; 
  signal MD_26_OUTMUX : STD_LOGIC; 
  signal MD_26_OD : STD_LOGIC; 
  signal MD_19_ENABLE : STD_LOGIC; 
  signal MD_19_TORGTS : STD_LOGIC; 
  signal MD_19_OUTMUX : STD_LOGIC; 
  signal MD_19_OD : STD_LOGIC; 
  signal MD_27_ENABLE : STD_LOGIC; 
  signal MD_27_TORGTS : STD_LOGIC; 
  signal MD_27_OUTMUX : STD_LOGIC; 
  signal MD_27_OD : STD_LOGIC; 
  signal MD_28_ENABLE : STD_LOGIC; 
  signal MD_28_TORGTS : STD_LOGIC; 
  signal MD_28_OUTMUX : STD_LOGIC; 
  signal MD_28_OD : STD_LOGIC; 
  signal MD_29_ENABLE : STD_LOGIC; 
  signal MD_29_TORGTS : STD_LOGIC; 
  signal MD_29_OUTMUX : STD_LOGIC; 
  signal MD_29_OD : STD_LOGIC; 
  signal MA_0_ENABLE : STD_LOGIC; 
  signal MA_0_TORGTS : STD_LOGIC; 
  signal MA_0_OUTMUX : STD_LOGIC; 
  signal MA_0_OD : STD_LOGIC; 
  signal MA_1_ENABLE : STD_LOGIC; 
  signal MA_1_TORGTS : STD_LOGIC; 
  signal MA_1_OUTMUX : STD_LOGIC; 
  signal MA_1_OD : STD_LOGIC; 
  signal MA_2_ENABLE : STD_LOGIC; 
  signal MA_2_TORGTS : STD_LOGIC; 
  signal MA_2_OUTMUX : STD_LOGIC; 
  signal MA_2_OD : STD_LOGIC; 
  signal MA_3_ENABLE : STD_LOGIC; 
  signal MA_3_TORGTS : STD_LOGIC; 
  signal MA_3_OUTMUX : STD_LOGIC; 
  signal MA_3_OD : STD_LOGIC; 
  signal MA_4_ENABLE : STD_LOGIC; 
  signal MA_4_TORGTS : STD_LOGIC; 
  signal MA_4_OUTMUX : STD_LOGIC; 
  signal MA_4_OD : STD_LOGIC; 
  signal MA_5_ENABLE : STD_LOGIC; 
  signal MA_5_TORGTS : STD_LOGIC; 
  signal MA_5_OUTMUX : STD_LOGIC; 
  signal MA_5_OD : STD_LOGIC; 
  signal MA_6_ENABLE : STD_LOGIC; 
  signal MA_6_TORGTS : STD_LOGIC; 
  signal MA_6_OUTMUX : STD_LOGIC; 
  signal MA_6_OD : STD_LOGIC; 
  signal MA_7_ENABLE : STD_LOGIC; 
  signal MA_7_TORGTS : STD_LOGIC; 
  signal MA_7_OUTMUX : STD_LOGIC; 
  signal MA_7_OD : STD_LOGIC; 
  signal MA_8_ENABLE : STD_LOGIC; 
  signal MA_8_TORGTS : STD_LOGIC; 
  signal MA_8_OUTMUX : STD_LOGIC; 
  signal MA_8_OD : STD_LOGIC; 
  signal mac_control_phyaddr_9_FFY_RST : STD_LOGIC; 
  signal MA_9_ENABLE : STD_LOGIC; 
  signal MA_9_TORGTS : STD_LOGIC; 
  signal MA_9_OUTMUX : STD_LOGIC; 
  signal MA_9_OD : STD_LOGIC; 
  signal PHYRESET_ENABLE : STD_LOGIC; 
  signal PHYRESET_TORGTS : STD_LOGIC; 
  signal PHYRESET_OUTMUX : STD_LOGIC; 
  signal mac_control_PHYRESET_OBUF : STD_LOGIC; 
  signal PHYRESET_OD : STD_LOGIC; 
  signal MD_0_ENABLE : STD_LOGIC; 
  signal MD_0_TORGTS : STD_LOGIC; 
  signal MD_0_OUTMUX : STD_LOGIC; 
  signal MD_0_OD : STD_LOGIC; 
  signal MD_1_ENABLE : STD_LOGIC; 
  signal MD_1_TORGTS : STD_LOGIC; 
  signal MD_1_OUTMUX : STD_LOGIC; 
  signal MD_1_OD : STD_LOGIC; 
  signal rx_input_fifo_fifo_N15_FFX_RST : STD_LOGIC; 
  signal MD_2_ENABLE : STD_LOGIC; 
  signal MD_2_TORGTS : STD_LOGIC; 
  signal MD_2_OUTMUX : STD_LOGIC; 
  signal MD_2_OD : STD_LOGIC; 
  signal MD_3_ENABLE : STD_LOGIC; 
  signal MD_3_TORGTS : STD_LOGIC; 
  signal MD_3_OUTMUX : STD_LOGIC; 
  signal MD_3_OD : STD_LOGIC; 
  signal MD_4_ENABLE : STD_LOGIC; 
  signal MD_4_TORGTS : STD_LOGIC; 
  signal MD_4_OUTMUX : STD_LOGIC; 
  signal MD_4_OD : STD_LOGIC; 
  signal MD_5_ENABLE : STD_LOGIC; 
  signal MD_5_TORGTS : STD_LOGIC; 
  signal MD_5_OUTMUX : STD_LOGIC; 
  signal MD_5_OD : STD_LOGIC; 
  signal MD_6_ENABLE : STD_LOGIC; 
  signal MD_6_TORGTS : STD_LOGIC; 
  signal MD_6_OUTMUX : STD_LOGIC; 
  signal MD_6_OD : STD_LOGIC; 
  signal MD_7_ENABLE : STD_LOGIC; 
  signal MD_7_TORGTS : STD_LOGIC; 
  signal MD_7_OUTMUX : STD_LOGIC; 
  signal MD_7_OD : STD_LOGIC; 
  signal MD_8_ENABLE : STD_LOGIC; 
  signal MD_8_TORGTS : STD_LOGIC; 
  signal MD_8_OUTMUX : STD_LOGIC; 
  signal MD_8_OD : STD_LOGIC; 
  signal MD_9_ENABLE : STD_LOGIC; 
  signal MD_9_TORGTS : STD_LOGIC; 
  signal MD_9_OUTMUX : STD_LOGIC; 
  signal MD_9_OD : STD_LOGIC; 
  signal GTX_CLK_ENABLE : STD_LOGIC; 
  signal GTX_CLK_TORGTS : STD_LOGIC; 
  signal GTX_CLK_OUTMUX : STD_LOGIC; 
  signal clkio_dll_LOCKED : STD_LOGIC; 
  signal clkio_dll_CLKDV : STD_LOGIC; 
  signal clkio_dll_CLK2X180 : STD_LOGIC; 
  signal clkio_dll_CLK2X : STD_LOGIC; 
  signal clkio_dll_CLK270 : STD_LOGIC; 
  signal clkio_dll_CLK180 : STD_LOGIC; 
  signal clkio_dll_CLK90 : STD_LOGIC; 
  signal clk_dll_LOCKED : STD_LOGIC; 
  signal clk_dll_CLK2X180 : STD_LOGIC; 
  signal clk_dll_CLK2X : STD_LOGIC; 
  signal clk_dll_CLK270 : STD_LOGIC; 
  signal clk_dll_CLK180 : STD_LOGIC; 
  signal clk_dll_CLK90 : STD_LOGIC; 
  signal clkrx_dll_LOCKED : STD_LOGIC; 
  signal clkrx_dll_CLKDV : STD_LOGIC; 
  signal clkrx_dll_CLK2X180 : STD_LOGIC; 
  signal clkrx_dll_CLK2X : STD_LOGIC; 
  signal clkrx_dll_CLK270 : STD_LOGIC; 
  signal clkrx_dll_CLK180 : STD_LOGIC; 
  signal clkrx_dll_CLK90 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOB9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA15 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA14 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA13 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA12 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA11 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA10 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA9 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA8 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA7 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA6 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA5 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA4 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA3 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA2 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_DOA0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRB3 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRB2 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRB1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRB0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRA3 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRA2 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRA1 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_ADDRA0 : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_fifo_B7_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA15 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA14 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA13 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA12 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA11 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA10 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA9 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA8 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA7 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA6 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA5 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA4 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA3 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA2 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA1 : STD_LOGIC; 
  signal rx_output_fifo_B7_DOA0 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRB3 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRB2 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRB1 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRB0 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRA3 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRA2 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRA1 : STD_LOGIC; 
  signal rx_output_fifo_B7_ADDRA0 : STD_LOGIC; 
  signal rx_output_fifo_B7_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_B7_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_N81880 : STD_LOGIC; 
  signal mac_control_dout_19_rt : STD_LOGIC; 
  signal mac_control_N81872 : STD_LOGIC; 
  signal mac_control_dout_20_rt : STD_LOGIC; 
  signal mac_control_N81896 : STD_LOGIC; 
  signal mac_control_dout_21_rt : STD_LOGIC; 
  signal mac_control_N81884 : STD_LOGIC; 
  signal mac_control_dout_29_rt : STD_LOGIC; 
  signal mac_control_N81856 : STD_LOGIC; 
  signal mac_control_dout_22_rt : STD_LOGIC; 
  signal mac_control_N81900 : STD_LOGIC; 
  signal mac_control_dout_15_rt : STD_LOGIC; 
  signal rx_input_fifo_fifo_N1599_FFX_RST : STD_LOGIC; 
  signal mac_control_N81852 : STD_LOGIC; 
  signal mac_control_dout_23_rt : STD_LOGIC; 
  signal mac_control_N81876 : STD_LOGIC; 
  signal mac_control_dout_24_rt : STD_LOGIC; 
  signal mac_control_N81904 : STD_LOGIC; 
  signal mac_control_dout_16_rt : STD_LOGIC; 
  signal mac_control_N81908 : STD_LOGIC; 
  signal mac_control_dout_25_rt : STD_LOGIC; 
  signal mac_control_N81868 : STD_LOGIC; 
  signal mac_control_dout_17_rt : STD_LOGIC; 
  signal mac_control_N81892 : STD_LOGIC; 
  signal mac_control_dout_18_rt : STD_LOGIC; 
  signal mac_control_N81860 : STD_LOGIC; 
  signal mac_control_dout_26_rt : STD_LOGIC; 
  signal mac_control_N81888 : STD_LOGIC; 
  signal mac_control_dout_27_rt : STD_LOGIC; 
  signal mac_control_N81864 : STD_LOGIC; 
  signal mac_control_dout_28_rt : STD_LOGIC; 
  signal mac_control_phyaddr_9_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81848 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81846 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE977_F5MUX : STD_LOGIC; 
  signal memcontroller_N81728 : STD_LOGIC; 
  signal memcontroller_N81726 : STD_LOGIC; 
  signal memcontroller_addrn_0_F5MUX : STD_LOGIC; 
  signal memcontroller_N81688 : STD_LOGIC; 
  signal memcontroller_N81686 : STD_LOGIC; 
  signal memcontroller_addrn_8_F5MUX : STD_LOGIC; 
  signal memcontroller_N81723 : STD_LOGIC; 
  signal memcontroller_N81721 : STD_LOGIC; 
  signal memcontroller_addrn_1_F5MUX : STD_LOGIC; 
  signal memcontroller_N81683 : STD_LOGIC; 
  signal memcontroller_N81681 : STD_LOGIC; 
  signal memcontroller_addrn_9_F5MUX : STD_LOGIC; 
  signal memcontroller_N81718 : STD_LOGIC; 
  signal memcontroller_N81716 : STD_LOGIC; 
  signal memcontroller_addrn_2_F5MUX : STD_LOGIC; 
  signal memcontroller_N81678 : STD_LOGIC; 
  signal memcontroller_N81676 : STD_LOGIC; 
  signal memcontroller_addrn_10_F5MUX : STD_LOGIC; 
  signal memcontroller_N81713 : STD_LOGIC; 
  signal memcontroller_N81711 : STD_LOGIC; 
  signal memcontroller_addrn_3_F5MUX : STD_LOGIC; 
  signal memcontroller_N81673 : STD_LOGIC; 
  signal memcontroller_N81671 : STD_LOGIC; 
  signal memcontroller_addrn_11_F5MUX : STD_LOGIC; 
  signal memcontroller_N81708 : STD_LOGIC; 
  signal memcontroller_N81706 : STD_LOGIC; 
  signal memcontroller_addrn_4_F5MUX : STD_LOGIC; 
  signal memcontroller_N81668 : STD_LOGIC; 
  signal memcontroller_N81666 : STD_LOGIC; 
  signal memcontroller_addrn_12_F5MUX : STD_LOGIC; 
  signal memcontroller_N81703 : STD_LOGIC; 
  signal memcontroller_N81701 : STD_LOGIC; 
  signal memcontroller_addrn_5_F5MUX : STD_LOGIC; 
  signal memcontroller_N81608 : STD_LOGIC; 
  signal memcontroller_N81606 : STD_LOGIC; 
  signal memcontroller_addrn_13_F5MUX : STD_LOGIC; 
  signal memcontroller_N81698 : STD_LOGIC; 
  signal memcontroller_N81696 : STD_LOGIC; 
  signal memcontroller_addrn_6_F5MUX : STD_LOGIC; 
  signal memcontroller_N81603 : STD_LOGIC; 
  signal memcontroller_N81601 : STD_LOGIC; 
  signal memcontroller_addrn_14_F5MUX : STD_LOGIC; 
  signal memcontroller_N81693 : STD_LOGIC; 
  signal memcontroller_N81691 : STD_LOGIC; 
  signal memcontroller_addrn_7_F5MUX : STD_LOGIC; 
  signal memcontroller_N81613 : STD_LOGIC; 
  signal memcontroller_N81611 : STD_LOGIC; 
  signal memcontroller_addrn_15_F5MUX : STD_LOGIC; 
  signal memcontroller_addrn_16_FROM : STD_LOGIC; 
  signal memcontroller_addrn_16_GROM : STD_LOGIC; 
  signal memcontroller_addrn_16_F5MUX : STD_LOGIC; 
  signal memcontroller_N81828 : STD_LOGIC; 
  signal memcontroller_N81826 : STD_LOGIC; 
  signal memcontroller_dnl1_10_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81783 : STD_LOGIC; 
  signal memcontroller_N81781 : STD_LOGIC; 
  signal memcontroller_dnl1_1_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81833 : STD_LOGIC; 
  signal memcontroller_N81831 : STD_LOGIC; 
  signal memcontroller_dnl1_11_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81778 : STD_LOGIC; 
  signal memcontroller_N81776 : STD_LOGIC; 
  signal memcontroller_dnl1_0_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_validucast_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0052 : STD_LOGIC; 
  signal rx_input_memio_addrchk_validucast_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpen_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_destok_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0053 : STD_LOGIC; 
  signal rx_input_memio_destok_CEMUXNOT : STD_LOGIC; 
  signal rx_output_cs_FFd10_FROM : STD_LOGIC; 
  signal rx_output_cs_FFd10_In : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_26_Xo_1_GROM : STD_LOGIC; 
  signal tx_output_crcl_18_FROM : STD_LOGIC; 
  signal tx_output_n0034_18_Q : STD_LOGIC; 
  signal tx_output_crcl_26_FROM : STD_LOGIC; 
  signal tx_output_n0034_26_Q : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_19_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_19_Q : STD_LOGIC; 
  signal rx_input_memio_crcl_13_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_13_Q : STD_LOGIC; 
  signal tx_output_crcl_27_FROM : STD_LOGIC; 
  signal tx_output_n0034_27_Q : STD_LOGIC; 
  signal rx_output_cs_FFd6_FROM : STD_LOGIC; 
  signal rx_output_cs_FFd6_In : STD_LOGIC; 
  signal rx_input_memio_crcl_30_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_30_1_O : STD_LOGIC; 
  signal rx_input_memio_crcl_14_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_14_Q : STD_LOGIC; 
  signal tx_input_cs_FFd12_FROM : STD_LOGIC; 
  signal tx_input_cs_FFd12_In : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_5_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_9_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_11_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_21_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_13_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_13_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_31_CEMUXNOT : STD_LOGIC; 
  signal tx_input_fifofulll_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_23_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_15_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_41_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_33_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_33_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_25_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_17_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_43_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_43_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81838 : STD_LOGIC; 
  signal memcontroller_N81836 : STD_LOGIC; 
  signal memcontroller_dnl1_12_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81653 : STD_LOGIC; 
  signal memcontroller_N81651 : STD_LOGIC; 
  signal memcontroller_dnl1_20_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81788 : STD_LOGIC; 
  signal memcontroller_N81786 : STD_LOGIC; 
  signal memcontroller_dnl1_2_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81658 : STD_LOGIC; 
  signal memcontroller_N81656 : STD_LOGIC; 
  signal memcontroller_dnl1_21_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81843 : STD_LOGIC; 
  signal memcontroller_N81841 : STD_LOGIC; 
  signal memcontroller_dnl1_13_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81738 : STD_LOGIC; 
  signal memcontroller_N81736 : STD_LOGIC; 
  signal memcontroller_dnl1_30_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81663 : STD_LOGIC; 
  signal memcontroller_N81661 : STD_LOGIC; 
  signal memcontroller_dnl1_22_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_dout_1_FFY_RST : STD_LOGIC; 
  signal memcontroller_N81623 : STD_LOGIC; 
  signal memcontroller_N81621 : STD_LOGIC; 
  signal memcontroller_dnl1_14_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81773 : STD_LOGIC; 
  signal memcontroller_N81771 : STD_LOGIC; 
  signal memcontroller_dnl1_31_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81628 : STD_LOGIC; 
  signal memcontroller_N81626 : STD_LOGIC; 
  signal memcontroller_dnl1_15_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81618 : STD_LOGIC; 
  signal memcontroller_N81616 : STD_LOGIC; 
  signal memcontroller_dnl1_23_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81793 : STD_LOGIC; 
  signal memcontroller_N81791 : STD_LOGIC; 
  signal memcontroller_dnl1_3_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81798 : STD_LOGIC; 
  signal memcontroller_N81796 : STD_LOGIC; 
  signal memcontroller_dnl1_4_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81768 : STD_LOGIC; 
  signal memcontroller_N81766 : STD_LOGIC; 
  signal memcontroller_dnl1_24_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81633 : STD_LOGIC; 
  signal memcontroller_N81631 : STD_LOGIC; 
  signal memcontroller_dnl1_16_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81803 : STD_LOGIC; 
  signal memcontroller_N81801 : STD_LOGIC; 
  signal memcontroller_dnl1_5_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81763 : STD_LOGIC; 
  signal memcontroller_N81761 : STD_LOGIC; 
  signal memcontroller_dnl1_25_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81638 : STD_LOGIC; 
  signal memcontroller_N81636 : STD_LOGIC; 
  signal memcontroller_dnl1_17_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_11_FFY_RST : STD_LOGIC; 
  signal memcontroller_N81808 : STD_LOGIC; 
  signal memcontroller_N81806 : STD_LOGIC; 
  signal memcontroller_dnl1_6_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81758 : STD_LOGIC; 
  signal memcontroller_N81756 : STD_LOGIC; 
  signal memcontroller_dnl1_26_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_dout_1_FFX_RST : STD_LOGIC; 
  signal memcontroller_N81643 : STD_LOGIC; 
  signal memcontroller_N81641 : STD_LOGIC; 
  signal memcontroller_dnl1_18_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81813 : STD_LOGIC; 
  signal memcontroller_N81811 : STD_LOGIC; 
  signal memcontroller_dnl1_7_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81753 : STD_LOGIC; 
  signal memcontroller_N81751 : STD_LOGIC; 
  signal memcontroller_dnl1_27_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81648 : STD_LOGIC; 
  signal memcontroller_N81646 : STD_LOGIC; 
  signal memcontroller_dnl1_19_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81818 : STD_LOGIC; 
  signal memcontroller_N81816 : STD_LOGIC; 
  signal memcontroller_dnl1_8_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81748 : STD_LOGIC; 
  signal memcontroller_N81746 : STD_LOGIC; 
  signal memcontroller_dnl1_28_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81823 : STD_LOGIC; 
  signal memcontroller_N81821 : STD_LOGIC; 
  signal memcontroller_dnl1_9_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_N81743 : STD_LOGIC; 
  signal memcontroller_N81741 : STD_LOGIC; 
  signal memcontroller_dnl1_29_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0076_inst_lut2_127 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_1_CYMUXG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_1_XORG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_1_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_181 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_1_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_2_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_2_XORF : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_2_CYMUXG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_2_XORG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_2_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_183 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_2_CYINIT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_4_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_4_XORF : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_4_XORG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_5_rt : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_185 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_n0076_4_CYINIT : STD_LOGIC; 
  signal txfbbp_11_FFX_RST : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_lut2_0 : STD_LOGIC; 
  signal addr2ext_0_CYMUXG : STD_LOGIC; 
  signal addr2ext_0_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_0 : STD_LOGIC; 
  signal addr2ext_0_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_2_FROM : STD_LOGIC; 
  signal addr2ext_2_CYMUXG : STD_LOGIC; 
  signal addr2ext_2_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_2_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_2 : STD_LOGIC; 
  signal addr2ext_2_CYINIT : STD_LOGIC; 
  signal addr2ext_4_FROM : STD_LOGIC; 
  signal addr2ext_4_CYMUXG : STD_LOGIC; 
  signal addr2ext_4_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_4_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_4 : STD_LOGIC; 
  signal addr2ext_4_CYINIT : STD_LOGIC; 
  signal addr2ext_6_FROM : STD_LOGIC; 
  signal addr2ext_6_CYMUXG : STD_LOGIC; 
  signal addr2ext_6_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_6_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_6 : STD_LOGIC; 
  signal addr2ext_6_CYINIT : STD_LOGIC; 
  signal addr2ext_8_FROM : STD_LOGIC; 
  signal addr2ext_8_CYMUXG : STD_LOGIC; 
  signal addr2ext_8_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_8_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_8 : STD_LOGIC; 
  signal addr2ext_8_CYINIT : STD_LOGIC; 
  signal addr2ext_10_FROM : STD_LOGIC; 
  signal addr2ext_10_CYMUXG : STD_LOGIC; 
  signal addr2ext_10_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_10_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_10 : STD_LOGIC; 
  signal addr2ext_10_CYINIT : STD_LOGIC; 
  signal addr2ext_12_FROM : STD_LOGIC; 
  signal addr2ext_12_CYMUXG : STD_LOGIC; 
  signal addr2ext_12_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_12_GROM : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_12 : STD_LOGIC; 
  signal addr2ext_12_CYINIT : STD_LOGIC; 
  signal addr2ext_14_LOGIC_ZERO : STD_LOGIC; 
  signal addr2ext_14_FROM : STD_LOGIC; 
  signal addr2ext_15_rt : STD_LOGIC; 
  signal tx_output_addr_Madd_n0000_inst_cy_14 : STD_LOGIC; 
  signal addr2ext_14_CYINIT : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_2_rt : STD_LOGIC; 
  signal rx_input_memio_bcnt_86_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_72 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_270 : STD_LOGIC; 
  signal rx_input_memio_bcnt_86_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_235 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_73 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_236 : STD_LOGIC; 
  signal rx_input_memio_bcnt_87_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_87_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_87_XORG : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_74 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_272 : STD_LOGIC; 
  signal rx_input_memio_bcnt_87_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_75 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_238 : STD_LOGIC; 
  signal rx_input_memio_bcnt_89_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_89_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_76 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_274 : STD_LOGIC; 
  signal rx_input_memio_bcnt_89_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_239 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_77 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_240 : STD_LOGIC; 
  signal rx_input_memio_bcnt_91_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_91_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_78 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_276 : STD_LOGIC; 
  signal rx_input_memio_bcnt_91_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_241 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_79 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_242 : STD_LOGIC; 
  signal rx_input_memio_bcnt_93_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_93_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_80 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_278 : STD_LOGIC; 
  signal rx_input_memio_bcnt_93_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_243 : STD_LOGIC; 
  signal rx_input_memio_dout_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_81 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_244 : STD_LOGIC; 
  signal rx_input_memio_bcnt_95_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_95_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_82 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_280 : STD_LOGIC; 
  signal rx_input_memio_bcnt_95_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_245 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_83 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_246 : STD_LOGIC; 
  signal rx_input_memio_bcnt_97_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_97_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_84 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_282 : STD_LOGIC; 
  signal rx_input_memio_bcnt_97_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_247 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_85 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_248 : STD_LOGIC; 
  signal rx_input_memio_bcnt_99_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_bcnt_99_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_86 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_cy_284 : STD_LOGIC; 
  signal rx_input_memio_bcnt_99_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_249 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_lut3_87 : STD_LOGIC; 
  signal rx_input_memio_bcnt_inst_sum_250 : STD_LOGIC; 
  signal rx_input_memio_bcnt_101_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_lut2_4811_O : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_49_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_lut2_491_O : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_48 : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_49_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_2_FROM : STD_LOGIC; 
  signal rx_output_n0060_2_XORF : STD_LOGIC; 
  signal rx_output_n0060_2_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_2_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_2_XORG : STD_LOGIC; 
  signal rx_output_n0060_2_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_50 : STD_LOGIC; 
  signal rx_output_n0060_2_CYINIT : STD_LOGIC; 
  signal rx_output_n0060_4_FROM : STD_LOGIC; 
  signal rx_output_n0060_4_XORF : STD_LOGIC; 
  signal rx_output_n0060_4_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_4_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_4_XORG : STD_LOGIC; 
  signal rx_output_n0060_4_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_52 : STD_LOGIC; 
  signal rx_output_n0060_4_CYINIT : STD_LOGIC; 
  signal rx_input_memio_dout_5_FFY_RST : STD_LOGIC; 
  signal rx_output_n0060_6_FROM : STD_LOGIC; 
  signal rx_output_n0060_6_XORF : STD_LOGIC; 
  signal rx_output_n0060_6_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_6_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_6_XORG : STD_LOGIC; 
  signal rx_output_n0060_6_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_54 : STD_LOGIC; 
  signal rx_output_n0060_6_CYINIT : STD_LOGIC; 
  signal rx_output_n0060_8_FROM : STD_LOGIC; 
  signal rx_output_n0060_8_XORF : STD_LOGIC; 
  signal rx_output_n0060_8_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_8_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_8_XORG : STD_LOGIC; 
  signal rx_output_n0060_8_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_56 : STD_LOGIC; 
  signal rx_output_n0060_8_CYINIT : STD_LOGIC; 
  signal rx_output_n0060_10_FROM : STD_LOGIC; 
  signal rx_output_n0060_10_XORF : STD_LOGIC; 
  signal rx_output_n0060_10_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_10_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_10_XORG : STD_LOGIC; 
  signal rx_output_n0060_10_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_58 : STD_LOGIC; 
  signal rx_output_n0060_10_CYINIT : STD_LOGIC; 
  signal rx_output_n0060_12_FROM : STD_LOGIC; 
  signal rx_output_n0060_12_XORF : STD_LOGIC; 
  signal rx_output_n0060_12_CYMUXG : STD_LOGIC; 
  signal rx_output_n0060_12_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_12_XORG : STD_LOGIC; 
  signal rx_output_n0060_12_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_60 : STD_LOGIC; 
  signal rx_output_n0060_12_CYINIT : STD_LOGIC; 
  signal txfbbp_13_FFX_RST : STD_LOGIC; 
  signal rx_output_n0060_14_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0060_14_FROM : STD_LOGIC; 
  signal rx_output_n0060_14_XORF : STD_LOGIC; 
  signal rx_output_n0060_14_XORG : STD_LOGIC; 
  signal rx_output_len_15_rt : STD_LOGIC; 
  signal rx_output_Madd_n0060_inst_cy_62 : STD_LOGIC; 
  signal rx_output_n0060_14_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_4_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0036_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_4_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_18_CYINIT : STD_LOGIC; 
  signal rx_input_memio_dout_5_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_31_rt : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_rxcrcerr_cnt_30_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_0_FROM : STD_LOGIC; 
  signal rx_input_memio_bp_0_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_134 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_221 : STD_LOGIC; 
  signal rx_input_memio_bp_0_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_0_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_bp_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_135 : STD_LOGIC; 
  signal rx_input_memio_bp_2_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_136 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_223 : STD_LOGIC; 
  signal rx_input_memio_bp_2_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_137 : STD_LOGIC; 
  signal rx_input_memio_bp_4_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_138 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_225 : STD_LOGIC; 
  signal rx_input_memio_bp_4_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_6_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_139 : STD_LOGIC; 
  signal rx_input_memio_bp_6_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_140 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_227 : STD_LOGIC; 
  signal rx_input_memio_bp_6_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_8_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_141 : STD_LOGIC; 
  signal rx_input_memio_bp_8_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_142 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_229 : STD_LOGIC; 
  signal rx_input_memio_bp_8_CYINIT : STD_LOGIC; 
  signal txfbbp_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_10_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_143 : STD_LOGIC; 
  signal rx_input_memio_bp_10_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_144 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_231 : STD_LOGIC; 
  signal rx_input_memio_bp_10_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_12_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_145 : STD_LOGIC; 
  signal rx_input_memio_bp_12_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_146 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_233 : STD_LOGIC; 
  signal rx_input_memio_bp_12_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bp_14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_147 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_lut2_148 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0043_inst_cy_235 : STD_LOGIC; 
  signal rx_input_memio_bp_14_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_14_CYINIT : STD_LOGIC; 
  signal rx_input_memio_dout_9_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_16_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_7 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_102 : STD_LOGIC; 
  signal addr3ext_7_CYMUXG : STD_LOGIC; 
  signal addr3ext_7_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_8 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_109 : STD_LOGIC; 
  signal addr3ext_7_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_103 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_9 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_104 : STD_LOGIC; 
  signal addr3ext_9_CYMUXG : STD_LOGIC; 
  signal addr3ext_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_10 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_111 : STD_LOGIC; 
  signal addr3ext_9_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_105 : STD_LOGIC; 
  signal rx_input_data_5_FFY_RST : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_11 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_106 : STD_LOGIC; 
  signal addr3ext_11_CYMUXG : STD_LOGIC; 
  signal addr3ext_11_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_12 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_113 : STD_LOGIC; 
  signal addr3ext_11_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_107 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_13 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_108 : STD_LOGIC; 
  signal addr3ext_13_CYMUXG : STD_LOGIC; 
  signal addr3ext_13_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_14 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_115 : STD_LOGIC; 
  signal addr3ext_13_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_109 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_15 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_110 : STD_LOGIC; 
  signal addr3ext_15_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_diff_0_rt : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_SIG_21 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_151 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut4_8 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut4_9 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_153 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT : STD_LOGIC; 
  signal tx_output_cs_FFd4_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut4_10 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut4_11 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_155 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_diff_13_rt : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_SIG_22 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_157 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut3_32 : STD_LOGIC; 
  signal rx_fifocheck_n0003_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_lut3_33 : STD_LOGIC; 
  signal rx_fifocheck_Mcompar_n0003_inst_cy_159 : STD_LOGIC; 
  signal rx_fifocheck_n0003_LOGIC_ONE : STD_LOGIC; 
  signal rx_fifocheck_n0003_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_0_rt : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_SIG_23 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_151 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut4_8 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut4_9 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_153 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut4_10 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut4_11 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_155 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_13_rt : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_SIG_24 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_157 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut3_32 : STD_LOGIC; 
  signal tx_fifocheck_n0003_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_lut3_33 : STD_LOGIC; 
  signal tx_fifocheck_Mcompar_n0003_inst_cy_159 : STD_LOGIC; 
  signal tx_fifocheck_n0003_LOGIC_ONE : STD_LOGIC; 
  signal tx_fifocheck_n0003_CYINIT : STD_LOGIC; 
  signal mac_control_N53144_rt : STD_LOGIC; 
  signal mac_control_phyrstcnt_110_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_192 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_294 : STD_LOGIC; 
  signal mac_control_phyrstcnt_110_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_257 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_193 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_258 : STD_LOGIC; 
  signal mac_control_phyrstcnt_111_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_111_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_194 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_296 : STD_LOGIC; 
  signal mac_control_phyrstcnt_111_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_259 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_195 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_260 : STD_LOGIC; 
  signal mac_control_phyrstcnt_113_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_113_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_196 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_298 : STD_LOGIC; 
  signal mac_control_phyrstcnt_113_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_261 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_197 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_262 : STD_LOGIC; 
  signal mac_control_phyrstcnt_115_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_115_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_198 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_300 : STD_LOGIC; 
  signal mac_control_phyrstcnt_115_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_263 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_199 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_264 : STD_LOGIC; 
  signal mac_control_phyrstcnt_117_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_117_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_200 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_302 : STD_LOGIC; 
  signal mac_control_phyrstcnt_117_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_265 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_201 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_266 : STD_LOGIC; 
  signal mac_control_phyrstcnt_119_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_119_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_202 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_304 : STD_LOGIC; 
  signal mac_control_phyrstcnt_119_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_267 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_203 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_268 : STD_LOGIC; 
  signal mac_control_phyrstcnt_121_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_121_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_204 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_306 : STD_LOGIC; 
  signal mac_control_phyrstcnt_121_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_269 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_205 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_270 : STD_LOGIC; 
  signal mac_control_phyrstcnt_123_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_123_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_206 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_308 : STD_LOGIC; 
  signal mac_control_phyrstcnt_123_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_271 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_207 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_272 : STD_LOGIC; 
  signal mac_control_phyrstcnt_125_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_125_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_208 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_310 : STD_LOGIC; 
  signal mac_control_phyrstcnt_125_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_273 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_209 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_274 : STD_LOGIC; 
  signal mac_control_phyrstcnt_127_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_127_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_210 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_312 : STD_LOGIC; 
  signal mac_control_phyrstcnt_127_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_275 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_211 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_276 : STD_LOGIC; 
  signal mac_control_phyrstcnt_129_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_129_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_212 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_314 : STD_LOGIC; 
  signal mac_control_phyrstcnt_129_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_277 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_213 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_278 : STD_LOGIC; 
  signal mac_control_phyrstcnt_131_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_131_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_214 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_316 : STD_LOGIC; 
  signal mac_control_phyrstcnt_131_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_279 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_215 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_280 : STD_LOGIC; 
  signal mac_control_phyrstcnt_133_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_133_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_216 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_318 : STD_LOGIC; 
  signal mac_control_phyrstcnt_133_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_281 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_217 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_282 : STD_LOGIC; 
  signal mac_control_phyrstcnt_135_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_135_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_218 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_320 : STD_LOGIC; 
  signal mac_control_phyrstcnt_135_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_283 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_219 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_284 : STD_LOGIC; 
  signal mac_control_phyrstcnt_137_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_137_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_220 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_322 : STD_LOGIC; 
  signal mac_control_phyrstcnt_137_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_285 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_221 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_286 : STD_LOGIC; 
  signal mac_control_phyrstcnt_139_CYMUXG : STD_LOGIC; 
  signal mac_control_phyrstcnt_139_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_222 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_cy_324 : STD_LOGIC; 
  signal mac_control_phyrstcnt_139_CYINIT : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_287 : STD_LOGIC; 
  signal rx_input_data_6_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_lut3_223 : STD_LOGIC; 
  signal mac_control_phyrstcnt_inst_sum_288 : STD_LOGIC; 
  signal mac_control_phyrstcnt_141_CYINIT : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_1_rt : STD_LOGIC; 
  signal rx_input_memio_macnt_70_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_56 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_253 : STD_LOGIC; 
  signal rx_input_memio_macnt_70_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_219 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_57 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_220 : STD_LOGIC; 
  signal rx_input_memio_macnt_71_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_71_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_71_XORG : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_58 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_255 : STD_LOGIC; 
  signal rx_input_memio_macnt_71_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_59 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_222 : STD_LOGIC; 
  signal rx_input_memio_macnt_73_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_73_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_60 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_257 : STD_LOGIC; 
  signal rx_input_memio_macnt_73_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_223 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_18_CYINIT : STD_LOGIC; 
  signal rx_input_memio_dout_7_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_31_rt : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_rxoferr_cnt_30_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_rst_rt : STD_LOGIC; 
  signal mac_control_ledrx_cnt_154_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_236 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_340 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_154_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_301 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_237 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_302 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_238 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_342 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_303 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_239 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_304 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_240 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_344 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_305 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_241 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_306 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_242 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_346 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_307 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_243 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_308 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_244 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_348 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_309 : STD_LOGIC; 
  signal rx_input_memio_dout_9_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_245 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_310 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163_CYMUXG : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_246 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_cy_350 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163_CYINIT : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_311 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_lut3_247 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_inst_sum_312 : STD_LOGIC; 
  signal mac_control_ledrx_cnt_165_CYINIT : STD_LOGIC; 
  signal tx_output_bcntl_1_rt : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_195_CYMUXG : STD_LOGIC; 
  signal tx_output_SIG_19 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_194 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut1_61_O : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_197_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut1_71_O : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_196 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_197_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_197_CYINIT : STD_LOGIC; 
  signal tx_output_bcntl_3_rt : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_199_CYMUXG : STD_LOGIC; 
  signal tx_output_SIG_20 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_198 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_199_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_199_CYINIT : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut4_161_O : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_201_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut4_171_O : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_200 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_201_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_201_CYINIT : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut4_18 : STD_LOGIC; 
  signal tx_output_n0035_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_lut4_19 : STD_LOGIC; 
  signal tx_output_Mcompar_n0035_inst_cy_202 : STD_LOGIC; 
  signal tx_output_n0035_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_n0035_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_20_CYINIT : STD_LOGIC; 
  signal rx_output_cs_FFd5_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_31_rt : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_rxphyerr_cnt_30_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_18_CYINIT : STD_LOGIC; 
  signal rx_input_data_0_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_31_rt : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_rxfifowerr_cnt_30_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_31_rt : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_txfifowerr_cnt_30_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_2_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0042_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_2_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_2_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_79 : STD_LOGIC; 
  signal rx_output_bp_0_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_80 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_86 : STD_LOGIC; 
  signal rx_output_bp_0_CYINIT : STD_LOGIC; 
  signal rx_output_bp_0_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_81 : STD_LOGIC; 
  signal rx_output_bp_2_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_82 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_88 : STD_LOGIC; 
  signal rx_output_bp_2_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_83 : STD_LOGIC; 
  signal rx_output_bp_4_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_84 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_90 : STD_LOGIC; 
  signal rx_output_bp_4_CYINIT : STD_LOGIC; 
  signal rx_input_data_1_FFY_RST : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_85 : STD_LOGIC; 
  signal rx_output_bp_6_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_86 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_92 : STD_LOGIC; 
  signal rx_output_bp_6_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_87 : STD_LOGIC; 
  signal rx_output_bp_8_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_88 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_94 : STD_LOGIC; 
  signal rx_output_bp_8_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_89 : STD_LOGIC; 
  signal rx_output_bp_10_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_90 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_96 : STD_LOGIC; 
  signal rx_output_bp_10_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_91 : STD_LOGIC; 
  signal rx_output_bp_12_CYMUXG : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_lut2_92 : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_98 : STD_LOGIC; 
  signal rx_output_bp_12_CYINIT : STD_LOGIC; 
  signal rx_output_bp_14_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_bp_14_FROM : STD_LOGIC; 
  signal rx_output_bp_15_rt : STD_LOGIC; 
  signal rx_output_Madd_lbp_inst_cy_100 : STD_LOGIC; 
  signal rx_output_bp_14_CYINIT : STD_LOGIC; 
  signal tx_output_cs_FFd12_rt : STD_LOGIC; 
  signal tx_output_bcnt_38_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_40 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_204 : STD_LOGIC; 
  signal tx_output_bcnt_38_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_171 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_41 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_172 : STD_LOGIC; 
  signal tx_output_bcnt_39_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_39_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_42 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_206 : STD_LOGIC; 
  signal tx_output_bcnt_39_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_173 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_43 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_174 : STD_LOGIC; 
  signal tx_output_bcnt_41_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_41_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_44 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_208 : STD_LOGIC; 
  signal tx_output_bcnt_41_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_175 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_45 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_176 : STD_LOGIC; 
  signal tx_output_bcnt_43_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_43_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_46 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_210 : STD_LOGIC; 
  signal tx_output_bcnt_43_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_177 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_47 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_178 : STD_LOGIC; 
  signal tx_output_bcnt_45_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_45_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_48 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_212 : STD_LOGIC; 
  signal tx_output_bcnt_45_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_179 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_49 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_180 : STD_LOGIC; 
  signal tx_output_bcnt_47_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_47_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_50 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_214 : STD_LOGIC; 
  signal tx_output_bcnt_47_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_181 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_51 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_182 : STD_LOGIC; 
  signal tx_output_bcnt_49_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_49_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_52 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_216 : STD_LOGIC; 
  signal tx_output_bcnt_49_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_183 : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_53 : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_184 : STD_LOGIC; 
  signal tx_output_bcnt_51_CYMUXG : STD_LOGIC; 
  signal tx_output_bcnt_51_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_bcnt_inst_lut3_54 : STD_LOGIC; 
  signal tx_output_bcnt_inst_cy_218 : STD_LOGIC; 
  signal tx_output_bcnt_51_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_inst_sum_185 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_3_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0039_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_3_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_3_CYINIT : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_0 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_79_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_1 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_78 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_2 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_81_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_3 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_80 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_81_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_81_CYINIT : STD_LOGIC; 
  signal rx_input_data_2_FFY_RST : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_4 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_83_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_5 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_82 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_83_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_83_CYINIT : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_6 : STD_LOGIC; 
  signal rx_output_n0017_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_lut4_7 : STD_LOGIC; 
  signal rx_output_Mcompar_n0017_inst_cy_84 : STD_LOGIC; 
  signal rx_output_n0017_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0017_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_111 : STD_LOGIC; 
  signal rx_fifocheck_diff_0_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_112 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_161 : STD_LOGIC; 
  signal rx_fifocheck_diff_0_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_diff_0_LOGIC_ONE : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_113 : STD_LOGIC; 
  signal rx_fifocheck_diff_2_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_114 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_163 : STD_LOGIC; 
  signal rx_fifocheck_diff_2_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_115 : STD_LOGIC; 
  signal rx_fifocheck_diff_4_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_116 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_165 : STD_LOGIC; 
  signal rx_fifocheck_diff_4_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_117 : STD_LOGIC; 
  signal rx_fifocheck_diff_6_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_118 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_167 : STD_LOGIC; 
  signal rx_fifocheck_diff_6_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_119 : STD_LOGIC; 
  signal rx_fifocheck_diff_8_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_120 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_169 : STD_LOGIC; 
  signal rx_fifocheck_diff_8_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_121 : STD_LOGIC; 
  signal rx_fifocheck_diff_10_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_122 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_171 : STD_LOGIC; 
  signal rx_fifocheck_diff_10_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_123 : STD_LOGIC; 
  signal rx_fifocheck_diff_12_CYMUXG : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_124 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_173 : STD_LOGIC; 
  signal rx_fifocheck_diff_12_CYINIT : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_125 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_lut2_126 : STD_LOGIC; 
  signal rx_fifocheck_Msub_n0001_inst_cy_175 : STD_LOGIC; 
  signal rx_fifocheck_diff_14_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_111 : STD_LOGIC; 
  signal tx_fifocheck_diff_0_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_112 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_161 : STD_LOGIC; 
  signal tx_fifocheck_diff_0_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_0_LOGIC_ONE : STD_LOGIC; 
  signal tx_fifocheck_diff_2_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_113 : STD_LOGIC; 
  signal tx_fifocheck_diff_2_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_114 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_163 : STD_LOGIC; 
  signal tx_fifocheck_diff_2_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_4_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_115 : STD_LOGIC; 
  signal tx_fifocheck_diff_4_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_116 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_165 : STD_LOGIC; 
  signal tx_fifocheck_diff_4_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_6_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_117 : STD_LOGIC; 
  signal tx_fifocheck_diff_6_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_118 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_167 : STD_LOGIC; 
  signal tx_fifocheck_diff_6_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_8_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_119 : STD_LOGIC; 
  signal tx_fifocheck_diff_8_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_120 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_169 : STD_LOGIC; 
  signal tx_fifocheck_diff_8_CYINIT : STD_LOGIC; 
  signal rx_input_data_3_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_10_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_121 : STD_LOGIC; 
  signal tx_fifocheck_diff_10_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_122 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_171 : STD_LOGIC; 
  signal tx_fifocheck_diff_10_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_12_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_123 : STD_LOGIC; 
  signal tx_fifocheck_diff_12_CYMUXG : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_124 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_173 : STD_LOGIC; 
  signal tx_fifocheck_diff_12_CYINIT : STD_LOGIC; 
  signal tx_fifocheck_diff_14_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_125 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_lut2_126 : STD_LOGIC; 
  signal tx_fifocheck_Msub_n0001_inst_cy_175 : STD_LOGIC; 
  signal tx_fifocheck_diff_14_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_142_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_rst_rt : STD_LOGIC; 
  signal mac_control_ledtx_cnt_142_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_224 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_327 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_142_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_289 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_225 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_290 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_226 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_329 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_291 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_227 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_292 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_228 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_331 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_293 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_229 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_294 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_230 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_333 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_295 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_231 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_296 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_232 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_335 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_297 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_233 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_298 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151_CYMUXG : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_234 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_cy_337 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151_CYINIT : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_299 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_lut3_235 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_inst_sum_300 : STD_LOGIC; 
  signal mac_control_ledtx_cnt_153_CYINIT : STD_LOGIC; 
  signal tx_output_bcnt_53_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1912 : STD_LOGIC; 
  signal rx_output_fifo_N1904 : STD_LOGIC; 
  signal rx_output_fifo_N17_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N17_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1914 : STD_LOGIC; 
  signal rx_output_fifo_N17_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N17_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N1905 : STD_LOGIC; 
  signal rx_output_fifo_N15_FROM : STD_LOGIC; 
  signal rx_output_fifo_N1906 : STD_LOGIC; 
  signal rx_output_fifo_N15_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N15_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1924 : STD_LOGIC; 
  signal rx_output_fifo_N15_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N1907 : STD_LOGIC; 
  signal rx_output_fifo_N13_FROM : STD_LOGIC; 
  signal rx_output_fifo_N1908 : STD_LOGIC; 
  signal rx_output_fifo_N13_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N13_GROM : STD_LOGIC; 
  signal rx_output_fifo_N1934 : STD_LOGIC; 
  signal rx_output_fifo_N13_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N1909 : STD_LOGIC; 
  signal rx_output_fifo_N11_FROM : STD_LOGIC; 
  signal rx_output_fifo_N1910 : STD_LOGIC; 
  signal rx_output_fifo_N10_rt : STD_LOGIC; 
  signal rx_output_fifo_N1944 : STD_LOGIC; 
  signal rx_output_fifo_N11_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N1911 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_95 : STD_LOGIC; 
  signal tx_input_n0074_0_XORF : STD_LOGIC; 
  signal tx_input_n0074_0_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_0_XORG : STD_LOGIC; 
  signal tx_input_n0074_0_GROM : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_118 : STD_LOGIC; 
  signal tx_input_n0074_0_CYINIT : STD_LOGIC; 
  signal tx_input_n0074_0_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_97 : STD_LOGIC; 
  signal tx_input_n0074_2_XORF : STD_LOGIC; 
  signal tx_input_n0074_2_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_2_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_98 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_120 : STD_LOGIC; 
  signal tx_input_n0074_2_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_99 : STD_LOGIC; 
  signal tx_input_n0074_4_XORF : STD_LOGIC; 
  signal tx_input_n0074_4_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_4_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_100 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_122 : STD_LOGIC; 
  signal tx_input_n0074_4_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_101 : STD_LOGIC; 
  signal tx_input_n0074_6_XORF : STD_LOGIC; 
  signal tx_input_n0074_6_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_6_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_102 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_124 : STD_LOGIC; 
  signal tx_input_n0074_6_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_103 : STD_LOGIC; 
  signal tx_input_n0074_8_XORF : STD_LOGIC; 
  signal tx_input_n0074_8_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_8_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_104 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_126 : STD_LOGIC; 
  signal tx_input_n0074_8_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_105 : STD_LOGIC; 
  signal tx_input_n0074_10_XORF : STD_LOGIC; 
  signal tx_input_n0074_10_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_10_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_106 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_128 : STD_LOGIC; 
  signal tx_input_n0074_10_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_107 : STD_LOGIC; 
  signal tx_input_n0074_12_XORF : STD_LOGIC; 
  signal tx_input_n0074_12_CYMUXG : STD_LOGIC; 
  signal tx_input_n0074_12_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_108 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_130 : STD_LOGIC; 
  signal tx_input_n0074_12_CYINIT : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_109 : STD_LOGIC; 
  signal tx_input_n0074_14_XORF : STD_LOGIC; 
  signal tx_input_n0074_14_XORG : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_lut2_110 : STD_LOGIC; 
  signal tx_input_Msub_n0034_inst_cy_132 : STD_LOGIC; 
  signal tx_input_n0074_14_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_1_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0045_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_1_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_1_CYINIT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd5_rt : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_32_CYMUXG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_34 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_187 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_32_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_165 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_35 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_166 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33_CYMUXG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_36 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_189 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33_CYINIT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_167 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_37 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_168 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35_CYMUXG : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_38 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_191 : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35_CYINIT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_169 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_0 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_79_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_1 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_78 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_2 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_81_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_3 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_80 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_81_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_81_CYINIT : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_4 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_83_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_5 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_82 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_83_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_83_CYINIT : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_6 : STD_LOGIC; 
  signal rx_output_n0018_CYMUXG : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_lut4_7 : STD_LOGIC; 
  signal rx_output_Mcompar_n0018_inst_cy_84 : STD_LOGIC; 
  signal rx_output_n0018_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0018_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_txf_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_txf_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_txf_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_txf_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_txf_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_txf_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_txf_cnt_10_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_txf_cnt_12_CYINIT : STD_LOGIC; 
  signal tx_output_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_txf_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_txf_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_txf_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_txf_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_txf_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_txf_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_txf_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_txf_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_txf_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_txf_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_txf_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_txf_cnt_31_rt : STD_LOGIC; 
  signal mac_control_txf_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_txf_cnt_30_CYINIT : STD_LOGIC; 
  signal rx_output_cs_FFd19_rt : STD_LOGIC; 
  signal addr3ext_0_CYMUXG : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_0 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_101 : STD_LOGIC; 
  signal addr3ext_0_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_95 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_1 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_96 : STD_LOGIC; 
  signal addr3ext_1_CYMUXG : STD_LOGIC; 
  signal addr3ext_1_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_2 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_103 : STD_LOGIC; 
  signal addr3ext_1_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_97 : STD_LOGIC; 
  signal rx_input_data_4_FFY_RST : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_3 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_98 : STD_LOGIC; 
  signal addr3ext_3_CYMUXG : STD_LOGIC; 
  signal addr3ext_3_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_4 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_105 : STD_LOGIC; 
  signal addr3ext_3_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_99 : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_5 : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_100 : STD_LOGIC; 
  signal addr3ext_5_CYMUXG : STD_LOGIC; 
  signal addr3ext_5_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_macnt_inst_lut3_6 : STD_LOGIC; 
  signal rx_output_macnt_inst_cy_107 : STD_LOGIC; 
  signal addr3ext_5_CYINIT : STD_LOGIC; 
  signal rx_output_macnt_inst_sum_101 : STD_LOGIC; 
  signal tx_output_data_0_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_61 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_224 : STD_LOGIC; 
  signal rx_input_memio_macnt_75_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_75_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_62 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_259 : STD_LOGIC; 
  signal rx_input_memio_macnt_75_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_225 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_63 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_226 : STD_LOGIC; 
  signal rx_input_memio_macnt_77_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_77_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_64 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_261 : STD_LOGIC; 
  signal rx_input_memio_macnt_77_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_227 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_65 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_228 : STD_LOGIC; 
  signal rx_input_memio_macnt_79_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_79_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_66 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_263 : STD_LOGIC; 
  signal rx_input_memio_macnt_79_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_229 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_67 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_230 : STD_LOGIC; 
  signal rx_input_memio_macnt_81_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_81_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_68 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_265 : STD_LOGIC; 
  signal rx_input_memio_macnt_81_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_231 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_69 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_232 : STD_LOGIC; 
  signal rx_input_memio_macnt_83_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_macnt_83_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_70 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_cy_267 : STD_LOGIC; 
  signal rx_input_memio_macnt_83_CYINIT : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_233 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_lut3_71 : STD_LOGIC; 
  signal rx_input_memio_macnt_inst_sum_234 : STD_LOGIC; 
  signal rx_input_memio_macnt_85_CYINIT : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_lut2_641_O : STD_LOGIC; 
  signal rx_output_n0070_2_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_2_XORG : STD_LOGIC; 
  signal rx_output_n0070_2_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_63 : STD_LOGIC; 
  signal rx_output_n0070_2_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_3_FROM : STD_LOGIC; 
  signal rx_output_n0070_3_XORF : STD_LOGIC; 
  signal rx_output_n0070_3_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_3_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_3_XORG : STD_LOGIC; 
  signal rx_output_n0070_3_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_65 : STD_LOGIC; 
  signal rx_output_n0070_3_CYINIT : STD_LOGIC; 
  signal rx_output_n0070_5_FROM : STD_LOGIC; 
  signal rx_output_n0070_5_XORF : STD_LOGIC; 
  signal rx_output_n0070_5_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_5_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_5_XORG : STD_LOGIC; 
  signal rx_output_n0070_5_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_67 : STD_LOGIC; 
  signal rx_output_n0070_5_CYINIT : STD_LOGIC; 
  signal rx_output_n0070_7_FROM : STD_LOGIC; 
  signal rx_output_n0070_7_XORF : STD_LOGIC; 
  signal rx_output_n0070_7_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_7_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_7_XORG : STD_LOGIC; 
  signal rx_output_n0070_7_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_69 : STD_LOGIC; 
  signal rx_output_n0070_7_CYINIT : STD_LOGIC; 
  signal rx_output_n0070_9_FROM : STD_LOGIC; 
  signal rx_output_n0070_9_XORF : STD_LOGIC; 
  signal rx_output_n0070_9_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_9_XORG : STD_LOGIC; 
  signal rx_output_n0070_9_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_71 : STD_LOGIC; 
  signal rx_output_n0070_9_CYINIT : STD_LOGIC; 
  signal rx_output_n0070_11_FROM : STD_LOGIC; 
  signal rx_output_n0070_11_XORF : STD_LOGIC; 
  signal rx_output_n0070_11_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_11_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_11_XORG : STD_LOGIC; 
  signal rx_output_n0070_11_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_73 : STD_LOGIC; 
  signal rx_output_n0070_11_CYINIT : STD_LOGIC; 
  signal rx_output_n0070_13_FROM : STD_LOGIC; 
  signal rx_output_n0070_13_XORF : STD_LOGIC; 
  signal rx_output_n0070_13_CYMUXG : STD_LOGIC; 
  signal rx_output_n0070_13_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_n0070_13_XORG : STD_LOGIC; 
  signal rx_output_n0070_13_GROM : STD_LOGIC; 
  signal rx_output_Madd_n0047_inst_cy_75 : STD_LOGIC; 
  signal rx_output_n0070_13_CYINIT : STD_LOGIC; 
  signal rx_output_SIG_38 : STD_LOGIC; 
  signal rx_output_n0070_15_XORF : STD_LOGIC; 
  signal rx_output_n0070_15_CYINIT : STD_LOGIC; 
  signal rx_input_data_7_FFY_RST : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_0 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_79_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_1 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_78 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ONE : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_2 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_81_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_3 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_80 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_81_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_81_CYINIT : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_4 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_83_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_5 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_82 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_83_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_83_CYINIT : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_6 : STD_LOGIC; 
  signal tx_output_n0006_CYMUXG : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_lut4_7 : STD_LOGIC; 
  signal tx_output_Mcompar_n0006_inst_cy_84 : STD_LOGIC; 
  signal tx_output_n0006_LOGIC_ZERO : STD_LOGIC; 
  signal tx_output_n0006_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_0_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0048_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_0_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_0_CYINIT : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_149 : STD_LOGIC; 
  signal rx_input_memio_bcntl_0_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_150 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_237 : STD_LOGIC; 
  signal rx_input_memio_bcntl_0_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_0_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_bcntl_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_2_FROM : STD_LOGIC; 
  signal rx_input_memio_bcntl_2_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_152 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_239 : STD_LOGIC; 
  signal rx_input_memio_bcntl_2_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_153 : STD_LOGIC; 
  signal rx_input_memio_bcntl_4_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_154 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_241 : STD_LOGIC; 
  signal rx_input_memio_bcntl_4_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_6_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_155 : STD_LOGIC; 
  signal rx_input_memio_bcntl_6_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_156 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_243 : STD_LOGIC; 
  signal rx_input_memio_bcntl_6_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_8_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_157 : STD_LOGIC; 
  signal rx_input_memio_bcntl_8_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_158 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_245 : STD_LOGIC; 
  signal rx_input_memio_bcntl_8_CYINIT : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_10_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_159 : STD_LOGIC; 
  signal rx_input_memio_bcntl_10_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_160 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_247 : STD_LOGIC; 
  signal rx_input_memio_bcntl_10_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_12_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_161 : STD_LOGIC; 
  signal rx_input_memio_bcntl_12_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_162 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_249 : STD_LOGIC; 
  signal rx_input_memio_bcntl_12_CYINIT : STD_LOGIC; 
  signal rx_input_memio_bcntl_14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_163 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_lut2_164 : STD_LOGIC; 
  signal rx_input_memio_Msub_n0042_inst_cy_251 : STD_LOGIC; 
  signal rx_input_memio_bcntl_14_CYINIT : STD_LOGIC; 
  signal tx_input_addr_16_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd12_rt : STD_LOGIC; 
  signal tx_input_addr_16_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_16 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_134 : STD_LOGIC; 
  signal tx_input_addr_16_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_sum_127 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_17 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_128 : STD_LOGIC; 
  signal tx_input_addr_17_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_17_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_18 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_136 : STD_LOGIC; 
  signal tx_input_addr_17_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_129 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_19 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_130 : STD_LOGIC; 
  signal tx_input_addr_19_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_19_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_20 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_138 : STD_LOGIC; 
  signal tx_input_addr_19_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_131 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_21 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_132 : STD_LOGIC; 
  signal tx_input_addr_21_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_21_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_22 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_140 : STD_LOGIC; 
  signal tx_input_addr_21_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_133 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_23 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_134 : STD_LOGIC; 
  signal tx_input_addr_23_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_23_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_24 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_142 : STD_LOGIC; 
  signal tx_input_addr_23_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_135 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_25 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_136 : STD_LOGIC; 
  signal tx_input_addr_25_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_25_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_26 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_144 : STD_LOGIC; 
  signal tx_input_addr_25_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_137 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_27 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_138 : STD_LOGIC; 
  signal tx_input_addr_27_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_27_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_28 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_146 : STD_LOGIC; 
  signal tx_input_addr_27_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_139 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_29 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_140 : STD_LOGIC; 
  signal tx_input_addr_29_CYMUXG : STD_LOGIC; 
  signal tx_input_addr_29_LOGIC_ZERO : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_30 : STD_LOGIC; 
  signal tx_input_addr_inst_cy_148 : STD_LOGIC; 
  signal tx_input_addr_29_CYINIT : STD_LOGIC; 
  signal tx_input_addr_inst_sum_141 : STD_LOGIC; 
  signal tx_input_addr_inst_lut3_31 : STD_LOGIC; 
  signal tx_input_addr_inst_sum_142 : STD_LOGIC; 
  signal tx_input_addr_31_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_lut2_16 : STD_LOGIC; 
  signal mac_control_rxf_cnt_0_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_0_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_16 : STD_LOGIC; 
  signal mac_control_rxf_cnt_0_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_2_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_2_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_2_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_2_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_18 : STD_LOGIC; 
  signal mac_control_rxf_cnt_2_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_4_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_4_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_4_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_4_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_20 : STD_LOGIC; 
  signal mac_control_rxf_cnt_4_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_6_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_6_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_6_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_6_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_22 : STD_LOGIC; 
  signal mac_control_rxf_cnt_6_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_8_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_8_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_8_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_8_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_24 : STD_LOGIC; 
  signal mac_control_rxf_cnt_8_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_10_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_10_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_10_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_10_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_26 : STD_LOGIC; 
  signal mac_control_rxf_cnt_10_CYINIT : STD_LOGIC; 
  signal rx_output_cs_FFd9_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cnt_12_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_12_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_12_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_12_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_28 : STD_LOGIC; 
  signal mac_control_rxf_cnt_12_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_14_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_14_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_14_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_14_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_30 : STD_LOGIC; 
  signal mac_control_rxf_cnt_14_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_16_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_16_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_16_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_16_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_32 : STD_LOGIC; 
  signal mac_control_rxf_cnt_16_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_18_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_18_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_18_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_18_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_34 : STD_LOGIC; 
  signal mac_control_rxf_cnt_18_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_20_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_20_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_20_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_20_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_36 : STD_LOGIC; 
  signal mac_control_rxf_cnt_20_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_22_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_22_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_22_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_22_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_38 : STD_LOGIC; 
  signal mac_control_rxf_cnt_22_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_24_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_24_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_24_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_24_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_40 : STD_LOGIC; 
  signal mac_control_rxf_cnt_24_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_26_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_26_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_26_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_26_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_42 : STD_LOGIC; 
  signal mac_control_rxf_cnt_26_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_28_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_28_CYMUXG : STD_LOGIC; 
  signal mac_control_rxf_cnt_28_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_28_GROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_44 : STD_LOGIC; 
  signal mac_control_rxf_cnt_28_CYINIT : STD_LOGIC; 
  signal mac_control_rxf_cnt_30_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_rxf_cnt_30_FROM : STD_LOGIC; 
  signal mac_control_rxf_cnt_31_rt : STD_LOGIC; 
  signal mac_control_rxf_cnt_Madd_n0000_inst_cy_46 : STD_LOGIC; 
  signal mac_control_rxf_cnt_30_CYINIT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_4_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_2_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_4_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_6_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_8_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_8_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_10_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_12 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_13 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_177 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ONE : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_14 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_5_CYMUXG : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_15 : STD_LOGIC; 
  signal rx_input_memio_addrchk_Mcompar_n0033_inst_cy_179 : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_5_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_5_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N2840 : STD_LOGIC; 
  signal rx_output_fifo_N2832 : STD_LOGIC; 
  signal rx_output_fifo_N9_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N9_GROM : STD_LOGIC; 
  signal rx_output_fifo_N2842 : STD_LOGIC; 
  signal rx_output_fifo_N9_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N2833 : STD_LOGIC; 
  signal rx_output_fifo_N7_FROM : STD_LOGIC; 
  signal rx_output_fifo_N2834 : STD_LOGIC; 
  signal rx_output_fifo_N7_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N7_GROM : STD_LOGIC; 
  signal rx_output_fifo_N2852 : STD_LOGIC; 
  signal rx_output_fifo_N7_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N2835 : STD_LOGIC; 
  signal rx_output_fifo_N5_FROM : STD_LOGIC; 
  signal rx_output_fifo_N2836 : STD_LOGIC; 
  signal rx_output_fifo_N5_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N5_GROM : STD_LOGIC; 
  signal rx_output_fifo_N2862 : STD_LOGIC; 
  signal rx_output_fifo_N5_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N2837 : STD_LOGIC; 
  signal rx_output_fifo_N3_FROM : STD_LOGIC; 
  signal rx_output_fifo_N2838 : STD_LOGIC; 
  signal rx_output_fifo_N2_rt : STD_LOGIC; 
  signal rx_output_fifo_N2872 : STD_LOGIC; 
  signal rx_output_fifo_N3_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N2839 : STD_LOGIC; 
  signal rx_output_fifo_N2569 : STD_LOGIC; 
  signal rx_output_fifo_N2576_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N2568 : STD_LOGIC; 
  signal rx_output_fifo_N2577 : STD_LOGIC; 
  signal rx_output_fifo_N2576_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N2576_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_fifo_N2567 : STD_LOGIC; 
  signal rx_output_fifo_N2574_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N2566 : STD_LOGIC; 
  signal rx_output_fifo_N2575 : STD_LOGIC; 
  signal rx_output_fifo_N2574_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N2574_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N2565 : STD_LOGIC; 
  signal rx_output_fifo_N2572_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N2564 : STD_LOGIC; 
  signal rx_output_fifo_N2573 : STD_LOGIC; 
  signal rx_output_fifo_N2572_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N2572_CYINIT : STD_LOGIC; 
  signal tx_output_crcl_6_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N2563 : STD_LOGIC; 
  signal rx_output_fifo_BU172_O_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N2562 : STD_LOGIC; 
  signal rx_output_fifo_N2571 : STD_LOGIC; 
  signal rx_output_fifo_BU172_O_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_BU172_O_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_empty_FROM : STD_LOGIC; 
  signal rx_output_fifo_N2580 : STD_LOGIC; 
  signal rx_output_fifo_empty_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N3607 : STD_LOGIC; 
  signal rx_output_fifo_N3614_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N3606 : STD_LOGIC; 
  signal rx_output_fifo_N3615 : STD_LOGIC; 
  signal rx_output_fifo_N3614_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N3614_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_fifo_N3605 : STD_LOGIC; 
  signal rx_output_fifo_N3612_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N3604 : STD_LOGIC; 
  signal rx_output_fifo_N3613 : STD_LOGIC; 
  signal rx_output_fifo_N3612_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N3612_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N3603 : STD_LOGIC; 
  signal rx_output_fifo_N3610_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N3602 : STD_LOGIC; 
  signal rx_output_fifo_N3611 : STD_LOGIC; 
  signal rx_output_fifo_N3610_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_N3610_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N3601 : STD_LOGIC; 
  signal rx_output_fifo_BU351_O_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N3600 : STD_LOGIC; 
  signal rx_output_fifo_N3609 : STD_LOGIC; 
  signal rx_output_fifo_BU351_O_LOGIC_ZERO : STD_LOGIC; 
  signal rx_output_fifo_BU351_O_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_full_FROM : STD_LOGIC; 
  signal rx_output_fifo_N3618 : STD_LOGIC; 
  signal rx_output_fifo_full_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N4756 : STD_LOGIC; 
  signal rx_output_fifo_N4763_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N4760 : STD_LOGIC; 
  signal rx_output_fifo_N4759 : STD_LOGIC; 
  signal rx_output_fifo_N4763_LOGIC_ONE : STD_LOGIC; 
  signal rx_output_fifo_N4764 : STD_LOGIC; 
  signal rx_output_fifo_N4771_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N4768 : STD_LOGIC; 
  signal rx_output_fifo_N4767 : STD_LOGIC; 
  signal rx_output_fifo_N4771_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N4772 : STD_LOGIC; 
  signal rx_output_fifo_N4779_CYMUXG : STD_LOGIC; 
  signal rx_output_fifo_N4776 : STD_LOGIC; 
  signal rx_output_fifo_N4775 : STD_LOGIC; 
  signal rx_output_fifo_N4779_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N4780 : STD_LOGIC; 
  signal rx_output_fifo_N4754 : STD_LOGIC; 
  signal rx_output_fifo_N4786 : STD_LOGIC; 
  signal rx_output_fifo_N4783 : STD_LOGIC; 
  signal rx_output_fifo_wrcount_0_CYINIT : STD_LOGIC; 
  signal rx_output_fifo_N4755 : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_103_rt : STD_LOGIC; 
  signal mac_control_bitcnt_104_CYMUXG : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_186 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_287 : STD_LOGIC; 
  signal mac_control_bitcnt_104_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_251 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_187 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_252 : STD_LOGIC; 
  signal mac_control_bitcnt_105_CYMUXG : STD_LOGIC; 
  signal mac_control_bitcnt_105_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_188 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_289 : STD_LOGIC; 
  signal mac_control_bitcnt_105_CYINIT : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_253 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_189 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_254 : STD_LOGIC; 
  signal mac_control_bitcnt_107_CYMUXG : STD_LOGIC; 
  signal mac_control_bitcnt_107_LOGIC_ZERO : STD_LOGIC; 
  signal mac_control_bitcnt_inst_lut3_190 : STD_LOGIC; 
  signal mac_control_bitcnt_inst_cy_291 : STD_LOGIC; 
  signal mac_control_bitcnt_107_CYINIT : STD_LOGIC; 
  signal mac_control_bitcnt_inst_sum_255 : STD_LOGIC; 
  signal tx_output_crc_loigc_n0115_0_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_n0115_0_GROM : STD_LOGIC; 
  signal rx_input_memio_n0048_15_1_O : STD_LOGIC; 
  signal rx_input_memio_n0048_12_1_O : STD_LOGIC; 
  signal rx_input_memio_n0048_31_Q : STD_LOGIC; 
  signal rx_input_memio_crcl_31_GROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O_GROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd15_FROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd15_In7_O : STD_LOGIC; 
  signal rx_input_memio_menl_FROM : STD_LOGIC; 
  signal rx_input_memio_menl_GROM : STD_LOGIC; 
  signal rx_input_memio_menl_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_n0019_SW0_O_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_n0019_SW0_O_GROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_n0115_0_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_n0115_0_GROM : STD_LOGIC; 
  signal tx_input_Ker3585921_O_FROM : STD_LOGIC; 
  signal tx_input_Ker3585921_O_GROM : STD_LOGIC; 
  signal rx_input_endf_GROM : STD_LOGIC; 
  signal tx_output_n0034_15_1_O : STD_LOGIC; 
  signal tx_output_n0034_5_1_O : STD_LOGIC; 
  signal tx_input_Ker35859120_O_FROM : STD_LOGIC; 
  signal tx_input_Ker35859120_O_GROM : STD_LOGIC; 
  signal rx_input_memio_n0048_22_Q : STD_LOGIC; 
  signal rx_input_memio_n0048_5_1_O : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_n0005_Result1_O_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_n0005_Result1_O_GROM : STD_LOGIC; 
  signal rx_output_lenr_10_FROM : STD_LOGIC; 
  signal rx_output_n0046_10_O : STD_LOGIC; 
  signal rx_output_lenr_10_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_11_FROM : STD_LOGIC; 
  signal rx_output_n0046_11_O : STD_LOGIC; 
  signal rx_output_lenr_11_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_12_FROM : STD_LOGIC; 
  signal rx_output_n0046_12_O : STD_LOGIC; 
  signal rx_output_lenr_12_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_13_FROM : STD_LOGIC; 
  signal rx_output_n0046_13_O : STD_LOGIC; 
  signal rx_output_lenr_13_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_14_FROM : STD_LOGIC; 
  signal rx_output_n0046_14_O : STD_LOGIC; 
  signal rx_output_lenr_14_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_15_FROM : STD_LOGIC; 
  signal rx_output_n0046_15_O : STD_LOGIC; 
  signal rx_output_lenr_15_CEMUXNOT : STD_LOGIC; 
  signal tx_input_N35872_FROM : STD_LOGIC; 
  signal tx_input_N35872_GROM : STD_LOGIC; 
  signal tx_output_crc_0_FROM : STD_LOGIC; 
  signal tx_output_crc_0_GROM : STD_LOGIC; 
  signal rx_output_lenr_2_FROM : STD_LOGIC; 
  signal rx_output_n0046_2_O : STD_LOGIC; 
  signal rx_output_lenr_2_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_3_FROM : STD_LOGIC; 
  signal rx_output_n0046_3_O : STD_LOGIC; 
  signal rx_output_lenr_3_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_4_FROM : STD_LOGIC; 
  signal rx_output_n0046_4_O : STD_LOGIC; 
  signal rx_output_lenr_4_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_5_FROM : STD_LOGIC; 
  signal rx_output_n0046_5_O : STD_LOGIC; 
  signal rx_output_lenr_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcenl_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcenl_FROM : STD_LOGIC; 
  signal tx_output_crcenl_GROM : STD_LOGIC; 
  signal rx_output_lenr_6_FROM : STD_LOGIC; 
  signal rx_output_n0046_6_O : STD_LOGIC; 
  signal rx_output_lenr_6_CEMUXNOT : STD_LOGIC; 
  signal macaddr_1_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_7_FROM : STD_LOGIC; 
  signal rx_output_n0046_7_O : STD_LOGIC; 
  signal rx_output_lenr_7_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_8_FROM : STD_LOGIC; 
  signal rx_output_n0046_8_O : STD_LOGIC; 
  signal rx_output_lenr_8_CEMUXNOT : STD_LOGIC; 
  signal rx_output_lenr_9_FROM : STD_LOGIC; 
  signal rx_output_n0046_9_O : STD_LOGIC; 
  signal rx_output_lenr_9_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_n001618_O_FROM : STD_LOGIC; 
  signal rx_input_memio_n001618_O_GROM : STD_LOGIC; 
  signal rx_output_n0043_SW1_O_FROM : STD_LOGIC; 
  signal rx_output_n0043_SW1_O_GROM : STD_LOGIC; 
  signal mac_control_n0085_FROM : STD_LOGIC; 
  signal mac_control_n0085_GROM : STD_LOGIC; 
  signal tx_input_cs_FFd6_In : STD_LOGIC; 
  signal tx_input_cs_FFd5_In1_O : STD_LOGIC; 
  signal macaddr_1_FFX_RST : STD_LOGIC; 
  signal tx_input_cs_FFd8_In1_O : STD_LOGIC; 
  signal tx_input_cs_FFd7_In1_O : STD_LOGIC; 
  signal rx_input_memio_crc_0_FROM : STD_LOGIC; 
  signal rx_input_memio_crc_0_GROM : STD_LOGIC; 
  signal rx_input_fifo_rd_en_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_rd_en_FROM : STD_LOGIC; 
  signal rx_input_fifo_rd_en_GROM : STD_LOGIC; 
  signal mac_control_phyaddr_31_GROM : STD_LOGIC; 
  signal tx_output_addrinc_SW0_O_FROM : STD_LOGIC; 
  signal tx_output_addrinc_SW0_O_GROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O_FROM : STD_LOGIC; 
  signal tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O_GROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_n0005_Result1_O_FROM : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_n0005_Result1_O_GROM : STD_LOGIC; 
  signal mac_control_n0046 : STD_LOGIC; 
  signal mac_control_n0048 : STD_LOGIC; 
  signal mac_control_txf_rst_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd4_In : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd3_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd10_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd9_In : STD_LOGIC; 
  signal macaddr_3_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd5_In : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd4_In : STD_LOGIC; 
  signal macaddr_5_FFX_RST : STD_LOGIC; 
  signal macaddr_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_n0048_21_Q : STD_LOGIC; 
  signal rx_input_memio_n0048_20_Q : STD_LOGIC; 
  signal memcontroller_clknum_1_2_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_1_2_GROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd12_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd11_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd14_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd13_In : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_1_GROM : STD_LOGIC; 
  signal mac_control_n0049 : STD_LOGIC; 
  signal mac_control_n0051 : STD_LOGIC; 
  signal mac_control_rxfifowerr_rst_CEMUXNOT : STD_LOGIC; 
  signal mac_control_n0047 : STD_LOGIC; 
  signal mac_control_rxf_rst_CEMUXNOT : STD_LOGIC; 
  signal macaddr_7_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_11_CEMUXNOT : STD_LOGIC; 
  signal macaddr_9_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_13_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_15_CEMUXNOT : STD_LOGIC; 
  signal tx_input_enableintl_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_enableintl_GSHIFT : STD_LOGIC; 
  signal tx_input_enableintl_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd2_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd1_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd4_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd3_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd6_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd5_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd8_In : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd7_In : STD_LOGIC; 
  signal rx_input_memio_n0049 : STD_LOGIC; 
  signal rx_input_memio_crcen_CEMUXNOT : STD_LOGIC; 
  signal tx_input_lden : STD_LOGIC; 
  signal tx_input_den_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_endfin_FROM : STD_LOGIC; 
  signal rx_input_endfin_GROM : STD_LOGIC; 
  signal rx_output_invalid_FROM : STD_LOGIC; 
  signal rx_output_fifo_N1835 : STD_LOGIC; 
  signal rx_output_fifo_N2259 : STD_LOGIC; 
  signal rx_output_fifo_N2299 : STD_LOGIC; 
  signal tx_output_n0034_1_Q : STD_LOGIC; 
  signal tx_output_n0034_0_Q : STD_LOGIC; 
  signal mac_control_lsclkdelta : STD_LOGIC; 
  signal mac_control_sclkdelta_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_n0048_1_Q : STD_LOGIC; 
  signal rx_input_memio_n0048_0_Q : STD_LOGIC; 
  signal tx_output_cs_FFd16_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd16_GROM : STD_LOGIC; 
  signal mac_control_n0050 : STD_LOGIC; 
  signal mac_control_rxphyerr_rst_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_1_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_3_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_5_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_7_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifodin_9_CEMUXNOT : STD_LOGIC; 
  signal rx_output_n0051 : STD_LOGIC; 
  signal rx_output_fifo_full_CEMUXNOT : STD_LOGIC; 
  signal rx_input_GMII_N79913 : STD_LOGIC; 
  signal rx_input_GMII_N79916 : STD_LOGIC; 
  signal rx_input_GMII_N79922 : STD_LOGIC; 
  signal rx_input_GMII_N79919 : STD_LOGIC; 
  signal rx_input_GMII_N79901 : STD_LOGIC; 
  signal rx_input_GMII_N79910 : STD_LOGIC; 
  signal rx_input_GMII_N79907 : STD_LOGIC; 
  signal rx_input_GMII_N79904 : STD_LOGIC; 
  signal tx_input_dinint_11_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_11_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_13_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_13_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_13_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_15_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_15_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_15_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_oe_FFY_RST : STD_LOGIC; 
  signal memcontroller_wen : STD_LOGIC; 
  signal rx_input_memio_n0061 : STD_LOGIC; 
  signal rx_input_memio_n0060 : STD_LOGIC; 
  signal rxfifowerr_CEMUXNOT : STD_LOGIC; 
  signal rx_output_cs_FFd17_In : STD_LOGIC; 
  signal rx_output_cs_FFd4_In : STD_LOGIC; 
  signal rx_output_cs_FFd19_In : STD_LOGIC; 
  signal mac_control_dout_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_n0058 : STD_LOGIC; 
  signal rx_input_memio_n0057 : STD_LOGIC; 
  signal rxoferr_CEMUXNOT : STD_LOGIC; 
  signal tx_input_cs_FFd11_FROM : STD_LOGIC; 
  signal tx_input_cs_FFd11_In : STD_LOGIC; 
  signal mac_control_txf_cross_GROM : STD_LOGIC; 
  signal tx_output_cs_FFd5_GROM : STD_LOGIC; 
  signal tx_output_cs_FFd6_GROM : STD_LOGIC; 
  signal tx_input_dinint_1_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_1_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_3_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_3_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_5_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_5_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_7_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_7_CEMUXNOT : STD_LOGIC; 
  signal tx_input_dinint_9_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_dinint_9_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd2_In : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd1_In : STD_LOGIC; 
  signal mac_control_PHY_status_din_3_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd2_In : STD_LOGIC; 
  signal rx_output_cs_FFd1_In : STD_LOGIC; 
  signal rx_output_cs_FFd8_In : STD_LOGIC; 
  signal rx_output_cs_FFd7_In : STD_LOGIC; 
  signal rx_input_GMII_lince : STD_LOGIC; 
  signal tx_input_cs_FFd2_In : STD_LOGIC; 
  signal tx_input_cs_FFd3_In : STD_LOGIC; 
  signal tx_input_cs_FFd10_In_O : STD_LOGIC; 
  signal tx_input_cs_FFd9_In : STD_LOGIC; 
  signal mac_control_PHY_status_din_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_10_59_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_10_net14 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_10_59_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_11_58_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_11_net12 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_11_58_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_12_57_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_12_net10 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_12_57_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_13_56_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_13_net8 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_13_56_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_14_55_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_14_net6 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_14_55_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_15_54_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_15_net4 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_15_54_CEMUXNOT : STD_LOGIC; 
  signal mac_control_Mshreg_sinlll_102_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal mac_control_Mshreg_sinlll_net185 : STD_LOGIC; 
  signal mac_control_Mshreg_sinlll_102_CEMUXNOT : STD_LOGIC; 
  signal rx_output_fifo_N2339 : STD_LOGIC; 
  signal rx_output_fifo_N2379 : STD_LOGIC; 
  signal rx_output_fifo_N2419 : STD_LOGIC; 
  signal rx_output_fifo_N2459 : STD_LOGIC; 
  signal rx_output_fifo_N3267 : STD_LOGIC; 
  signal rx_output_fifo_N3307 : STD_LOGIC; 
  signal mac_control_PHY_status_din_3_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N3187 : STD_LOGIC; 
  signal rx_output_fifo_N3227 : STD_LOGIC; 
  signal rx_output_fifo_N3347 : STD_LOGIC; 
  signal rx_output_fifo_N3387 : STD_LOGIC; 
  signal rx_output_fifo_N1589_FROM : STD_LOGIC; 
  signal rx_output_fifo_N3971 : STD_LOGIC; 
  signal rx_output_fifo_N3973 : STD_LOGIC; 
  signal rx_output_fifo_N3968 : STD_LOGIC; 
  signal rx_output_fifo_N3969 : STD_LOGIC; 
  signal tx_output_cs_FFd8_In : STD_LOGIC; 
  signal tx_output_cs_FFd7_In : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_0_69_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_0_net34 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_0_69_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_1_68_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_1_net32 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_1_68_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_2_67_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_2_net30 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_2_67_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_3_66_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_3_net28 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_3_66_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_4_65_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_4_net26 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_4_65_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_din_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_5_64_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_5_net24 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_5_64_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_6_63_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_6_net22 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_6_63_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_7_62_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_7_net20 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_7_62_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_8_61_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_8_net18 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_8_61_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_9_60_SRMUX_OUTPUTNOT : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_9_net16 : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_9_60_CEMUXNOT : STD_LOGIC; 
  signal tx_input_newfint_LOGIC_ONE : STD_LOGIC; 
  signal tx_input_lnewfint : STD_LOGIC; 
  signal tx_input_newfint_CEMUXNOT : STD_LOGIC; 
  signal tx_output_n0034_21_Q : STD_LOGIC; 
  signal tx_output_n0034_20_Q : STD_LOGIC; 
  signal mac_control_PHY_status_din_9_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_22_FROM : STD_LOGIC; 
  signal tx_output_n0034_22_Q : STD_LOGIC; 
  signal tx_output_crcl_31_FROM : STD_LOGIC; 
  signal tx_output_n0034_31_Q : STD_LOGIC; 
  signal mac_control_PHY_status_din_7_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_19_FROM : STD_LOGIC; 
  signal tx_output_n0034_19_Q : STD_LOGIC; 
  signal tx_output_crcl_13_FROM : STD_LOGIC; 
  signal tx_output_n0034_13_Q : STD_LOGIC; 
  signal rx_input_memio_crcl_6_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_6_1_O : STD_LOGIC; 
  signal tx_output_crcsell_3_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_din_9_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_3_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_30_FROM : STD_LOGIC; 
  signal tx_output_n0034_30_1_O : STD_LOGIC; 
  signal memcontroller_dnl2_5_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_7_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_9_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_14_FROM : STD_LOGIC; 
  signal tx_output_n0034_14_Q : STD_LOGIC; 
  signal mac_control_sclkdeltal_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcl_7_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_7_Q : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4_FROM : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4_In : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_5_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_9_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_21_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_23_FROM : STD_LOGIC; 
  signal tx_output_n0034_23_Q : STD_LOGIC; 
  signal rx_input_memio_crcl_10_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_10_Q : STD_LOGIC; 
  signal rx_input_memio_crcl_8_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_8_1_O : STD_LOGIC; 
  signal memcontroller_dnl2_11_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_21_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_13_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_23_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_13_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_15_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_31_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_25_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_17_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_27_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_19_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_dnl2_29_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_datal_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_datal_3_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_datal_5_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_datal_7_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_0_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_0_rt : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_0_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_0_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_2_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_2_rt : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_2_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_2_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_4_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_lmaceq_4_rt : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_4_CYINIT : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_4_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_done_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_24_FROM : STD_LOGIC; 
  signal tx_output_n0034_24_Q : STD_LOGIC; 
  signal tx_output_crcl_16_FROM : STD_LOGIC; 
  signal tx_output_n0034_16_1_O : STD_LOGIC; 
  signal rx_input_memio_crcl_11_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_11_1_O : STD_LOGIC; 
  signal mac_control_PHY_status_n0011_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_1_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_1_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_9_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_9_Q : STD_LOGIC; 
  signal mac_control_sclkdeltall_CEMUXNOT : STD_LOGIC; 
  signal mac_control_phyaddr_13_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_21_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_15_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_23_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_30_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_25_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_19_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_27_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_11_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_25_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_35_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_35_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_27_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_19_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_45_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_45_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_37_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_37_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_29_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_47_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_47_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_39_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_39_CEMUXNOT : STD_LOGIC; 
  signal mac_control_CHOICE2745_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2745_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2348_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2348_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2085_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2085_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2181_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2181_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2753_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2753_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2586_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2586_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2494_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2494_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2497_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2497_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2089_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2089_GROM : STD_LOGIC; 
  signal tx_output_crcl_28_FROM : STD_LOGIC; 
  signal tx_output_n0034_28_Q : STD_LOGIC; 
  signal mac_control_CHOICE2315_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2315_GROM : STD_LOGIC; 
  signal tx_output_crcl_8_FFY_RST : STD_LOGIC; 
  signal mac_control_CHOICE2062_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2062_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2544_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2544_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2547_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2547_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2343_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2343_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2590_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2590_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2339_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2339_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2569_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2569_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2572_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2572_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2771_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2771_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2154_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2154_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2066_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2066_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2223_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2223_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2093_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2093_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2070_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2070_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2227_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2227_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2779_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2779_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2231_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2231_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2594_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2594_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2277_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2277_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2048_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2048_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2597_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2597_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2208_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2208_GROM : STD_LOGIC; 
  signal mac_control_CHOICE2269_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2269_GROM : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_3_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_5_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_7_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_9_CEMUXNOT : STD_LOGIC; 
  signal tx_output_ltxd_3_FROM : STD_LOGIC; 
  signal tx_output_ltxd_3_GROM : STD_LOGIC; 
  signal tx_output_ltxd_5_GROM : STD_LOGIC; 
  signal tx_output_crcl_25_FROM : STD_LOGIC; 
  signal tx_output_n0034_25_Q : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_17_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_17_FROM : STD_LOGIC; 
  signal tx_output_n0034_17_Q : STD_LOGIC; 
  signal memcontroller_clknum_0_1_BYMUXNOT : STD_LOGIC; 
  signal rx_input_memio_dout_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_13_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_12_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_15_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_27_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_17_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_validbcast_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_validbcast_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_n0051 : STD_LOGIC; 
  signal rx_input_memio_addrchk_validbcast_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_bp_12_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_14_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_154_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_0_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_4_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_0_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_2_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_0_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_2_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_0_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_6_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_2_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_4_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_155_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_157_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159_FFY_RST : STD_LOGIC; 
  signal mac_control_CHOICE2273_FROM : STD_LOGIC; 
  signal mac_control_CHOICE2273_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_23_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_23_Q : STD_LOGIC; 
  signal mac_control_CHOICE2254_GROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxallfl_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_CHOICE1112_GROM : STD_LOGIC; 
  signal tx_output_crcl_29_FROM : STD_LOGIC; 
  signal tx_output_n0034_29_Q : STD_LOGIC; 
  signal rx_input_memio_crcll_11_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_13_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_21_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_15_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_31_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_23_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_17_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_25_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_27_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_19_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcll_29_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcl_24_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_24_Q : STD_LOGIC; 
  signal rx_input_memio_crcl_16_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_16_1_O : STD_LOGIC; 
  signal mac_control_N53132_FROM : STD_LOGIC; 
  signal mac_control_N53132_GROM : STD_LOGIC; 
  signal mac_control_N53204_FROM : STD_LOGIC; 
  signal mac_control_N53204_GROM : STD_LOGIC; 
  signal mac_control_N53125_FROM : STD_LOGIC; 
  signal mac_control_N53125_GROM : STD_LOGIC; 
  signal mac_control_N53118_FROM : STD_LOGIC; 
  signal mac_control_N53118_GROM : STD_LOGIC; 
  signal mac_control_N53154_FROM : STD_LOGIC; 
  signal mac_control_N53154_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_phyaddrws_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_phyaddrws_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_phyaddrws_BYMUXNOT : STD_LOGIC; 
  signal mac_control_dout_31_FROM : STD_LOGIC; 
  signal mac_control_rxcrcerr_rst_FROM : STD_LOGIC; 
  signal mac_control_n0052 : STD_LOGIC; 
  signal mac_control_rxcrcerr_rst_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE963_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE963_GROM : STD_LOGIC; 
  signal rx_input_memio_crcequal_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE980_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_CHOICE980_GROM : STD_LOGIC; 
  signal tx_output_bpl_1_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_3_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_5_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_7_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_9_CEMUXNOT : STD_LOGIC; 
  signal macaddr_13_FFY_RST : STD_LOGIC; 
  signal macaddr_21_FFY_RST : STD_LOGIC; 
  signal macaddr_31_FFY_RST : STD_LOGIC; 
  signal macaddr_23_FFY_RST : STD_LOGIC; 
  signal macaddr_15_FFY_RST : STD_LOGIC; 
  signal macaddr_33_FFY_RST : STD_LOGIC; 
  signal macaddr_41_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_4_FFY_RST : STD_LOGIC; 
  signal macaddr_25_FFY_RST : STD_LOGIC; 
  signal macaddr_17_FFY_RST : STD_LOGIC; 
  signal macaddr_27_FFY_RST : STD_LOGIC; 
  signal macaddr_35_FFY_RST : STD_LOGIC; 
  signal macaddr_19_FFY_RST : STD_LOGIC; 
  signal macaddr_29_FFY_RST : STD_LOGIC; 
  signal macaddr_37_FFY_RST : STD_LOGIC; 
  signal macaddr_45_FFY_RST : STD_LOGIC; 
  signal macaddr_39_FFY_RST : STD_LOGIC; 
  signal macaddr_47_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_addrl_1_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_addrl_4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_25_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_25_Q : STD_LOGIC; 
  signal tx_output_outsell_1_FROM : STD_LOGIC; 
  signal tx_output_outsel_1_Q : STD_LOGIC; 
  signal tx_output_outsell_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcl_17_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_17_Q : STD_LOGIC; 
  signal tx_output_outsell_0_FROM : STD_LOGIC; 
  signal tx_output_outsel_0_Q : STD_LOGIC; 
  signal tx_output_outsell_0_CEMUXNOT : STD_LOGIC; 
  signal memcontroller_oel_BYMUXNOT : STD_LOGIC; 
  signal memcontroller_oel_CEMUXNOT : STD_LOGIC; 
  signal rx_output_cs_FFd18_FROM : STD_LOGIC; 
  signal rx_output_cs_FFd18_In : STD_LOGIC; 
  signal tx_input_CHOICE2029_FROM : STD_LOGIC; 
  signal tx_input_CHOICE2029_GROM : STD_LOGIC; 
  signal tx_input_CHOICE2022_GROM : STD_LOGIC; 
  signal rx_output_fifo_nearfull_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd6_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd6_In : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd6_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd6_In : STD_LOGIC; 
  signal rx_input_memio_crccomb_Mxor_CO_26_Xo_1_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_18_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_18_Q : STD_LOGIC; 
  signal rx_input_memio_crcl_26_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_26_Q : STD_LOGIC; 
  signal memcontroller_clknum_1_BYMUXNOT : STD_LOGIC; 
  signal txfbbp_1_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_3_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_5_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_7_CEMUXNOT : STD_LOGIC; 
  signal txfbbp_9_CEMUXNOT : STD_LOGIC; 
  signal mac_control_dout_5_FFY_RST : STD_LOGIC; 
  signal addr4ext_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_3_FFY_RST : STD_LOGIC; 
  signal addr4ext_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_9_rt : STD_LOGIC; 
  signal addr4ext_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_control_d0_9_rt : STD_LOGIC; 
  signal rx_input_fifo_control_d2_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_control_d1_9_rt : STD_LOGIC; 
  signal rx_input_fifo_control_d3_9_LOGIC_ZERO : STD_LOGIC; 
  signal rx_input_fifo_control_d2_9_rt : STD_LOGIC; 
  signal addr4ext_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_27_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_27_Q : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_11_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_21_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_13_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_31_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_23_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_15_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_25_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_17_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_27_CEMUXNOT : STD_LOGIC; 
  signal addr4ext_5_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_19_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_29_CEMUXNOT : STD_LOGIC; 
  signal mac_control_PHY_status_miirw_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_miirw_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_cell_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_crcl_28_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_28_Q : STD_LOGIC; 
  signal mac_control_PHY_status_N43105_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_N43105_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_0_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_2_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_2_GROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_4_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_miiaddr_4_GROM : STD_LOGIC; 
  signal addr4ext_7_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1918_GROM : STD_LOGIC; 
  signal rx_input_memio_crcl_29_FROM : STD_LOGIC; 
  signal rx_input_memio_n0048_29_Q : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1925_GROM : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1940_GROM : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1941_FROM : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1941_GROM : STD_LOGIC; 
  signal tx_fifocheck_CHOICE1933_GROM : STD_LOGIC; 
  signal rx_input_fifo_control_celll_CEMUXNOT : STD_LOGIC; 
  signal d4_1_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_11_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_21_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_13_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_23_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_15_CEMUXNOT : STD_LOGIC; 
  signal addr4ext_9_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_31_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_17_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_25_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_19_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_27_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_29_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_cs_FFd3_FROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd3_In : STD_LOGIC; 
  signal mac_control_ledrx_rst_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_validmcast_CEMUXNOT : STD_LOGIC; 
  signal mac_control_ledtx_rst_CEMUXNOT : STD_LOGIC; 
  signal d4_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd4_FROM : STD_LOGIC; 
  signal rx_input_memio_cs_FFd4_In : STD_LOGIC; 
  signal rxallf_FFY_RST : STD_LOGIC; 
  signal d4_23_FFY_RST : STD_LOGIC; 
  signal d4_31_FFY_RST : STD_LOGIC; 
  signal d4_3_FFX_RST : STD_LOGIC; 
  signal d4_17_FFY_RST : STD_LOGIC; 
  signal d4_29_FFY_RST : STD_LOGIC; 
  signal rxfifofull_LOGIC_ONE : STD_LOGIC; 
  signal mac_control_rxf_cntl_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_5_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxf_cntl_9_CEMUXNOT : STD_LOGIC; 
  signal d4_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxbcastl_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_11_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_21_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_13_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_31_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_23_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_15_CEMUXNOT : STD_LOGIC; 
  signal d4_9_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_25_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_17_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_27_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_19_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_29_CEMUXNOT : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_1_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_5_FFY_RST : STD_LOGIC; 
  signal mac_control_CHOICE1407_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1407_GROM : STD_LOGIC; 
  signal d4_7_FFX_RST : STD_LOGIC; 
  signal mac_control_CHOICE1356_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1364_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1373_FROM : STD_LOGIC; 
  signal mac_control_CHOICE1373_GROM : STD_LOGIC; 
  signal mac_control_CHOICE1371_GROM : STD_LOGIC; 
  signal mac_control_N80967_FROM : STD_LOGIC; 
  signal mac_control_N80967_GROM : STD_LOGIC; 
  signal mac_control_n0086_FROM : STD_LOGIC; 
  signal mac_control_n0086_GROM : STD_LOGIC; 
  signal d4_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxmcastl_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_1_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_3_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_5_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_7_CEMUXNOT : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_9_CEMUXNOT : STD_LOGIC; 
  signal mac_control_n00851_1_FROM : STD_LOGIC; 
  signal mac_control_n00851_1_GROM : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxucastl_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd1_FROM : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd1_In : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_13_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_15_FFX_RST : STD_LOGIC; 
  signal rxbp_11_CEMUXNOT : STD_LOGIC; 
  signal rxbp_13_CEMUXNOT : STD_LOGIC; 
  signal rxbp_15_CEMUXNOT : STD_LOGIC; 
  signal rx_output_cs_FFd12_FFX_RST : STD_LOGIC; 
  signal rx_output_ceinl_FFX_RST : STD_LOGIC; 
  signal tx_output_N80951_GROM : STD_LOGIC; 
  signal tx_output_bpl_11_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_13_CEMUXNOT : STD_LOGIC; 
  signal tx_output_bpl_15_CEMUXNOT : STD_LOGIC; 
  signal rx_output_cs_FFd14_FFX_RST : STD_LOGIC; 
  signal tx_output_outsell_2_FROM : STD_LOGIC; 
  signal tx_output_outsel_3_Q : STD_LOGIC; 
  signal tx_output_outsell_2_CEMUXNOT : STD_LOGIC; 
  signal rx_input_memio_fifofulll_CEMUXNOT : STD_LOGIC; 
  signal rx_output_nfl_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_1_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_3_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_5_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_7_CEMUXNOT : STD_LOGIC; 
  signal mac_control_txf_cntl_9_CEMUXNOT : STD_LOGIC; 
  signal rx_output_cs_FFd16_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81171_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81171_GROM : STD_LOGIC; 
  signal tx_output_crcl_3_FROM : STD_LOGIC; 
  signal tx_output_n0034_3_Q : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81405_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81405_GROM : STD_LOGIC; 
  signal mac_control_dout_6_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_RESET_1_GROM : STD_LOGIC; 
  signal rxf_CEMUXNOT : STD_LOGIC; 
  signal tx_output_crcl_4_FROM : STD_LOGIC; 
  signal tx_output_n0034_4_1_O : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81167_FROM : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_N81167_GROM : STD_LOGIC; 
  signal mac_control_dout_7_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cross_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_5_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_7_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_2_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd14_FFX_RST : STD_LOGIC; 
  signal tx_output_data_2_FFY_RST : STD_LOGIC; 
  signal tx_output_data_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd7_FFX_SET : STD_LOGIC; 
  signal tx_output_data_6_FFY_RST : STD_LOGIC; 
  signal tx_output_data_7_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_2_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_2_FFX_RST : STD_LOGIC; 
  signal tx_output_bcntl_4_FFX_RST : STD_LOGIC; 
  signal tx_output_bcntl_6_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_11_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_13_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_15_FFX_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_1_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_2_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_3_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_8_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_1_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_1_FFX_RST : STD_LOGIC; 
  signal tx_input_dh_3_FFX_RST : STD_LOGIC; 
  signal tx_input_dh_5_FFX_RST : STD_LOGIC; 
  signal tx_input_dh_7_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_7_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_1_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_9_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_9_FFX_RST : STD_LOGIC; 
  signal txbp_9_FFY_RST : STD_LOGIC; 
  signal txbp_9_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_1_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_1_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_3_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_5_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_7_FFX_RST : STD_LOGIC; 
  signal rxbp_1_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_9_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_15_FFX_RST : STD_LOGIC; 
  signal tx_output_ltxen3_FFY_RST : STD_LOGIC; 
  signal tx_output_ltxen3_FFX_RST : STD_LOGIC; 
  signal tx_input_DONE_FFY_RST : STD_LOGIC; 
  signal MD_13_OFF_RST : STD_LOGIC; 
  signal MD_22_IFF_RST : STD_LOGIC; 
  signal MD_22_OFF_RST : STD_LOGIC; 
  signal MD_14_IFF_RST : STD_LOGIC; 
  signal MD_14_OFF_RST : STD_LOGIC; 
  signal MD_30_IFF_RST : STD_LOGIC; 
  signal MD_23_IFF_RST : STD_LOGIC; 
  signal MD_30_OFF_RST : STD_LOGIC; 
  signal tx_input_dl_1_FFX_RST : STD_LOGIC; 
  signal txbp_1_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_3_FFX_RST : STD_LOGIC; 
  signal txbp_3_FFY_RST : STD_LOGIC; 
  signal txbp_3_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_5_FFX_RST : STD_LOGIC; 
  signal txbp_5_FFY_RST : STD_LOGIC; 
  signal txbp_5_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_7_FFX_RST : STD_LOGIC; 
  signal txbp_7_FFY_RST : STD_LOGIC; 
  signal txbp_7_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_0_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_25_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_17_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_27_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_19_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_29_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_10_FFY_RST : STD_LOGIC; 
  signal DOUT_3_OFF_RST : STD_LOGIC; 
  signal DOUT_4_OFF_RST : STD_LOGIC; 
  signal DOUT_5_OFF_RST : STD_LOGIC; 
  signal DOUT_6_OFF_RST : STD_LOGIC; 
  signal DOUT_7_OFF_RST : STD_LOGIC; 
  signal tx_output_outselll_1_FFX_RST : STD_LOGIC; 
  signal tx_output_outselll_1_FFY_SET : STD_LOGIC; 
  signal tx_output_outselll_3_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_11_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_11_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_21_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_13_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_11_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_21_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_13_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_31_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_23_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_25_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_15_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1603_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N1607_FFX_SET : STD_LOGIC; 
  signal mac_control_phystat_25_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_17_FFX_RST : STD_LOGIC; 
  signal q3_31_FFX_RST : STD_LOGIC; 
  signal q3_15_FFY_RST : STD_LOGIC; 
  signal q3_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_mcast_0_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_0_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_11_FFY_RST : STD_LOGIC; 
  signal addr2ext_4_FFX_RST : STD_LOGIC; 
  signal addr2ext_6_FFX_RST : STD_LOGIC; 
  signal addr2ext_8_FFY_RST : STD_LOGIC; 
  signal addr2ext_10_FFY_RST : STD_LOGIC; 
  signal addr2ext_12_FFY_RST : STD_LOGIC; 
  signal addr2ext_14_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_87_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_89_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_91_FFY_RST : STD_LOGIC; 
  signal tx_output_data_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_3_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_5_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_7_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_7_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_11_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_13_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_13_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_15_FFY_RST : STD_LOGIC; 
  signal rxucast_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_11_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_12_FFX_RST : STD_LOGIC; 
  signal tx_output_crcsell_0_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_1_FFY_RST : STD_LOGIC; 
  signal tx_output_crcsell_0_FFX_SET : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_1_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd15_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd12_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd14_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_4_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_5_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_6_FFY_RST : STD_LOGIC; 
  signal tx_output_ncrcbytel_7_FFY_RST : STD_LOGIC; 
  signal rxmcast_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_11_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_21_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_13_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_31_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_23_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_15_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_25_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_25_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_17_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_27_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_19_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_29_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_1_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_fbbpl_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd8_FFX_RST : STD_LOGIC; 
  signal mac_control_bitcnt_109_FFX_RST : STD_LOGIC; 
  signal tx_output_data_4_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_12_FFY_RST : STD_LOGIC; 
  signal tx_output_bcntl_12_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_0_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_bcast_2_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_13_FFY_RST : STD_LOGIC; 
  signal mac_control_Mshreg_scslll_103_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_11_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_3_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_5_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_7_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_rwl_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_2_FFY_RST : STD_LOGIC; 
  signal TXD_4_OFF_RST : STD_LOGIC; 
  signal TXD_5_OFF_RST : STD_LOGIC; 
  signal TXD_6_OFF_RST : STD_LOGIC; 
  signal TXD_7_OFF_RST : STD_LOGIC; 
  signal LEDDPX_OFF_RST : STD_LOGIC; 
  signal rxfbbp_1_FFX_RST : STD_LOGIC; 
  signal tx_output_bcntl_8_FFX_RST : STD_LOGIC; 
  signal rxfbbp_3_FFX_RST : STD_LOGIC; 
  signal tx_output_datal_1_FFX_RST : STD_LOGIC; 
  signal tx_output_bcntl_10_FFX_RST : STD_LOGIC; 
  signal rxfbbp_5_FFX_RST : STD_LOGIC; 
  signal tx_output_datal_3_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1610_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N1563_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1627_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1567_FFX_RST : STD_LOGIC; 
  signal q2_11_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1627_FFX_RST : STD_LOGIC; 
  signal q2_11_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1569_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1565_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1605_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N1609_FFX_SET : STD_LOGIC; 
  signal mac_control_phystat_21_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_13_FFX_RST : STD_LOGIC; 
  signal q2_27_FFX_RST : STD_LOGIC; 
  signal q2_19_FFX_RST : STD_LOGIC; 
  signal q3_11_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1585_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_79_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_81_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_83_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_85_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1579_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1579_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1583_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1583_FFX_RST : STD_LOGIC; 
  signal q3_23_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_27_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_27_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_19_FFX_RST : STD_LOGIC; 
  signal q3_25_FFX_RST : STD_LOGIC; 
  signal q3_17_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_29_FFX_RST : STD_LOGIC; 
  signal rxfbbp_7_FFX_RST : STD_LOGIC; 
  signal tx_output_datal_5_FFX_RST : STD_LOGIC; 
  signal rxfbbp_9_FFX_RST : STD_LOGIC; 
  signal rxfbbp_9_FFY_RST : STD_LOGIC; 
  signal tx_output_datal_7_FFX_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_3_FFX_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_5_FFY_RST : STD_LOGIC; 
  signal q3_27_FFX_RST : STD_LOGIC; 
  signal q3_19_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1581_FFX_RST : STD_LOGIC; 
  signal q3_29_FFX_RST : STD_LOGIC; 
  signal rx_output_ceinll_FFY_RST : STD_LOGIC; 
  signal tx_output_data_5_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd3_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_23_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_31_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_15_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1571_FFX_RST : STD_LOGIC; 
  signal q2_29_FFX_RST : STD_LOGIC; 
  signal q3_21_FFX_RST : STD_LOGIC; 
  signal q3_13_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1586_FFX_SET : STD_LOGIC; 
  signal LEDACT_OFF_RST : STD_LOGIC; 
  signal TXD_0_OFF_RST : STD_LOGIC; 
  signal TXD_1_OFF_RST : STD_LOGIC; 
  signal TXD_2_OFF_RST : STD_LOGIC; 
  signal TXD_3_OFF_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_31_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_23_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_15_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_25_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_27_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_17_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_19_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_27_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_27_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_19_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_29_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd10_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd3_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd10_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_3_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_19_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_29_FFX_RST : STD_LOGIC; 
  signal MDIO_IFF_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_37_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_10_FFY_RST : STD_LOGIC; 
  signal rx_output_len_11_FFY_RST : STD_LOGIC; 
  signal rx_output_len_11_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_11_FFX_RST : STD_LOGIC; 
  signal rx_output_len_13_FFY_RST : STD_LOGIC; 
  signal rx_output_len_13_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_21_FFX_RST : STD_LOGIC; 
  signal LED1000_OFF_RST : STD_LOGIC; 
  signal TX_EN_OFF_RST : STD_LOGIC; 
  signal DOUTEN_OFF_RST : STD_LOGIC; 
  signal MWE_OFF_SET : STD_LOGIC; 
  signal NEXTFRAME_IFF_RST : STD_LOGIC; 
  signal rx_output_mdl_13_FFX_RST : STD_LOGIC; 
  signal rx_output_len_15_FFY_RST : STD_LOGIC; 
  signal rx_output_len_15_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_31_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_23_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_15_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_25_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_25_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_17_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_7_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_27_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_19_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_8_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_28_FFX_RST : STD_LOGIC; 
  signal DOUT_10_OFF_RST : STD_LOGIC; 
  signal DOUT_11_OFF_RST : STD_LOGIC; 
  signal DOUT_12_OFF_RST : STD_LOGIC; 
  signal DOUT_13_OFF_RST : STD_LOGIC; 
  signal DOUT_14_OFF_RST : STD_LOGIC; 
  signal rx_output_len_5_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_5_FFX_RST : STD_LOGIC; 
  signal rx_output_len_7_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_7_FFX_RST : STD_LOGIC; 
  signal rx_output_len_9_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_4_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_5_FFX_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_7_FFX_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_cntl_9_FFX_RST : STD_LOGIC; 
  signal rx_output_len_1_FFY_RST : STD_LOGIC; 
  signal rx_output_len_1_FFX_RST : STD_LOGIC; 
  signal rx_output_mdl_1_FFX_RST : STD_LOGIC; 
  signal rx_output_len_3_FFX_RST : STD_LOGIC; 
  signal rx_output_len_5_FFY_RST : STD_LOGIC; 
  signal rx_output_mdl_3_FFX_RST : STD_LOGIC; 
  signal DOUT_15_OFF_RST : STD_LOGIC; 
  signal LED100_OFF_RST : STD_LOGIC; 
  signal NEWFRAME_IFF_RST : STD_LOGIC; 
  signal MD_28_OFF_RST : STD_LOGIC; 
  signal MD_29_IFF_RST : STD_LOGIC; 
  signal MD_29_OFF_RST : STD_LOGIC; 
  signal MA_0_OFF_RST : STD_LOGIC; 
  signal MA_1_OFF_RST : STD_LOGIC; 
  signal MA_2_OFF_RST : STD_LOGIC; 
  signal MD_23_OFF_RST : STD_LOGIC; 
  signal MD_15_IFF_RST : STD_LOGIC; 
  signal MD_15_OFF_RST : STD_LOGIC; 
  signal MD_31_IFF_RST : STD_LOGIC; 
  signal MD_31_OFF_RST : STD_LOGIC; 
  signal MD_24_IFF_RST : STD_LOGIC; 
  signal MA_3_OFF_RST : STD_LOGIC; 
  signal MA_4_OFF_RST : STD_LOGIC; 
  signal MA_5_OFF_RST : STD_LOGIC; 
  signal MA_6_OFF_RST : STD_LOGIC; 
  signal MA_7_OFF_RST : STD_LOGIC; 
  signal MD_18_OFF_RST : STD_LOGIC; 
  signal MD_26_IFF_RST : STD_LOGIC; 
  signal MD_26_OFF_RST : STD_LOGIC; 
  signal MD_19_IFF_RST : STD_LOGIC; 
  signal MD_19_OFF_RST : STD_LOGIC; 
  signal MD_27_IFF_RST : STD_LOGIC; 
  signal MD_28_IFF_RST : STD_LOGIC; 
  signal MD_27_OFF_RST : STD_LOGIC; 
  signal RXD_0_IFF_RST : STD_LOGIC; 
  signal RXD_1_IFF_RST : STD_LOGIC; 
  signal RXD_2_IFF_RST : STD_LOGIC; 
  signal RXD_3_IFF_RST : STD_LOGIC; 
  signal RXD_4_IFF_RST : STD_LOGIC; 
  signal RXD_5_IFF_RST : STD_LOGIC; 
  signal RXD_6_IFF_RST : STD_LOGIC; 
  signal RXD_7_IFF_RST : STD_LOGIC; 
  signal DIN_10_IFF_RST : STD_LOGIC; 
  signal DIN_11_IFF_RST : STD_LOGIC; 
  signal DIN_12_IFF_RST : STD_LOGIC; 
  signal DIN_13_IFF_RST : STD_LOGIC; 
  signal DIN_14_IFF_RST : STD_LOGIC; 
  signal DIN_15_IFF_RST : STD_LOGIC; 
  signal DOUT_0_OFF_RST : STD_LOGIC; 
  signal DOUT_1_OFF_RST : STD_LOGIC; 
  signal DOUT_2_OFF_RST : STD_LOGIC; 
  signal DIN_8_IFF_RST : STD_LOGIC; 
  signal DIN_9_IFF_RST : STD_LOGIC; 
  signal RX_ER_IFF_RST : STD_LOGIC; 
  signal RX_DV_IFF_RST : STD_LOGIC; 
  signal MA_10_OFF_RST : STD_LOGIC; 
  signal MA_11_OFF_RST : STD_LOGIC; 
  signal MA_12_OFF_RST : STD_LOGIC; 
  signal MA_13_OFF_RST : STD_LOGIC; 
  signal DOUT_8_OFF_RST : STD_LOGIC; 
  signal DOUT_9_OFF_RST : STD_LOGIC; 
  signal SOUT_OFF_RST : STD_LOGIC; 
  signal SCLK_IFF_RST : STD_LOGIC; 
  signal LEDRX_OFF_RST : STD_LOGIC; 
  signal MA_14_OFF_RST : STD_LOGIC; 
  signal MA_15_OFF_RST : STD_LOGIC; 
  signal MA_16_OFF_RST : STD_LOGIC; 
  signal MD_10_IFF_RST : STD_LOGIC; 
  signal MD_10_OFF_RST : STD_LOGIC; 
  signal MD_11_IFF_RST : STD_LOGIC; 
  signal LEDTX_OFF_RST : STD_LOGIC; 
  signal DIN_0_IFF_RST : STD_LOGIC; 
  signal DIN_1_IFF_RST : STD_LOGIC; 
  signal DIN_2_IFF_RST : STD_LOGIC; 
  signal DIN_3_IFF_RST : STD_LOGIC; 
  signal DIN_4_IFF_RST : STD_LOGIC; 
  signal DIN_5_IFF_RST : STD_LOGIC; 
  signal DIN_6_IFF_RST : STD_LOGIC; 
  signal DIN_7_IFF_RST : STD_LOGIC; 
  signal MD_9_OFF_RST : STD_LOGIC; 
  signal mac_control_dout_30_FFX_RST : STD_LOGIC; 
  signal MD_1_OFF_RST : STD_LOGIC; 
  signal MD_2_IFF_RST : STD_LOGIC; 
  signal MD_2_OFF_RST : STD_LOGIC; 
  signal MD_3_IFF_RST : STD_LOGIC; 
  signal MD_3_OFF_RST : STD_LOGIC; 
  signal MD_4_IFF_RST : STD_LOGIC; 
  signal MD_5_IFF_RST : STD_LOGIC; 
  signal MD_4_OFF_RST : STD_LOGIC; 
  signal MA_8_OFF_RST : STD_LOGIC; 
  signal MA_9_OFF_RST : STD_LOGIC; 
  signal PHYRESET_OFF_RST : STD_LOGIC; 
  signal MD_0_IFF_RST : STD_LOGIC; 
  signal MD_0_OFF_RST : STD_LOGIC; 
  signal MD_1_IFF_RST : STD_LOGIC; 
  signal MD_16_IFF_RST : STD_LOGIC; 
  signal MD_24_OFF_RST : STD_LOGIC; 
  signal MD_16_OFF_RST : STD_LOGIC; 
  signal MD_17_IFF_RST : STD_LOGIC; 
  signal MD_17_OFF_RST : STD_LOGIC; 
  signal MD_25_IFF_RST : STD_LOGIC; 
  signal MD_25_OFF_RST : STD_LOGIC; 
  signal MD_18_IFF_RST : STD_LOGIC; 
  signal MD_11_OFF_RST : STD_LOGIC; 
  signal MD_20_IFF_RST : STD_LOGIC; 
  signal MD_20_OFF_RST : STD_LOGIC; 
  signal MD_12_IFF_RST : STD_LOGIC; 
  signal MD_12_OFF_RST : STD_LOGIC; 
  signal MD_21_IFF_RST : STD_LOGIC; 
  signal MD_13_IFF_RST : STD_LOGIC; 
  signal MD_21_OFF_RST : STD_LOGIC; 
  signal addr2ext_8_FFX_RST : STD_LOGIC; 
  signal addr2ext_10_FFX_RST : STD_LOGIC; 
  signal addr2ext_12_FFX_RST : STD_LOGIC; 
  signal addr2ext_14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_86_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_21_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_22_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_23_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_20_FFX_RST : STD_LOGIC; 
  signal MD_5_OFF_RST : STD_LOGIC; 
  signal MD_6_IFF_RST : STD_LOGIC; 
  signal MD_6_OFF_RST : STD_LOGIC; 
  signal MD_7_IFF_RST : STD_LOGIC; 
  signal MD_7_OFF_RST : STD_LOGIC; 
  signal MD_8_IFF_RST : STD_LOGIC; 
  signal MD_9_IFF_RST : STD_LOGIC; 
  signal MD_8_OFF_RST : STD_LOGIC; 
  signal memcontroller_dnl1_20_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_2_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_21_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_13_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_30_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_16_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_24_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_25_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_17_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_10_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_1_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_11_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_0_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_12_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_25_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_17_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_6_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_26_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_18_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_22_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_14_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_31_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_15_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_23_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_18_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_26_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_19_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_27_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_28_FFX_RST : STD_LOGIC; 
  signal mac_control_dout_29_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_3_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_4_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_24_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_16_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_47_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_3_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_1_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_5_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_3_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_7_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_9_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_9_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_7_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_7_FFX_RST : STD_LOGIC; 
  signal mac_control_phystat_9_FFY_RST : STD_LOGIC; 
  signal mac_control_phystat_9_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_25_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_17_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_0_1_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_1_3_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_29_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_5_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_7_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_8_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d0_9_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_control_d0_9_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_5_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_1_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_1_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_3_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_3_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_5_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_5_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_7_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_7_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_9_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_9_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_13_FFY_RST : STD_LOGIC; 
  signal addr2ext_0_FFY_RST : STD_LOGIC; 
  signal addr2ext_2_FFY_RST : STD_LOGIC; 
  signal addr2ext_6_FFY_RST : STD_LOGIC; 
  signal addr2ext_0_FFX_RST : STD_LOGIC; 
  signal addr2ext_2_FFX_RST : STD_LOGIC; 
  signal addr2ext_4_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_89_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_91_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_93_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_93_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_95_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_97_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl1_9_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl1_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_6_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_8_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_10_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_0_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_95_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_97_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_99_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_101_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_99_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_0_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_2_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bp_4_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_165_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_159_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_161_FFX_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_cnt_163_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N17_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_151_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_153_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_10_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_12_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_14_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_4_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_6_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_8_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_39_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_39_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_41_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_45_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_41_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_43_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_8_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_10_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_12_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_0_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_12_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_14_FFY_RST : STD_LOGIC; 
  signal addr3ext_1_FFY_RST : STD_LOGIC; 
  signal addr3ext_0_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_117_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_119_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_121_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_125_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_121_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_123_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_10_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_12_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_14_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_14_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_38_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_43_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_45_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_47_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_51_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_47_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_49_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_4_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_6_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_8_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_12_FFY_RST : STD_LOGIC; 
  signal rx_output_bp_8_FFX_RST : STD_LOGIC; 
  signal rx_output_bp_10_FFY_RST : STD_LOGIC; 
  signal tx_output_bcnt_49_FFX_RST : STD_LOGIC; 
  signal tx_output_bcnt_51_FFX_RST : STD_LOGIC; 
  signal addr3ext_7_FFX_RST : STD_LOGIC; 
  signal addr3ext_9_FFY_RST : STD_LOGIC; 
  signal addr3ext_9_FFX_RST : STD_LOGIC; 
  signal addr3ext_11_FFY_RST : STD_LOGIC; 
  signal addr3ext_13_FFY_RST : STD_LOGIC; 
  signal addr3ext_11_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_2_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_4_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_6_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_10_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_6_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_8_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N13_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N11_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_diff_14_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_0_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_diff_2_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_32_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_129_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_131_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_133_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_133_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_135_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_33_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_mdccnt_35_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_143_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_149_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_145_FFX_RST : STD_LOGIC; 
  signal mac_control_ledtx_cnt_147_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N17_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N15_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N15_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N13_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N11_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_139_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_70_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_77_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_71_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_73_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_75_FFY_RST : STD_LOGIC; 
  signal tx_input_addr_17_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_19_FFY_RST : STD_LOGIC; 
  signal tx_input_addr_19_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_21_FFY_RST : STD_LOGIC; 
  signal tx_input_addr_23_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_111_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_110_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_113_FFY_RST : STD_LOGIC; 
  signal addr3ext_1_FFX_RST : STD_LOGIC; 
  signal addr3ext_3_FFY_RST : STD_LOGIC; 
  signal addr3ext_3_FFX_RST : STD_LOGIC; 
  signal addr3ext_5_FFY_RST : STD_LOGIC; 
  signal addr3ext_7_FFY_RST : STD_LOGIC; 
  signal addr3ext_5_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_123_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_125_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_127_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_131_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_127_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_129_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_0_FFY_RST : STD_LOGIC; 
  signal addr3ext_13_FFX_RST : STD_LOGIC; 
  signal addr3ext_15_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_135_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_137_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_137_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_139_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_141_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_111_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_113_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_115_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_119_FFY_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_115_FFX_RST : STD_LOGIC; 
  signal mac_control_phyrstcnt_117_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_73_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_83_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_75_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_77_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_79_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_81_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_6_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_8_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_21_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_23_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_25_FFY_RST : STD_LOGIC; 
  signal tx_input_addr_25_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_27_FFY_RST : STD_LOGIC; 
  signal tx_input_addr_29_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_rst_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd4_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd10_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd10_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_1_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_3_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_1_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_3_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_5_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_statecnt_5_FFX_RST : STD_LOGIC; 
  signal addr1ext_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_0_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_2_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_4_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_27_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_29_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_10_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_12_FFX_RST : STD_LOGIC; 
  signal tx_input_addr_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcntl_14_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N5_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N3_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_empty_FFX_SET : STD_LOGIC; 
  signal rx_input_endf_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_15_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_15_FFY_RST : STD_LOGIC; 
  signal rx_input_endf_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_22_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_22_FFX_RST : STD_LOGIC; 
  signal rx_output_lenr_10_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_menl_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_2_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_3_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_4_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_5_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_6_FFY_RST : STD_LOGIC; 
  signal tx_output_crcenl_FFX_RST : STD_LOGIC; 
  signal mac_control_bitcnt_105_FFY_RST : STD_LOGIC; 
  signal mac_control_bitcnt_105_FFX_RST : STD_LOGIC; 
  signal mac_control_bitcnt_107_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_15_FFY_RST : STD_LOGIC; 
  signal mac_control_bitcnt_107_FFX_RST : STD_LOGIC; 
  signal d1_11_FFX_RST : STD_LOGIC; 
  signal d1_21_FFX_RST : STD_LOGIC; 
  signal d1_21_FFY_RST : STD_LOGIC; 
  signal d1_13_FFY_RST : STD_LOGIC; 
  signal d1_13_FFX_RST : STD_LOGIC; 
  signal d1_31_FFX_RST : STD_LOGIC; 
  signal d1_31_FFY_RST : STD_LOGIC; 
  signal d1_23_FFY_RST : STD_LOGIC; 
  signal d1_23_FFX_RST : STD_LOGIC; 
  signal d1_25_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N9_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N9_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N7_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N7_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N5_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N3_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_full_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_wrcount_0_FFY_RST : STD_LOGIC; 
  signal mac_control_bitcnt_104_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_wrcount_0_FFX_RST : STD_LOGIC; 
  signal rx_output_lenr_11_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_12_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_13_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_14_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_15_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd6_FFX_RST : STD_LOGIC; 
  signal tx_input_cs_FFd8_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_rd_en_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_31_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_rst_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal addr1ext_3_FFX_RST : STD_LOGIC; 
  signal addr1ext_1_FFX_RST : STD_LOGIC; 
  signal addr1ext_3_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd5_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd5_FFY_RST : STD_LOGIC; 
  signal addr1ext_5_FFY_RST : STD_LOGIC; 
  signal addr1ext_7_FFX_RST : STD_LOGIC; 
  signal addr1ext_5_FFX_RST : STD_LOGIC; 
  signal addr1ext_7_FFY_RST : STD_LOGIC; 
  signal addr1ext_9_FFY_RST : STD_LOGIC; 
  signal d1_15_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_1_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_3_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_5_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_5_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_7_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_7_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_9_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_9_FFY_RST : STD_LOGIC; 
  signal rx_input_endfin_FFY_RST : STD_LOGIC; 
  signal rx_output_invalid_FFY_RST : STD_LOGIC; 
  signal addr1ext_9_FFX_RST : STD_LOGIC; 
  signal d1_15_FFX_RST : STD_LOGIC; 
  signal d1_14_FFX_RST : STD_LOGIC; 
  signal d1_14_FFY_RST : STD_LOGIC; 
  signal d1_3_FFX_RST : STD_LOGIC; 
  signal d1_3_FFY_RST : STD_LOGIC; 
  signal d1_5_FFX_RST : STD_LOGIC; 
  signal d1_5_FFY_RST : STD_LOGIC; 
  signal d1_7_FFX_RST : STD_LOGIC; 
  signal d1_7_FFY_RST : STD_LOGIC; 
  signal d1_9_FFY_RST : STD_LOGIC; 
  signal mac_control_rxfifowerr_rst_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_1_FFX_SET : STD_LOGIC; 
  signal addr1ext_11_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_rst_FFY_RST : STD_LOGIC; 
  signal addr1ext_11_FFX_RST : STD_LOGIC; 
  signal addr1ext_13_FFX_RST : STD_LOGIC; 
  signal addr1ext_13_FFY_RST : STD_LOGIC; 
  signal addr1ext_15_FFX_RST : STD_LOGIC; 
  signal addr1ext_15_FFY_RST : STD_LOGIC; 
  signal d1_11_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1553_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_1_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1553_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_1_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_sclkdelta_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_rst_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_1_FFX_RST : STD_LOGIC; 
  signal rx_output_lenr_7_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_8_FFY_RST : STD_LOGIC; 
  signal rx_output_lenr_9_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_9_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_full_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_11_FFY_RST : STD_LOGIC; 
  signal d1_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd12_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_1_2_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd12_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd14_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd14_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_1_FFY_SET : STD_LOGIC; 
  signal mac_control_rxfifowerr_rst_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_11_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_13_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_15_FFX_RST : STD_LOGIC; 
  signal rxfifowerr_FFY_RST : STD_LOGIC; 
  signal rxfifowerr_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd17_FFY_RST : STD_LOGIC; 
  signal d1_25_FFX_RST : STD_LOGIC; 
  signal d1_17_FFY_RST : STD_LOGIC; 
  signal d1_17_FFX_RST : STD_LOGIC; 
  signal d1_27_FFY_RST : STD_LOGIC; 
  signal d1_27_FFX_RST : STD_LOGIC; 
  signal d1_19_FFY_RST : STD_LOGIC; 
  signal d1_19_FFX_RST : STD_LOGIC; 
  signal d1_29_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_11_FFY_RST : STD_LOGIC; 
  signal d1_29_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd16_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_1_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_1_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_3_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_3_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_5_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_5_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_7_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_7_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_7_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_7_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd6_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bcnt_88_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_10_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_3_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_1_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_11_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_13_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_13_FFX_RST : STD_LOGIC; 
  signal rx_output_fifodin_15_FFY_RST : STD_LOGIC; 
  signal rx_output_fifodin_15_FFX_RST : STD_LOGIC; 
  signal tx_input_enableintl_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd4_FFY_SET : STD_LOGIC; 
  signal rx_output_cs_FFd4_FFX_RST : STD_LOGIC; 
  signal rxoferr_FFY_RST : STD_LOGIC; 
  signal rxoferr_FFX_RST : STD_LOGIC; 
  signal tx_input_cs_FFd11_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cross_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_11_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_11_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_13_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_13_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_15_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd4_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd6_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_cs_FFd8_FFX_SET : STD_LOGIC; 
  signal rx_input_memio_crcen_FFY_RST : STD_LOGIC; 
  signal tx_input_den_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_1_FFY_RST : STD_LOGIC; 
  signal tx_input_CNT_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_7_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_wbpl_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_13_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_27_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_30_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_5_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_7_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_7_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_9_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_9_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal rx_output_cs_FFd2_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd2_FFX_RST : STD_LOGIC; 
  signal tx_input_CNT_15_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd5_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_1_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal tx_output_cs_FFd5_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd6_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_1_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_3_FFY_RST : STD_LOGIC; 
  signal tx_input_dinint_3_FFX_RST : STD_LOGIC; 
  signal tx_input_dinint_5_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd8_FFX_RST : STD_LOGIC; 
  signal rx_input_ince_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd4_FFX_RST : STD_LOGIC; 
  signal txfifowerr_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd10_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd10_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_10_59_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_11_58_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1589_FFX_SET : STD_LOGIC; 
  signal rx_output_fifo_N1593_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1593_FFX_SET : STD_LOGIC; 
  signal tx_output_cs_FFd8_FFX_RST : STD_LOGIC; 
  signal tx_output_cs_FFd8_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_0_69_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_1_68_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_2_67_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_3_66_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_9_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_13_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_6_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_11_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_11_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_13_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_13_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_15_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_15_FFX_RST : STD_LOGIC; 
  signal tx_output_crcsell_3_FFY_RST : STD_LOGIC; 
  signal tx_output_crcsell_3_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_1_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1549_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1615_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1617_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1617_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1613_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1613_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1589_FFY_SET : STD_LOGIC; 
  signal rx_output_fifo_N1588_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_12_57_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_13_56_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_14_55_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_15_54_FFY_RST : STD_LOGIC; 
  signal mac_control_Mshreg_sinlll_102_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1551_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1551_FFX_RST : STD_LOGIC; 
  signal rx_output_fifo_N1615_FFY_RST : STD_LOGIC; 
  signal rx_output_fifo_N1549_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_1_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_3_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_3_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_30_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_5_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_5_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_7_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_7_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_9_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_9_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_14_FFY_RST : STD_LOGIC; 
  signal mac_control_sclkdeltal_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_4_65_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_5_64_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_6_63_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_7_62_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_8_61_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_Mshreg_lbpout4_9_60_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_21_FFY_RST : STD_LOGIC; 
  signal tx_input_newfint_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_21_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_22_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_31_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_1_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_1_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_3_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_3_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_5_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_5_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_7_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_7_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_bpl_9_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_23_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_15_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_14_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_17_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_27_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_7_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_cs_FFd4_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_9_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_1_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_15_FFX_RST : STD_LOGIC; 
  signal txbp_15_FFY_RST : STD_LOGIC; 
  signal txbp_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxucastl_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd1_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_11_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_11_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_13_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_21_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_21_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_13_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_23_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_23_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_27_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_35_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_35_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_43_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_43_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_37_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_37_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_45_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_45_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_39_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_39_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_47_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_1_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_3_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_3_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_5_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_5_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_7_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_7_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_9_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_1_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_3_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_3_FFX_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd1_FFY_RST : STD_LOGIC; 
  signal mac_control_txfifowerr_cntl_5_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_1_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_3_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_5_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_5_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_7_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_7_FFX_RST : STD_LOGIC; 
  signal mac_control_phydo_9_FFY_RST : STD_LOGIC; 
  signal mac_control_phydo_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_8_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_11_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_11_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_21_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_21_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_13_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_19_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_29_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_datal_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_datal_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_datal_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_datal_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_datal_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_datal_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_datal_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_datal_7_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_0_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_0_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_13_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_23_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_23_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_15_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_15_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_31_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_31_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_25_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_25_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_17_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_17_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_27_FFY_RST : STD_LOGIC; 
  signal memcontroller_dnl2_27_FFX_RST : STD_LOGIC; 
  signal memcontroller_dnl2_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_sclkdeltall_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_11_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_11_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_13_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_21_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_23_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_23_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_41_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_33_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_33_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_41_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_17_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_2_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_maceq_4_FFX_RST : STD_LOGIC; 
  signal tx_output_crcl_24_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_16_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_11_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_11_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_13_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_13_FFX_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_15_FFY_RST : STD_LOGIC; 
  signal rx_fifocheck_fbbpl_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_13_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_dreg_12_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_dout_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_dout_31_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_17_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_23_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_17_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_25_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_19_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_27_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_13_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_datal_21_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_3_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_5_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_5_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_7_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_7_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_9_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_9_FFX_RST : STD_LOGIC; 
  signal macaddr_11_FFY_RST : STD_LOGIC; 
  signal macaddr_11_FFX_RST : STD_LOGIC; 
  signal macaddr_13_FFX_RST : STD_LOGIC; 
  signal macaddr_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_45_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_37_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_47_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_39_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_1_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_validucast_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_3_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_3_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_5_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_5_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_7_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_7_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_9_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpen_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_destok_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd10_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_18_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_26_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_5_FFY_RST : STD_LOGIC; 
  signal mac_control_lrxallf_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_doutl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_14_FFY_RST : STD_LOGIC; 
  signal tx_input_cs_FFd12_FFY_SET : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_1_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_3_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_3_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_5_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_5_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_7_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_7_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_23_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_41_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_phyaddrws_FFY_RST : STD_LOGIC; 
  signal mac_control_dout_31_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_rst_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_1_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_3_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_41_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_33_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_17_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_43_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_35_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_27_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_macaddrl_19_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_28_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxallfl_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_23_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_17_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_25_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_addrl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_addrl_3_FFX_RST : STD_LOGIC; 
  signal tx_output_outsell_1_FFY_RST : STD_LOGIC; 
  signal mac_control_din_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_17_FFY_RST : STD_LOGIC; 
  signal mac_control_din_1_FFY_RST : STD_LOGIC; 
  signal mac_control_din_3_FFY_RST : STD_LOGIC; 
  signal mac_control_din_3_FFX_RST : STD_LOGIC; 
  signal mac_control_din_5_FFY_RST : STD_LOGIC; 
  signal mac_control_din_7_FFY_RST : STD_LOGIC; 
  signal mac_control_din_5_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_11_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_21_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_21_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_13_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_13_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_23_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_23_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_15_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_15_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_31_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_31_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_17_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_25_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_17_FFX_RST : STD_LOGIC; 
  signal mac_control_lrxmcast_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_11_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_11_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_21_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_21_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_13_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_13_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_31_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_31_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_23_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_23_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_15_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_25_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_27_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_29_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcll_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_24_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_16_FFY_RST : STD_LOGIC; 
  signal mac_control_din_7_FFX_RST : STD_LOGIC; 
  signal tx_output_outsell_0_FFY_SET : STD_LOGIC; 
  signal memcontroller_oel_FFY_RST : STD_LOGIC; 
  signal mac_control_din_9_FFY_RST : STD_LOGIC; 
  signal mac_control_din_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_macnt_72_FFY_RST : STD_LOGIC; 
  signal rx_output_cs_FFd18_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_11_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_21_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_11_FFX_RST : STD_LOGIC; 
  signal macaddr_31_FFX_RST : STD_LOGIC; 
  signal macaddr_23_FFX_RST : STD_LOGIC; 
  signal macaddr_15_FFX_RST : STD_LOGIC; 
  signal macaddr_33_FFX_RST : STD_LOGIC; 
  signal macaddr_41_FFX_RST : STD_LOGIC; 
  signal macaddr_25_FFX_RST : STD_LOGIC; 
  signal macaddr_17_FFX_RST : STD_LOGIC; 
  signal macaddr_27_FFX_RST : STD_LOGIC; 
  signal macaddr_43_FFY_RST : STD_LOGIC; 
  signal mac_control_din_21_FFX_RST : STD_LOGIC; 
  signal mac_control_din_15_FFY_RST : STD_LOGIC; 
  signal mac_control_din_15_FFX_RST : STD_LOGIC; 
  signal mac_control_din_23_FFY_RST : STD_LOGIC; 
  signal mac_control_din_23_FFX_RST : STD_LOGIC; 
  signal mac_control_din_31_FFY_RST : STD_LOGIC; 
  signal mac_control_din_31_FFX_RST : STD_LOGIC; 
  signal mac_control_din_17_FFY_RST : STD_LOGIC; 
  signal mac_control_din_17_FFX_RST : STD_LOGIC; 
  signal mac_control_din_25_FFY_RST : STD_LOGIC; 
  signal mac_control_din_25_FFX_RST : STD_LOGIC; 
  signal mac_control_din_19_FFY_RST : STD_LOGIC; 
  signal mac_control_din_19_FFX_RST : STD_LOGIC; 
  signal mac_control_din_27_FFY_RST : STD_LOGIC; 
  signal mac_control_din_27_FFX_RST : STD_LOGIC; 
  signal mac_control_din_29_FFY_RST : STD_LOGIC; 
  signal macaddr_35_FFX_RST : STD_LOGIC; 
  signal macaddr_43_FFX_RST : STD_LOGIC; 
  signal macaddr_19_FFX_RST : STD_LOGIC; 
  signal macaddr_29_FFX_RST : STD_LOGIC; 
  signal macaddr_37_FFX_RST : STD_LOGIC; 
  signal macaddr_45_FFX_RST : STD_LOGIC; 
  signal macaddr_39_FFX_RST : STD_LOGIC; 
  signal macaddr_47_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_addrl_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxmcastl_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_5_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_7_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_9_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_dinl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_21_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_13_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_13_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_23_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_31_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_31_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_23_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_15_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_15_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_25_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_25_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_17_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_17_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_27_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_27_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_19_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_19_FFX_RST : STD_LOGIC; 
  signal mac_control_phydi_29_FFY_RST : STD_LOGIC; 
  signal mac_control_phydi_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_1_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_3_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_5_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_5_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_7_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_9_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_MII_Interface_cs_FFd6_FFY_SET : STD_LOGIC; 
  signal rx_input_memio_addrchk_cs_FFd6_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_11_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_11_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_13_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_13_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_15_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_din_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_18_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_26_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_1_FFY_RST : STD_LOGIC; 
  signal memcontroller_clknum_1_FFX_RST : STD_LOGIC; 
  signal txfbbp_1_FFY_RST : STD_LOGIC; 
  signal txfbbp_3_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_3_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_3_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_5_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_5_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_7_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_7_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_rxbcastl_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_11_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_11_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_21_FFY_RST : STD_LOGIC; 
  signal txfbbp_1_FFX_RST : STD_LOGIC; 
  signal txfbbp_3_FFX_RST : STD_LOGIC; 
  signal txfbbp_5_FFY_RST : STD_LOGIC; 
  signal txfbbp_5_FFX_RST : STD_LOGIC; 
  signal txfbbp_7_FFY_RST : STD_LOGIC; 
  signal txfbbp_7_FFX_RST : STD_LOGIC; 
  signal txfbbp_9_FFY_RST : STD_LOGIC; 
  signal txfbbp_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_11_FFX_RST : STD_LOGIC; 
  signal mac_control_lrxbcast_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_21_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_21_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_13_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_7_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_8_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_5_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_1_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_1_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d1_9_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_control_d1_9_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_7_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_31_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_31_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_23_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_23_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_15_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_25_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_25_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_17_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_17_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_27_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_19_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_19_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_doutl_29_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_7_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_3_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_3_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_5_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_8_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_5_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d2_9_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_control_d2_9_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_7_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_7_FFX_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_9_FFY_SET : STD_LOGIC; 
  signal rx_input_fifo_control_d3_9_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_d3_8_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_27_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_28_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_crcl_29_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_celll_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_11_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_25_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_17_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_17_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_27_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_27_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_19_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_19_FFX_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_29_FFY_RST : STD_LOGIC; 
  signal mac_control_rxoferr_cntl_29_FFX_RST : STD_LOGIC; 
  signal rx_input_GMII_rx_dvll_FFY_RST : STD_LOGIC; 
  signal mac_control_lrxucast_FFY_RST : STD_LOGIC; 
  signal rx_input_fifo_control_cell_FFY_RST : STD_LOGIC; 
  signal addr4ext_11_FFY_RST : STD_LOGIC; 
  signal addr4ext_11_FFX_RST : STD_LOGIC; 
  signal addr4ext_13_FFY_RST : STD_LOGIC; 
  signal addr4ext_13_FFX_RST : STD_LOGIC; 
  signal addr4ext_15_FFY_RST : STD_LOGIC; 
  signal addr4ext_15_FFX_RST : STD_LOGIC; 
  signal d4_11_FFY_RST : STD_LOGIC; 
  signal d4_11_FFX_RST : STD_LOGIC; 
  signal d4_21_FFY_RST : STD_LOGIC; 
  signal d4_21_FFX_RST : STD_LOGIC; 
  signal d4_13_FFY_RST : STD_LOGIC; 
  signal d4_13_FFX_RST : STD_LOGIC; 
  signal d4_15_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_21_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_13_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_13_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_31_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_31_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_23_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_23_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_15_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_15_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_25_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_25_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_17_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_17_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_27_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_25_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_19_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_19_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_27_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_27_FFX_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_29_FFY_RST : STD_LOGIC; 
  signal mac_control_rxcrcerr_cntl_29_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd3_FFY_RST : STD_LOGIC; 
  signal mac_control_ledrx_rst_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_addrchk_validmcast_FFY_RST : STD_LOGIC; 
  signal mac_control_ledtx_rst_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd4_FFY_RST : STD_LOGIC; 
  signal d4_23_FFX_RST : STD_LOGIC; 
  signal d4_15_FFX_RST : STD_LOGIC; 
  signal d4_31_FFX_RST : STD_LOGIC; 
  signal d4_17_FFX_RST : STD_LOGIC; 
  signal d4_25_FFY_RST : STD_LOGIC; 
  signal d4_25_FFX_RST : STD_LOGIC; 
  signal d4_19_FFY_RST : STD_LOGIC; 
  signal d4_19_FFX_RST : STD_LOGIC; 
  signal d4_27_FFY_RST : STD_LOGIC; 
  signal d4_27_FFX_RST : STD_LOGIC; 
  signal mac_control_rxf_cntl_1_FFY_RST : STD_LOGIC; 
  signal d4_29_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_7_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_9_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_9_FFX_RST : STD_LOGIC; 
  signal mac_control_addr_1_FFY_RST : STD_LOGIC; 
  signal mac_control_addr_1_FFX_RST : STD_LOGIC; 
  signal mac_control_addr_3_FFY_RST : STD_LOGIC; 
  signal mac_control_addr_3_FFX_RST : STD_LOGIC; 
  signal mac_control_addr_5_FFY_RST : STD_LOGIC; 
  signal mac_control_addr_5_FFX_RST : STD_LOGIC; 
  signal mac_control_din_11_FFY_RST : STD_LOGIC; 
  signal mac_control_addr_7_FFY_RST : STD_LOGIC; 
  signal mac_control_addr_7_FFX_RST : STD_LOGIC; 
  signal mac_control_din_11_FFX_RST : STD_LOGIC; 
  signal mac_control_din_13_FFY_RST : STD_LOGIC; 
  signal mac_control_din_13_FFX_RST : STD_LOGIC; 
  signal mac_control_din_21_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_27_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_19_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_19_FFX_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_29_FFY_RST : STD_LOGIC; 
  signal mac_control_rxphyerr_cntl_29_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_11_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_11_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_13_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_13_FFX_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_15_FFY_RST : STD_LOGIC; 
  signal tx_fifocheck_bpl_15_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_19_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_27_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_37_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_37_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_45_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_45_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_29_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_29_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_39_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_39_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_47_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_47_FFX_RST : STD_LOGIC; 
  signal rxbp_11_FFY_RST : STD_LOGIC; 
  signal rxbp_11_FFX_RST : STD_LOGIC; 
  signal rxbp_13_FFY_RST : STD_LOGIC; 
  signal rxbp_15_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_31_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_15_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_15_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_41_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_33_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_33_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_41_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_17_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_17_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_25_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_25_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_35_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_35_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_43_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_43_FFX_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_19_FFY_RST : STD_LOGIC; 
  signal mac_control_lmacaddr_27_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_11_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_11_FFX_RST : STD_LOGIC; 
  signal tx_input_dh_13_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_13_FFX_RST : STD_LOGIC; 
  signal tx_input_dh_15_FFY_RST : STD_LOGIC; 
  signal tx_input_dh_15_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_11_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_11_FFX_RST : STD_LOGIC; 
  signal txbp_11_FFY_RST : STD_LOGIC; 
  signal txbp_11_FFX_RST : STD_LOGIC; 
  signal tx_input_dl_13_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_13_FFX_RST : STD_LOGIC; 
  signal txbp_13_FFY_RST : STD_LOGIC; 
  signal tx_input_dl_15_FFY_RST : STD_LOGIC; 
  signal txbp_13_FFX_RST : STD_LOGIC; 
  signal tx_output_outsell_2_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_fifofulll_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_endbyte_1_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_endbyte_2_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_endbyte_1_FFX_RST : STD_LOGIC; 
  signal rx_output_nfl_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_1_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_1_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_3_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_3_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_5_FFY_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_5_FFX_RST : STD_LOGIC; 
  signal mac_control_txf_cntl_7_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_9_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_11_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_11_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_13_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_13_FFX_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_15_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_bpl_15_FFX_RST : STD_LOGIC; 
  signal rxf_FFY_RST : STD_LOGIC; 
  signal tx_output_crcl_4_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_1_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_1_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_3_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_5_FFY_RST : STD_LOGIC; 
  signal rxbp_13_FFX_RST : STD_LOGIC; 
  signal rxbp_15_FFX_RST : STD_LOGIC; 
  signal q2_1_FFY_RST : STD_LOGIC; 
  signal q2_1_FFX_RST : STD_LOGIC; 
  signal q2_2_FFY_RST : STD_LOGIC; 
  signal q2_3_FFY_RST : STD_LOGIC; 
  signal q2_5_FFY_RST : STD_LOGIC; 
  signal q2_5_FFX_RST : STD_LOGIC; 
  signal q3_1_FFY_RST : STD_LOGIC; 
  signal q3_1_FFX_RST : STD_LOGIC; 
  signal q2_7_FFY_RST : STD_LOGIC; 
  signal q2_7_FFX_RST : STD_LOGIC; 
  signal q3_2_FFY_RST : STD_LOGIC; 
  signal q3_3_FFY_RST : STD_LOGIC; 
  signal q2_9_FFY_RST : STD_LOGIC; 
  signal q2_9_FFX_RST : STD_LOGIC; 
  signal q3_5_FFY_RST : STD_LOGIC; 
  signal q3_5_FFX_RST : STD_LOGIC; 
  signal q3_7_FFY_RST : STD_LOGIC; 
  signal q3_7_FFX_RST : STD_LOGIC; 
  signal q3_9_FFY_RST : STD_LOGIC; 
  signal q3_9_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_11_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_11_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_13_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_13_FFX_RST : STD_LOGIC; 
  signal tx_output_bpl_15_FFY_RST : STD_LOGIC; 
  signal tx_output_bpl_15_FFX_RST : STD_LOGIC; 
  signal tx_output_outsell_2_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_3_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_5_FFX_RST : STD_LOGIC; 
  signal mac_control_phyaddr_7_FFY_RST : STD_LOGIC; 
  signal mac_control_phyaddr_7_FFX_RST : STD_LOGIC; 
  signal mac_control_din_29_FFX_RST : STD_LOGIC; 
  signal memcontroller_ts_0_FFY_SET : STD_LOGIC; 
  signal tx_output_crcl_3_FFY_RST : STD_LOGIC; 
  signal rx_input_memio_cs_FFd16_2_FFY_SET : STD_LOGIC; 
  signal mac_control_PHY_status_dout_1_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_1_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_3_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_3_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_5_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_5_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_7_FFY_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_7_FFX_RST : STD_LOGIC; 
  signal mac_control_PHY_status_dout_9_FFY_RST : STD_LOGIC; 
  signal clkio_bufg_CE : STD_LOGIC; 
  signal clk_bufg_CE : STD_LOGIC; 
  signal clkrx_bufg_CE : STD_LOGIC; 
  signal PWR_GND_0_GROM : STD_LOGIC; 
  signal PWR_GND_1_GROM : STD_LOGIC; 
  signal PWR_GND_2_GROM : STD_LOGIC; 
  signal PWR_GND_3_GROM : STD_LOGIC; 
  signal PWR_GND_4_GROM : STD_LOGIC; 
  signal PWR_GND_5_GROM : STD_LOGIC; 
  signal PWR_GND_6_GROM : STD_LOGIC; 
  signal PWR_GND_7_GROM : STD_LOGIC; 
  signal PWR_GND_8_GROM : STD_LOGIC; 
  signal PWR_GND_9_FROM : STD_LOGIC; 
  signal PWR_GND_9_GROM : STD_LOGIC; 
  signal PWR_GND_10_FROM : STD_LOGIC; 
  signal PWR_GND_10_GROM : STD_LOGIC; 
  signal PWR_GND_11_FROM : STD_LOGIC; 
  signal PWR_GND_11_GROM : STD_LOGIC; 
  signal PWR_GND_12_FROM : STD_LOGIC; 
  signal PWR_GND_12_GROM : STD_LOGIC; 
  signal PWR_GND_13_FROM : STD_LOGIC; 
  signal PWR_GND_13_GROM : STD_LOGIC; 
  signal PWR_GND_14_FROM : STD_LOGIC; 
  signal PWR_GND_14_GROM : STD_LOGIC; 
  signal PWR_GND_15_GROM : STD_LOGIC; 
  signal PWR_GND_16_GROM : STD_LOGIC; 
  signal PWR_GND_17_FROM : STD_LOGIC; 
  signal PWR_GND_17_GROM : STD_LOGIC; 
  signal PWR_GND_18_GROM : STD_LOGIC; 
  signal PWR_GND_19_FROM : STD_LOGIC; 
  signal PWR_GND_19_GROM : STD_LOGIC; 
  signal PWR_GND_20_GROM : STD_LOGIC; 
  signal PWR_GND_21_GROM : STD_LOGIC; 
  signal PWR_GND_22_GROM : STD_LOGIC; 
  signal PWR_GND_23_FROM : STD_LOGIC; 
  signal PWR_GND_23_GROM : STD_LOGIC; 
  signal PWR_GND_24_GROM : STD_LOGIC; 
  signal PWR_GND_25_FROM : STD_LOGIC; 
  signal PWR_GND_25_GROM : STD_LOGIC; 
  signal PWR_GND_26_GROM : STD_LOGIC; 
  signal PWR_GND_27_GROM : STD_LOGIC; 
  signal PWR_GND_28_GROM : STD_LOGIC; 
  signal PWR_GND_29_FROM : STD_LOGIC; 
  signal PWR_GND_29_GROM : STD_LOGIC; 
  signal PWR_GND_30_FROM : STD_LOGIC; 
  signal PWR_GND_30_GROM : STD_LOGIC; 
  signal PWR_GND_31_GROM : STD_LOGIC; 
  signal PWR_GND_32_GROM : STD_LOGIC; 
  signal PWR_GND_33_GROM : STD_LOGIC; 
  signal PWR_GND_34_GROM : STD_LOGIC; 
  signal PWR_GND_35_FROM : STD_LOGIC; 
  signal PWR_GND_35_GROM : STD_LOGIC; 
  signal PWR_GND_36_FROM : STD_LOGIC; 
  signal PWR_GND_36_GROM : STD_LOGIC; 
  signal PWR_GND_37_FROM : STD_LOGIC; 
  signal PWR_GND_37_GROM : STD_LOGIC; 
  signal PWR_GND_38_FROM : STD_LOGIC; 
  signal PWR_GND_38_GROM : STD_LOGIC; 
  signal PWR_GND_39_GROM : STD_LOGIC; 
  signal PWR_GND_40_FROM : STD_LOGIC; 
  signal PWR_GND_40_GROM : STD_LOGIC; 
  signal PWR_GND_41_GROM : STD_LOGIC; 
  signal PWR_GND_42_FROM : STD_LOGIC; 
  signal PWR_GND_42_GROM : STD_LOGIC; 
  signal PWR_GND_43_GROM : STD_LOGIC; 
  signal PWR_GND_44_FROM : STD_LOGIC; 
  signal PWR_GND_44_GROM : STD_LOGIC; 
  signal PWR_GND_45_FROM : STD_LOGIC; 
  signal PWR_GND_45_GROM : STD_LOGIC; 
  signal PWR_GND_46_FROM : STD_LOGIC; 
  signal PWR_GND_46_GROM : STD_LOGIC; 
  signal PWR_GND_47_GROM : STD_LOGIC; 
  signal PWR_GND_48_GROM : STD_LOGIC; 
  signal PWR_GND_49_GROM : STD_LOGIC; 
  signal PWR_GND_50_FROM : STD_LOGIC; 
  signal PWR_GND_50_GROM : STD_LOGIC; 
  signal PWR_VCC_0_FROM : STD_LOGIC; 
  signal PWR_VCC_1_FROM : STD_LOGIC; 
  signal PWR_VCC_2_FROM : STD_LOGIC; 
  signal PWR_VCC_3_FROM : STD_LOGIC; 
  signal PWR_VCC_4_FROM : STD_LOGIC; 
  signal PWR_VCC_5_FROM : STD_LOGIC; 
  signal PWR_VCC_6_FROM : STD_LOGIC; 
  signal PWR_VCC_7_FROM : STD_LOGIC; 
  signal PWR_VCC_8_FROM : STD_LOGIC; 
  signal PWR_VCC_9_FROM : STD_LOGIC; 
  signal PWR_VCC_10_FROM : STD_LOGIC; 
  signal PWR_VCC_11_FROM : STD_LOGIC; 
  signal PWR_VCC_12_FROM : STD_LOGIC; 
  signal VCC : STD_LOGIC; 
  signal GND : STD_LOGIC; 
  signal rx_input_fifo_dout : STD_LOGIC_VECTOR ( 9 downto 9 ); 
  signal mac_control_din : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_phyaddr : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_crcll : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_PHY_status_MII_Interface_statecnt : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal rx_input_data : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal rx_input_memio_dout : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal addr2ext : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal txfbbp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_PHY_status_din : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_fifo_control_d1 : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal rx_input_fifo_control_d0 : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal rx_input_fifo_control_d3 : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal rx_input_fifo_control_d2 : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal q2 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_fifo_control_ldata : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_18_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_crc_loigc_n0115 : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_crc_loigc_n0124 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_n0007_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_crcl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_addr : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal mac_control_lmacaddr : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal macaddr : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal tx_output_data : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal tx_output_crc_loigc_n0122 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_7_Xo : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal tx_output_crc_loigc_n0118 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal tx_input_CNT : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_phydo : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_dout : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_phydi : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_rxfifowerr_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_rxfifowerr_cntl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_crcl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_datal : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal rx_input_memio_crccomb_Mxor_CO_18_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_input_memio_crccomb_n0104 : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_input_memio_crccomb_Mxor_CO_23_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_input_memio_crccomb_n0122 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal tx_output_crc_loigc_n0104 : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_9_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_output_fifo_wrcount : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal addr4ext : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_input_dl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal d4 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal tx_fifocheck_fbbpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_rxphyerr_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_rxphyerr_cntl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_PHY_status_MII_Interface_dreg : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_input_dinint : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_input_dh : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_crccomb_n0118 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal rx_input_memio_crccomb_n0124 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal txbp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rxbp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_addrchk_macaddrl : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal memcontroller_clknum : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal mac_control_rxcrcerr_cntl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_rxf_cntl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_rxoferr_cntl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_txfifowerr_cntl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_txf_cntl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_phystat : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_crccomb_Mxor_CO_7_Xo : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal rx_input_memio_crccomb_Mxor_CO_9_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_crcsell : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rx_input_memio_addrchk_datal : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal rx_input_memio_addrchk_mcast : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_ncrcbytel : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal mac_control_PHY_status_dout : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_crccomb_Mxor_n0007_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal mac_control_rxf_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_fifocheck_diff : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_rxoferr_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_txfifowerr_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_addrchk_bcast : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal tx_output_bcntl : STD_LOGIC_VECTOR ( 15 downto 1 ); 
  signal rx_output_bp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rxfbbp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal memcontroller_qn : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal q3 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_output_mdl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_output_len : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_output_datal : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_23_Xo : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_outselll : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal tx_output_ltxd : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal rx_input_memio_crccomb_n0115 : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_outsell : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal mac_control_txf_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_output_fifodout : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_GMII_rxdl : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal tx_input_dinl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal memcontroller_addrn : STD_LOGIC_VECTOR ( 16 downto 0 ); 
  signal memcontroller_dnl2 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_ts : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal rx_input_fifoin : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal rx_input_fifo_fifodout : STD_LOGIC_VECTOR ( 8 downto 0 ); 
  signal rx_output_fifodin : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal addr3ext : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal addr1ext : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal d1 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_dnl1 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal mac_control_PHY_status_MII_Interface_n0076 : STD_LOGIC_VECTOR ( 5 downto 1 ); 
  signal rx_output_n0060 : STD_LOGIC_VECTOR ( 15 downto 2 ); 
  signal rx_input_memio_addrchk_lmaceq : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal mac_control_rxcrcerr_cnt : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_bp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_output_lenr : STD_LOGIC_VECTOR ( 15 downto 2 ); 
  signal rx_fifocheck_fbbpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_fifocheck_bpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_fifocheck_bpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_fifocheck_diff : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_input_n0074 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_output_n0070 : STD_LOGIC_VECTOR ( 15 downto 2 ); 
  signal tx_output_bpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_bcntl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_13_Xo : STD_LOGIC_VECTOR ( 2 downto 2 ); 
  signal rx_input_memio_crccomb_Mxor_CO_13_Xo : STD_LOGIC_VECTOR ( 2 downto 2 ); 
  signal rx_input_memio_bpl : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_doutl : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_endbyte : STD_LOGIC_VECTOR ( 2 downto 0 ); 
  signal rx_input_memio_addrchk_maceq : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal mac_control_PHY_status_addrl : STD_LOGIC_VECTOR ( 4 downto 0 ); 
  signal mac_control_PHY_status_miiaddr : STD_LOGIC_VECTOR ( 4 downto 0 ); 
  signal tx_output_crc_loigc_Mxor_CO_26_Xo : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal rx_input_memio_crccomb_Mxor_CO_26_Xo : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal rx_input_fifo_control_dinl : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal mac_control_n0016 : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_input_memio_addrchk_lmcast : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_ncrcbyte : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal tx_output_crcsel : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal tx_output_ldata : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal rx_input_memio_addrchk_lbcast : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal memcontroller_addr : STD_LOGIC_VECTOR ( 16 downto 0 ); 
  signal memcontroller_dnout : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_q : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal memcontroller_dn : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal tx_output_addr_n0000 : STD_LOGIC_VECTOR ( 15 downto 1 ); 
  signal mac_control_rxcrcerr_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal rx_input_memio_n0043 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_rxoferr_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal mac_control_rxphyerr_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal mac_control_rxfifowerr_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal mac_control_txfifowerr_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal rx_output_lbp : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_fifocheck_n0001 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_fifocheck_n0001 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_txf_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal rx_input_memio_n0042 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal mac_control_rxf_cnt_n0000 : STD_LOGIC_VECTOR ( 31 downto 1 ); 
  signal mac_control_PHY_status_MII_Interface_n0014 : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal rx_input_memio_lma : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal rx_input_memio_lmd : STD_LOGIC_VECTOR ( 31 downto 0 ); 
  signal rx_output_lma : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_input_n0032 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal tx_input_ldinint : STD_LOGIC_VECTOR ( 15 downto 0 ); 
begin
  rx_input_fifo_fifo_N1559_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1559_FFY_SET
    );
  rx_input_fifo_fifo_BU412 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N1552,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1559_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1559
    );
  rx_input_fifo_fifo_N1552_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1552_FFY_SET
    );
  rx_input_fifo_fifo_BU354 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N1524,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1552_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1552
    );
  rx_input_fifo_fifo_N1573_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1573_FFY_SET
    );
  rx_input_fifo_fifo_BU338 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1573_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1573
    );
  rx_input_fifo_fifo_N1538_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1538_FFY_SET
    );
  rx_input_fifo_fifo_BU289 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N1524,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N1538_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1538
    );
  rx_input_fifo_fifo_BU169 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_full,
      ADR1 => rx_input_ince,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N1497_FROM
    );
  rx_input_fifo_fifo_BU175 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_full,
      ADR1 => rx_input_ince,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N1497_GROM
    );
  rx_input_fifo_fifo_N1497_XUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1497_FROM,
      O => rx_input_fifo_fifo_N1497
    );
  rx_input_fifo_fifo_N1497_YUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1497_GROM,
      O => rx_input_fifo_fifo_N17
    );
  rx_input_fifo_fifo_full_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_full_FFY_SET
    );
  rx_input_fifo_fifo_BU321 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3374,
      CE => rx_input_fifo_fifo_N3373,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_full_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_full
    );
  rx_input_fifo_fifo_full_LOGIC_ZERO_4 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_full_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU317 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_full_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_full_CYINIT,
      SEL => rx_input_fifo_fifo_N3358,
      O => rx_input_fifo_fifo_BU317_O
    );
  rx_input_fifo_fifo_BU316 : X_LUT4
    generic map(
      INIT => X"E14B"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_full,
      ADR1 => rx_input_fifo_fifo_N1545,
      ADR2 => rx_input_fifo_fifo_N1580,
      ADR3 => rx_input_fifo_fifo_N1538,
      O => rx_input_fifo_fifo_N3358
    );
  rx_input_fifo_fifo_full_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_full_GROM
    );
  rx_input_fifo_fifo_BU320 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_BU317_O,
      I1 => rx_input_fifo_fifo_full_GROM,
      O => rx_input_fifo_fifo_N3374
    );
  rx_input_fifo_fifo_full_CYINIT_5 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3366,
      O => rx_input_fifo_fifo_full_CYINIT
    );
  rx_input_fifo_fifo_N1580_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1580_FFY_SET
    );
  rx_input_fifo_fifo_BU272 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3239,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1580_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1580
    );
  rx_input_fifo_fifo_BU271 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N2,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3239
    );
  rx_input_fifo_fifo_N2_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N2_FFX_RST
    );
  rx_input_fifo_fifo_BU221 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2690,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N2_FFX_RST,
      O => rx_input_fifo_fifo_N2
    );
  rx_input_fifo_fifo_BU219 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N2_CYINIT,
      I1 => rx_input_fifo_fifo_N2721,
      O => rx_input_fifo_fifo_N2690
    );
  rx_input_fifo_fifo_BU218 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N2,
      O => rx_input_fifo_fifo_N2721
    );
  rx_input_fifo_fifo_N2_CYINIT_6 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2718,
      O => rx_input_fifo_fifo_N2_CYINIT
    );
  rx_input_fifo_fifo_N1545_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1545_FFX_SET
    );
  rx_input_fifo_fifo_BU315 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N1538,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N1545_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1545
    );
  rx_input_fifo_fifo_N1545_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1545_FFY_RST
    );
  rx_input_fifo_fifo_BU312 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1539,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1545_FFY_RST,
      O => rx_input_fifo_fifo_N1546
    );
  rx_input_fifo_fifo_N1545_LOGIC_ZERO_7 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N1545_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU311 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1545_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N1545_CYINIT,
      SEL => rx_input_fifo_fifo_N3360,
      O => rx_input_fifo_fifo_N3367
    );
  rx_input_fifo_fifo_BU310 : X_LUT4
    generic map(
      INIT => X"A5C3"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1540,
      ADR1 => rx_input_fifo_fifo_N1547,
      ADR2 => rx_input_fifo_fifo_N1582,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N3360
    );
  rx_input_fifo_fifo_BU313 : X_LUT4
    generic map(
      INIT => X"C963"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_full,
      ADR1 => rx_input_fifo_fifo_N1581,
      ADR2 => rx_input_fifo_fifo_N1546,
      ADR3 => rx_input_fifo_fifo_N1539,
      O => rx_input_fifo_fifo_N3359
    );
  rx_input_fifo_fifo_N1545_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1545_CYMUXG,
      O => rx_input_fifo_fifo_N3366
    );
  rx_input_fifo_fifo_BU314 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1545_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N3367,
      SEL => rx_input_fifo_fifo_N3359,
      O => rx_input_fifo_fifo_N1545_CYMUXG
    );
  rx_input_fifo_fifo_N1545_CYINIT_8 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3368,
      O => rx_input_fifo_fifo_N1545_CYINIT
    );
  rx_input_rx_nearf_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_rx_nearf_FFX_RST
    );
  rx_input_fifo_fifo_BU443 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N4297,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_rx_nearf_FFX_RST,
      O => rx_input_rx_nearf
    );
  rx_input_fifo_fifo_BU441 : X_XOR2
    port map (
      I0 => rx_input_rx_nearf_CYINIT,
      I1 => rx_input_fifo_fifo_N4324,
      O => rx_input_fifo_fifo_N4297
    );
  rx_input_fifo_fifo_BU439 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1573,
      ADR1 => rx_input_fifo_fifo_N1559,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4324
    );
  rx_input_rx_nearf_CYINIT_9 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4321,
      O => rx_input_rx_nearf_CYINIT
    );
  rx_input_fifo_fifo_N1582_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1582_FFY_RST
    );
  rx_input_fifo_fifo_BU265 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3199,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1582_FFY_RST,
      O => rx_input_fifo_fifo_N1581
    );
  rx_input_fifo_fifo_BU257 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N4,
      O => rx_input_fifo_fifo_N3159
    );
  rx_input_fifo_fifo_BU264 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N2,
      ADR1 => rx_input_fifo_fifo_N3,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3199
    );
  rx_input_fifo_fifo_BU207 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N4,
      IB => rx_input_fifo_fifo_N4_CYINIT,
      SEL => rx_input_fifo_fifo_N2711,
      O => rx_input_fifo_fifo_N2713
    );
  rx_input_fifo_fifo_BU208 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N4_CYINIT,
      I1 => rx_input_fifo_fifo_N2711,
      O => rx_input_fifo_fifo_N2688
    );
  rx_input_fifo_fifo_BU206 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N4,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2711
    );
  rx_input_fifo_fifo_BU212 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2716
    );
  rx_input_fifo_fifo_N4_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4_CYMUXG,
      O => rx_input_fifo_fifo_N2718
    );
  rx_input_fifo_fifo_BU213 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N3,
      IB => rx_input_fifo_fifo_N2713,
      SEL => rx_input_fifo_fifo_N2716,
      O => rx_input_fifo_fifo_N4_CYMUXG
    );
  rx_input_fifo_fifo_BU214 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N2713,
      I1 => rx_input_fifo_fifo_N2716,
      O => rx_input_fifo_fifo_N2689
    );
  rx_input_fifo_fifo_N4_CYINIT_10 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2708,
      O => rx_input_fifo_fifo_N4_CYINIT
    );
  rx_input_fifo_fifo_N1547_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1547_FFY_RST
    );
  rx_input_fifo_fifo_BU306 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1541,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1547_FFY_RST,
      O => rx_input_fifo_fifo_N1548
    );
  rx_input_fifo_fifo_N1547_LOGIC_ZERO_11 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N1547_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU305 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1547_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N1547_CYINIT,
      SEL => rx_input_fifo_fifo_N3362,
      O => rx_input_fifo_fifo_N3369
    );
  rx_input_fifo_fifo_BU304 : X_LUT4
    generic map(
      INIT => X"E12D"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1549,
      ADR1 => rx_input_fifo_fifo_full,
      ADR2 => rx_input_fifo_fifo_N1584,
      ADR3 => rx_input_fifo_fifo_N1542,
      O => rx_input_fifo_fifo_N3362
    );
  rx_input_fifo_fifo_BU307 : X_LUT4
    generic map(
      INIT => X"C963"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_full,
      ADR1 => rx_input_fifo_fifo_N1583,
      ADR2 => rx_input_fifo_fifo_N1548,
      ADR3 => rx_input_fifo_fifo_N1541,
      O => rx_input_fifo_fifo_N3361
    );
  rx_input_fifo_fifo_N1547_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1547_CYMUXG,
      O => rx_input_fifo_fifo_N3368
    );
  rx_input_fifo_fifo_BU308 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1547_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N3369,
      SEL => rx_input_fifo_fifo_N3361,
      O => rx_input_fifo_fifo_N1547_CYMUXG
    );
  rx_input_fifo_fifo_N1547_CYINIT_12 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N3370,
      O => rx_input_fifo_fifo_N1547_CYINIT
    );
  rx_input_fifo_fifo_N1574_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1574_FFY_SET
    );
  rx_input_fifo_fifo_BU334 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N4,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1574_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1575
    );
  rx_input_fifo_fifo_BU431 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1575,
      IB => rx_input_fifo_fifo_N4321_CYINIT,
      SEL => rx_input_fifo_fifo_N4314,
      O => rx_input_fifo_fifo_N4317
    );
  rx_input_fifo_fifo_BU430 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1575,
      ADR1 => rx_input_fifo_fifo_N1561,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4314
    );
  rx_input_fifo_fifo_BU433 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1574,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N1560,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4318
    );
  rx_input_fifo_fifo_N4321_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4321_CYMUXG,
      O => rx_input_fifo_fifo_N4321
    );
  rx_input_fifo_fifo_BU434 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1574,
      IB => rx_input_fifo_fifo_N4317,
      SEL => rx_input_fifo_fifo_N4318,
      O => rx_input_fifo_fifo_N4321_CYMUXG
    );
  rx_input_fifo_fifo_N4321_CYINIT_13 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4313,
      O => rx_input_fifo_fifo_N4321_CYINIT
    );
  rx_input_fifo_fifo_BU366 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1552,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N1553,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3689
    );
  rx_input_fifo_fifo_BU372 : X_LUT4
    generic map(
      INIT => X"C33C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N1554,
      ADR2 => rx_input_fifo_fifo_N1553,
      ADR3 => rx_input_fifo_fifo_N1552,
      O => rx_input_fifo_fifo_N3688
    );
  rx_input_fifo_fifo_BU243 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N5,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N6,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N3079
    );
  rx_input_fifo_fifo_BU250 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N5,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N4,
      O => rx_input_fifo_fifo_N3119
    );
  rx_input_fifo_fifo_BU195 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N6,
      IB => rx_input_fifo_fifo_N6_CYINIT,
      SEL => rx_input_fifo_fifo_N2701,
      O => rx_input_fifo_fifo_N2703
    );
  rx_input_fifo_fifo_BU196 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N6_CYINIT,
      I1 => rx_input_fifo_fifo_N2701,
      O => rx_input_fifo_fifo_N2686
    );
  rx_input_fifo_fifo_BU194 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N6,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2701
    );
  rx_input_fifo_fifo_BU200 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N5,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2706
    );
  rx_input_fifo_fifo_N6_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N6_CYMUXG,
      O => rx_input_fifo_fifo_N2708
    );
  rx_input_fifo_fifo_BU201 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N5,
      IB => rx_input_fifo_fifo_N2703,
      SEL => rx_input_fifo_fifo_N2706,
      O => rx_input_fifo_fifo_N6_CYMUXG
    );
  rx_input_fifo_fifo_BU202 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N2703,
      I1 => rx_input_fifo_fifo_N2706,
      O => rx_input_fifo_fifo_N2687
    );
  rx_input_fifo_fifo_N6_CYINIT_14 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2698,
      O => rx_input_fifo_fifo_N6_CYINIT
    );
  rx_input_fifo_fifo_BU258 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3159,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1582_FFX_RST,
      O => rx_input_fifo_fifo_N1582
    );
  rx_input_fifo_fifo_N1582_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1582_FFX_RST
    );
  rx_input_fifo_fifo_N1549_LOGIC_ONE_15 : X_ONE
    port map (
      O => rx_input_fifo_fifo_N1549_LOGIC_ONE
    );
  rx_input_fifo_fifo_N1549_LOGIC_ZERO_16 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N1549_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU299 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1549_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N1549_LOGIC_ONE,
      SEL => rx_input_fifo_fifo_N3364,
      O => rx_input_fifo_fifo_N3371
    );
  rx_input_fifo_fifo_BU298 : X_LUT4
    generic map(
      INIT => X"C3A5"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1551,
      ADR1 => rx_input_fifo_fifo_N1544,
      ADR2 => rx_input_fifo_fifo_N1586,
      ADR3 => rx_input_fifo_fifo_full,
      O => rx_input_fifo_fifo_N3364
    );
  rx_input_fifo_fifo_BU301 : X_LUT4
    generic map(
      INIT => X"D287"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_full,
      ADR1 => rx_input_fifo_fifo_N1543,
      ADR2 => rx_input_fifo_fifo_N1585,
      ADR3 => rx_input_fifo_fifo_N1550,
      O => rx_input_fifo_fifo_N3363
    );
  rx_input_fifo_fifo_N1549_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1549_CYMUXG,
      O => rx_input_fifo_fifo_N3370
    );
  rx_input_fifo_fifo_BU302 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1549_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N3371,
      SEL => rx_input_fifo_fifo_N3363,
      O => rx_input_fifo_fifo_N1549_CYMUXG
    );
  rx_input_fifo_fifo_N1555_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1555_FFY_RST
    );
  rx_input_fifo_fifo_BU346 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1528,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1555_FFY_RST,
      O => rx_input_fifo_fifo_N1556
    );
  rx_input_fifo_fifo_N1576_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1576_FFY_SET
    );
  rx_input_fifo_fifo_BU330 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N6,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1576_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1577
    );
  rx_input_fifo_fifo_BU425 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1577,
      IB => rx_input_fifo_fifo_N4313_CYINIT,
      SEL => rx_input_fifo_fifo_N4306,
      O => rx_input_fifo_fifo_N4309
    );
  rx_input_fifo_fifo_BU424 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1577,
      ADR1 => rx_input_fifo_fifo_N1563,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4306
    );
  rx_input_fifo_fifo_BU427 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1576,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N1562,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4310
    );
  rx_input_fifo_fifo_N4313_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4313_CYMUXG,
      O => rx_input_fifo_fifo_N4313
    );
  rx_input_fifo_fifo_BU428 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1576,
      IB => rx_input_fifo_fifo_N4309,
      SEL => rx_input_fifo_fifo_N4310,
      O => rx_input_fifo_fifo_N4313_CYMUXG
    );
  rx_input_fifo_fifo_N4313_CYINIT_17 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4305,
      O => rx_input_fifo_fifo_N4313_CYINIT
    );
  rx_input_fifo_fifo_BU216 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2689,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N4_FFY_RST,
      O => rx_input_fifo_fifo_N3
    );
  rx_input_fifo_fifo_N4_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N4_FFY_RST
    );
  rx_input_fifo_fifo_BU378 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1553,
      ADR1 => rx_input_fifo_fifo_N1552,
      ADR2 => rx_input_fifo_fifo_N1554,
      ADR3 => rx_input_fifo_fifo_N1555,
      O => rx_input_fifo_fifo_N1562_FROM
    );
  rx_input_fifo_fifo_BU384 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N1556,
      ADR3 => rx_input_fifo_fifo_N3676,
      O => rx_input_fifo_fifo_N3686
    );
  rx_input_fifo_fifo_N1562_XUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1562_FROM,
      O => rx_input_fifo_fifo_N3676
    );
  rx_input_fifo_fifo_BU285 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1526,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1539_FFY_RST,
      O => rx_input_fifo_fifo_N1540
    );
  rx_input_fifo_fifo_N1539_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1539_FFY_RST
    );
  rx_input_fifo_fifo_BU229 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N7,
      ADR2 => rx_input_fifo_fifo_N8,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2999
    );
  rx_input_fifo_fifo_BU236 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N7,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N6,
      O => rx_input_fifo_fifo_N3039
    );
  rx_input_fifo_fifo_N8_LOGIC_ZERO_18 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N8_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU183 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N8,
      IB => rx_input_fifo_fifo_N8_CYINIT,
      SEL => rx_input_fifo_fifo_N2691,
      O => rx_input_fifo_fifo_N2693
    );
  rx_input_fifo_fifo_BU184 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N8_CYINIT,
      I1 => rx_input_fifo_fifo_N2691,
      O => rx_input_fifo_fifo_N2684
    );
  rx_input_fifo_fifo_BU182 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N8,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2691
    );
  rx_input_fifo_fifo_BU188 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N7,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2696
    );
  rx_input_fifo_fifo_N8_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N8_CYMUXG,
      O => rx_input_fifo_fifo_N2698
    );
  rx_input_fifo_fifo_BU189 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N7,
      IB => rx_input_fifo_fifo_N2693,
      SEL => rx_input_fifo_fifo_N2696,
      O => rx_input_fifo_fifo_N8_CYMUXG
    );
  rx_input_fifo_fifo_BU190 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N2693,
      I1 => rx_input_fifo_fifo_N2696,
      O => rx_input_fifo_fifo_N2685
    );
  rx_input_fifo_fifo_N8_CYINIT_19 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N8_LOGIC_ZERO,
      O => rx_input_fifo_fifo_N8_CYINIT
    );
  rx_input_fifo_fifo_BU292 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_full,
      ADR3 => rx_input_ince,
      O => rx_input_fifo_fifo_N1550_GROM
    );
  rx_input_fifo_fifo_N1550_YUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1550_GROM,
      O => rx_input_fifo_fifo_N3373
    );
  rx_input_fifo_fifo_N1578_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1578_FFY_SET
    );
  rx_input_fifo_fifo_BU326 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N8,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1578_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1579
    );
  rx_input_fifo_fifo_N4305_LOGIC_ONE_20 : X_ONE
    port map (
      O => rx_input_fifo_fifo_N4305_LOGIC_ONE
    );
  rx_input_fifo_fifo_BU419 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1579,
      IB => rx_input_fifo_fifo_N4305_LOGIC_ONE,
      SEL => rx_input_fifo_fifo_N4298,
      O => rx_input_fifo_fifo_N4301
    );
  rx_input_fifo_fifo_BU418 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1579,
      ADR1 => rx_input_fifo_fifo_N1565,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4298
    );
  rx_input_fifo_fifo_BU421 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1578,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N1564,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N4302
    );
  rx_input_fifo_fifo_N4305_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N4305_CYMUXG,
      O => rx_input_fifo_fifo_N4305
    );
  rx_input_fifo_fifo_BU422 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1578,
      IB => rx_input_fifo_fifo_N4301,
      SEL => rx_input_fifo_fifo_N4302,
      O => rx_input_fifo_fifo_N4305_CYMUXG
    );
  rx_input_fifo_fifo_BU396 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1556,
      ADR1 => rx_input_fifo_fifo_N1558,
      ADR2 => rx_input_fifo_fifo_N1557,
      ADR3 => rx_input_fifo_fifo_N3676,
      O => rx_input_fifo_fifo_N3684
    );
  rx_input_fifo_fifo_BU390 : X_LUT4
    generic map(
      INIT => X"C33C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N3676,
      ADR2 => rx_input_fifo_fifo_N1557,
      ADR3 => rx_input_fifo_fifo_N1556,
      O => rx_input_fifo_fifo_N3685
    );
  rx_input_fifo_fifo_BU16 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_rd_en,
      ADR3 => rx_input_fifo_fifo_empty,
      O => rx_input_fifo_fifo_N1495_FROM
    );
  rx_input_fifo_fifo_BU22 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_rd_en,
      ADR3 => rx_input_fifo_fifo_empty,
      O => rx_input_fifo_fifo_N1495_GROM
    );
  rx_input_fifo_fifo_N1495_XUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1495_FROM,
      O => rx_input_fifo_fifo_N1495
    );
  rx_input_fifo_fifo_N1495_YUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1495_GROM,
      O => rx_input_fifo_fifo_N16
    );
  rx_input_fifo_fifo_BU29 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_empty,
      ADR1 => rx_input_fifo_rd_en,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N1794
    );
  rx_input_fifo_fifo_empty_LOGIC_ZERO_21 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_empty_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU156 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_empty_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_empty_CYINIT,
      SEL => rx_input_fifo_fifo_N2434,
      O => rx_input_fifo_fifo_BU156_O
    );
  rx_input_fifo_fifo_BU155 : X_LUT4
    generic map(
      INIT => X"A5C3"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1580,
      ADR1 => rx_input_fifo_fifo_N1594,
      ADR2 => rx_input_fifo_fifo_N1524,
      ADR3 => rx_input_fifo_fifo_empty,
      O => rx_input_fifo_fifo_N2434
    );
  rx_input_fifo_fifo_empty_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_empty_GROM
    );
  rx_input_fifo_fifo_BU159 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_BU156_O,
      I1 => rx_input_fifo_fifo_empty_GROM,
      O => rx_input_fifo_fifo_N2450
    );
  rx_input_fifo_fifo_empty_CYINIT_22 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2442,
      O => rx_input_fifo_fifo_empty_CYINIT
    );
  rx_input_fifo_fifo_BU126 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N9,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2412
    );
  rx_input_fifo_fifo_BU74 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N9_CYINIT,
      I1 => rx_input_fifo_fifo_N1894,
      O => rx_input_fifo_fifo_N1863
    );
  rx_input_fifo_fifo_BU73 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N9,
      O => rx_input_fifo_fifo_N1894
    );
  rx_input_fifo_fifo_N9_CYINIT_23 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1891,
      O => rx_input_fifo_fifo_N9_CYINIT
    );
  rx_input_fifo_fifo_N1594_LOGIC_ZERO_24 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N1594_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU150 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1594_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N1594_CYINIT,
      SEL => rx_input_fifo_fifo_N2436,
      O => rx_input_fifo_fifo_N2443
    );
  rx_input_fifo_fifo_BU149 : X_LUT4
    generic map(
      INIT => X"CA35"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1596,
      ADR1 => rx_input_fifo_fifo_N1582,
      ADR2 => rx_input_fifo_fifo_empty,
      ADR3 => rx_input_fifo_fifo_N1526,
      O => rx_input_fifo_fifo_N2436
    );
  rx_input_fifo_fifo_BU152 : X_LUT4
    generic map(
      INIT => X"99C3"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1581,
      ADR1 => rx_input_fifo_fifo_N1525,
      ADR2 => rx_input_fifo_fifo_N1595,
      ADR3 => rx_input_fifo_fifo_empty,
      O => rx_input_fifo_fifo_N2435
    );
  rx_input_fifo_fifo_N1594_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1594_CYMUXG,
      O => rx_input_fifo_fifo_N2442
    );
  rx_input_fifo_fifo_BU153 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1594_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2443,
      SEL => rx_input_fifo_fifo_N2435,
      O => rx_input_fifo_fifo_N1594_CYMUXG
    );
  rx_input_fifo_fifo_N1594_CYINIT_25 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2444,
      O => rx_input_fifo_fifo_N1594_CYINIT
    );
  rx_input_fifo_fifo_BU119 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N10,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N9,
      O => rx_input_fifo_fifo_N2372
    );
  rx_input_fifo_fifo_BU112 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N11,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_fifo_N10,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2332
    );
  rx_input_fifo_fifo_BU62 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N11,
      IB => rx_input_fifo_fifo_N11_CYINIT,
      SEL => rx_input_fifo_fifo_N1884,
      O => rx_input_fifo_fifo_N1886
    );
  rx_input_fifo_fifo_BU63 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N11_CYINIT,
      I1 => rx_input_fifo_fifo_N1884,
      O => rx_input_fifo_fifo_N1861
    );
  rx_input_fifo_fifo_BU61 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N11,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N1884
    );
  rx_input_fifo_fifo_BU67 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N10,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N1889
    );
  rx_input_fifo_fifo_N11_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N11_CYMUXG,
      O => rx_input_fifo_fifo_N1891
    );
  rx_input_fifo_fifo_BU68 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N10,
      IB => rx_input_fifo_fifo_N1886,
      SEL => rx_input_fifo_fifo_N1889,
      O => rx_input_fifo_fifo_N11_CYMUXG
    );
  rx_input_fifo_fifo_BU69 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N1886,
      I1 => rx_input_fifo_fifo_N1889,
      O => rx_input_fifo_fifo_N1862
    );
  rx_input_fifo_fifo_N11_CYINIT_26 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1881,
      O => rx_input_fifo_fifo_N11_CYINIT
    );
  rx_input_fifo_fifo_N1596_LOGIC_ZERO_27 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N1596_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU144 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1596_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N1596_CYINIT,
      SEL => rx_input_fifo_fifo_N2438,
      O => rx_input_fifo_fifo_N2445
    );
  rx_input_fifo_fifo_BU143 : X_LUT4
    generic map(
      INIT => X"C939"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1598,
      ADR1 => rx_input_fifo_fifo_N1528,
      ADR2 => rx_input_fifo_fifo_empty,
      ADR3 => rx_input_fifo_fifo_N1584,
      O => rx_input_fifo_fifo_N2438
    );
  rx_input_fifo_fifo_BU146 : X_LUT4
    generic map(
      INIT => X"B847"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1583,
      ADR1 => rx_input_fifo_fifo_empty,
      ADR2 => rx_input_fifo_fifo_N1597,
      ADR3 => rx_input_fifo_fifo_N1527,
      O => rx_input_fifo_fifo_N2437
    );
  rx_input_fifo_fifo_N1596_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1596_CYMUXG,
      O => rx_input_fifo_fifo_N2444
    );
  rx_input_fifo_fifo_BU147 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1596_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2445,
      SEL => rx_input_fifo_fifo_N2437,
      O => rx_input_fifo_fifo_N1596_CYMUXG
    );
  rx_input_fifo_fifo_N1596_CYINIT_28 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N2446,
      O => rx_input_fifo_fifo_N1596_CYINIT
    );
  rx_input_fifo_fifo_BU105 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N11,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N12,
      O => rx_input_fifo_fifo_N2292
    );
  rx_input_fifo_fifo_BU98 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N12,
      ADR2 => rx_input_fifo_fifo_N13,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2252
    );
  rx_input_fifo_fifo_BU50 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N13,
      IB => rx_input_fifo_fifo_N13_CYINIT,
      SEL => rx_input_fifo_fifo_N1874,
      O => rx_input_fifo_fifo_N1876
    );
  rx_input_fifo_fifo_BU51 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N13_CYINIT,
      I1 => rx_input_fifo_fifo_N1874,
      O => rx_input_fifo_fifo_N1859
    );
  rx_input_fifo_fifo_BU49 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N13,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N1874
    );
  rx_input_fifo_fifo_BU55 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N12,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N1879
    );
  rx_input_fifo_fifo_N13_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N13_CYMUXG,
      O => rx_input_fifo_fifo_N1881
    );
  rx_input_fifo_fifo_BU56 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N12,
      IB => rx_input_fifo_fifo_N1876,
      SEL => rx_input_fifo_fifo_N1879,
      O => rx_input_fifo_fifo_N13_CYMUXG
    );
  rx_input_fifo_fifo_BU57 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N1876,
      I1 => rx_input_fifo_fifo_N1879,
      O => rx_input_fifo_fifo_N1860
    );
  rx_input_fifo_fifo_N13_CYINIT_29 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1871,
      O => rx_input_fifo_fifo_N13_CYINIT
    );
  rx_input_fifo_fifo_N1598_LOGIC_ONE_30 : X_ONE
    port map (
      O => rx_input_fifo_fifo_N1598_LOGIC_ONE
    );
  rx_input_fifo_fifo_N1598_LOGIC_ZERO_31 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N1598_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU138 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1598_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N1598_LOGIC_ONE,
      SEL => rx_input_fifo_fifo_N2440,
      O => rx_input_fifo_fifo_N2447
    );
  rx_input_fifo_fifo_BU137 : X_LUT4
    generic map(
      INIT => X"A965"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N1530,
      ADR1 => rx_input_fifo_fifo_empty,
      ADR2 => rx_input_fifo_fifo_N1600,
      ADR3 => rx_input_fifo_fifo_N1586,
      O => rx_input_fifo_fifo_N2440
    );
  rx_input_fifo_fifo_BU140 : X_LUT4
    generic map(
      INIT => X"C693"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_empty,
      ADR1 => rx_input_fifo_fifo_N1529,
      ADR2 => rx_input_fifo_fifo_N1585,
      ADR3 => rx_input_fifo_fifo_N1599,
      O => rx_input_fifo_fifo_N2439
    );
  rx_input_fifo_fifo_N1598_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1598_CYMUXG,
      O => rx_input_fifo_fifo_N2446
    );
  rx_input_fifo_fifo_BU141 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N1598_LOGIC_ZERO,
      IB => rx_input_fifo_fifo_N2447,
      SEL => rx_input_fifo_fifo_N2439,
      O => rx_input_fifo_fifo_N1598_CYMUXG
    );
  rx_input_fifo_fifo_BU84 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N15,
      ADR1 => rx_input_fifo_fifo_N14,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N2172
    );
  rx_input_fifo_fifo_BU91 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_fifo_N14,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_fifo_N13,
      O => rx_input_fifo_fifo_N2212
    );
  rx_input_fifo_fifo_N15_LOGIC_ZERO_32 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_N15_LOGIC_ZERO
    );
  rx_input_fifo_fifo_BU38 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N15,
      IB => rx_input_fifo_fifo_N15_CYINIT,
      SEL => rx_input_fifo_fifo_N1864,
      O => rx_input_fifo_fifo_N1866
    );
  rx_input_fifo_fifo_BU39 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N15_CYINIT,
      I1 => rx_input_fifo_fifo_N1864,
      O => rx_input_fifo_fifo_N1857
    );
  rx_input_fifo_fifo_BU37 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N15,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N1864
    );
  rx_input_fifo_fifo_BU43 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_N14,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N1869
    );
  rx_input_fifo_fifo_N15_COUTUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N15_CYMUXG,
      O => rx_input_fifo_fifo_N1871
    );
  rx_input_fifo_fifo_BU44 : X_MUX2
    port map (
      IA => rx_input_fifo_fifo_N14,
      IB => rx_input_fifo_fifo_N1866,
      SEL => rx_input_fifo_fifo_N1869,
      O => rx_input_fifo_fifo_N15_CYMUXG
    );
  rx_input_fifo_fifo_BU45 : X_XOR2
    port map (
      I0 => rx_input_fifo_fifo_N1866,
      I1 => rx_input_fifo_fifo_N1869,
      O => rx_input_fifo_fifo_N1858
    );
  rx_input_fifo_fifo_N15_CYINIT_33 : X_BUF
    port map (
      I => rx_input_fifo_fifo_N15_LOGIC_ZERO,
      O => rx_input_fifo_fifo_N15_CYINIT
    );
  rx_input_fifo_fifo_BU131 : X_LUT4
    generic map(
      INIT => X"EEEE"
    )
    port map (
      ADR0 => rx_input_fifo_fifo_empty,
      ADR1 => rx_input_fifo_rd_en,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_fifo_N1599_GROM
    );
  rx_input_fifo_fifo_N1599_YUSED : X_BUF
    port map (
      I => rx_input_fifo_fifo_N1599_GROM,
      O => rx_input_fifo_fifo_N2449
    );
  rx_input_memio_n0059126_SW0 : X_LUT4
    generic map(
      INIT => X"F7FF"
    )
    port map (
      ADR0 => rx_input_memio_crcll(25),
      ADR1 => rx_input_memio_crcll(24),
      ADR2 => rx_input_memio_crcll(27),
      ADR3 => rx_input_memio_crcll(26),
      O => rx_input_memio_N80955_GROM
    );
  rx_input_memio_N80955_YUSED : X_BUF
    port map (
      I => rx_input_memio_N80955_GROM,
      O => rx_input_memio_N80955
    );
  rx_input_fifo_fifo_BU350 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1526,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1553_FFY_RST,
      O => rx_input_fifo_fifo_N1554
    );
  rx_input_fifo_fifo_N1553_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1553_FFY_RST
    );
  rx_input_memio_crcrst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcrst_FFY_RST
    );
  rx_input_memio_crcrst_34 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd16_1,
      CE => rx_input_memio_crcrst_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcrst_FFY_RST,
      O => rx_input_memio_crcrst
    );
  rx_input_memio_crcrst_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcrst_CEMUXNOT
    );
  rx_input_fifo_fifo_BU210 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2688,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N4_FFX_RST,
      O => rx_input_fifo_fifo_N4
    );
  rx_input_fifo_fifo_N4_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N4_FFX_RST
    );
  mac_control_sclkll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_sclkll_FFY_RST
    );
  mac_control_sclkll_35 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_sclkl,
      CE => mac_control_sclkll_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_sclkll_FFY_RST,
      O => mac_control_sclkll
    );
  mac_control_sclkll_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_sclkll_CEMUXNOT
    );
  mac_control_PHY_status_MII_Interface_n0077_SW18 : X_LUT4
    generic map(
      INIT => X"77FF"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(5),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(0),
      O => mac_control_PHY_status_MII_Interface_CHOICE1101_FROM
    );
  mac_control_PHY_status_MII_Interface_n0004_SW0 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(5),
      O => mac_control_PHY_status_MII_Interface_CHOICE1101_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE1101_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE1101_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE1101
    );
  mac_control_PHY_status_MII_Interface_CHOICE1101_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE1101_GROM,
      O => mac_control_PHY_status_MII_Interface_N70497
    );
  txfbbp_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => txfbbp_11_CEMUXNOT
    );
  rx_input_memio_dout_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_3_FFY_RST
    );
  rx_input_memio_dout_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_3_FFY_RST,
      O => rx_input_memio_dout(2)
    );
  txfbbp_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_13_FFY_RST
    );
  tx_output_FBBP_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(12),
      CE => txfbbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_13_FFY_RST,
      O => txfbbp(12)
    );
  txfbbp_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => txfbbp_13_CEMUXNOT
    );
  txfbbp_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_15_FFY_RST
    );
  tx_output_FBBP_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(14),
      CE => txfbbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_15_FFY_RST,
      O => txfbbp(14)
    );
  txfbbp_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => txfbbp_15_CEMUXNOT
    );
  rx_input_memio_dout_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_7_FFY_RST
    );
  rx_input_memio_dout_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_7_FFY_RST,
      O => rx_input_memio_dout(6)
    );
  mac_control_PHY_status_MII_Interface_Ker386151 : X_LUT4
    generic map(
      INIT => X"8800"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(1),
      O => mac_control_PHY_status_MII_Interface_N38617_FROM
    );
  mac_control_PHY_status_MII_Interface_sout312 : X_LUT4
    generic map(
      INIT => X"AC00"
    )
    port map (
      ADR0 => mac_control_PHY_status_din(0),
      ADR1 => mac_control_PHY_status_din(8),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR3 => mac_control_PHY_status_MII_Interface_N38617,
      O => mac_control_PHY_status_MII_Interface_N38617_GROM
    );
  mac_control_PHY_status_MII_Interface_N38617_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N38617_FROM,
      O => mac_control_PHY_status_MII_Interface_N38617
    );
  mac_control_PHY_status_MII_Interface_N38617_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N38617_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE951
    );
  rx_input_fifo_control_ldata_6_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d0(6),
      ADR1 => rx_input_fifo_control_d1(6),
      ADR2 => rx_input_fifo_control_cs_FFd1,
      ADR3 => rx_input_fifo_control_cs_FFd2,
      O => rx_input_fifo_control_CHOICE1623_FROM
    );
  rx_input_fifo_control_ldata_0_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d1(0),
      ADR1 => rx_input_fifo_control_d0(0),
      ADR2 => rx_input_fifo_control_cs_FFd1,
      ADR3 => rx_input_fifo_control_cs_FFd2,
      O => rx_input_fifo_control_CHOICE1623_GROM
    );
  rx_input_fifo_control_CHOICE1623_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1623_FROM,
      O => rx_input_fifo_control_CHOICE1623
    );
  rx_input_fifo_control_CHOICE1623_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1623_GROM,
      O => rx_input_fifo_control_CHOICE1588
    );
  rx_output_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"0A00"
    )
    port map (
      ADR0 => rx_output_nf,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_full,
      ADR3 => rx_output_cs_FFd7,
      O => rx_output_cs_FFd5_In
    );
  rx_output_cs_FFd6_In0 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_full,
      ADR3 => rx_output_cs_FFd7,
      O => rx_output_cs_FFd5_GROM
    );
  rx_output_cs_FFd5_YUSED : X_BUF
    port map (
      I => rx_output_cs_FFd5_GROM,
      O => rx_output_CHOICE1106
    );
  rx_input_fifo_control_ldata_8_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_d1(8),
      ADR1 => rx_input_fifo_control_cs_FFd2,
      ADR2 => rx_input_fifo_control_d0(8),
      ADR3 => rx_input_fifo_control_cs_FFd1,
      O => rx_input_fifo_control_CHOICE1602_FROM
    );
  rx_input_fifo_control_ldata_1_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d1(1),
      ADR1 => rx_input_fifo_control_d0(1),
      ADR2 => rx_input_fifo_control_cs_FFd2,
      ADR3 => rx_input_fifo_control_cs_FFd1,
      O => rx_input_fifo_control_CHOICE1602_GROM
    );
  rx_input_fifo_control_CHOICE1602_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1602_FROM,
      O => rx_input_fifo_control_CHOICE1602
    );
  rx_input_fifo_control_CHOICE1602_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1602_GROM,
      O => rx_input_fifo_control_CHOICE1581
    );
  rx_input_fifo_control_ldata_0_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd4,
      ADR1 => rx_input_fifo_control_d3(0),
      ADR2 => rx_input_fifo_control_d2(0),
      ADR3 => rx_input_fifo_control_cs_FFd3,
      O => rx_input_data_0_FROM
    );
  rx_input_fifo_control_ldata_0_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1588,
      ADR3 => rx_input_fifo_control_CHOICE1591,
      O => rx_input_fifo_control_ldata(0)
    );
  rx_input_data_0_XUSED : X_BUF
    port map (
      I => rx_input_data_0_FROM,
      O => rx_input_fifo_control_CHOICE1591
    );
  rx_input_fifo_control_ldata_4_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd2,
      ADR1 => rx_input_fifo_control_d1(4),
      ADR2 => rx_input_fifo_control_d0(4),
      ADR3 => rx_input_fifo_control_cs_FFd1,
      O => rx_input_fifo_control_CHOICE1630_FROM
    );
  rx_input_fifo_control_ldata_2_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd2,
      ADR1 => rx_input_fifo_control_cs_FFd1,
      ADR2 => rx_input_fifo_control_d1(2),
      ADR3 => rx_input_fifo_control_d0(2),
      O => rx_input_fifo_control_CHOICE1630_GROM
    );
  rx_input_fifo_control_CHOICE1630_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1630_FROM,
      O => rx_input_fifo_control_CHOICE1630
    );
  rx_input_fifo_control_CHOICE1630_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1630_GROM,
      O => rx_input_fifo_control_CHOICE1644
    );
  rx_input_fifo_control_ldata_1_9 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd4,
      ADR1 => rx_input_fifo_control_cs_FFd3,
      ADR2 => rx_input_fifo_control_d2(1),
      ADR3 => rx_input_fifo_control_d3(1),
      O => rx_input_data_1_FROM
    );
  rx_input_fifo_control_ldata_1_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1581,
      ADR3 => rx_input_fifo_control_CHOICE1584,
      O => rx_input_fifo_control_ldata(1)
    );
  rx_input_data_1_XUSED : X_BUF
    port map (
      I => rx_input_data_1_FROM,
      O => rx_input_fifo_control_CHOICE1584
    );
  tx_output_n000724 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcnt_44,
      ADR1 => tx_output_bcnt_45,
      ADR2 => tx_output_bcnt_43,
      ADR3 => tx_output_bcnt_42,
      O => tx_output_CHOICE1871_GROM
    );
  tx_output_CHOICE1871_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1871_GROM,
      O => tx_output_CHOICE1871
    );
  rx_input_fifo_control_ldata_9_4 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd1,
      ADR1 => rx_input_fifo_control_d0(9),
      ADR2 => rx_input_fifo_control_d1(9),
      ADR3 => rx_input_fifo_control_cs_FFd2,
      O => rx_input_fifo_control_CHOICE1595_FROM
    );
  rx_input_fifo_control_ldata_3_4 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d0(3),
      ADR1 => rx_input_fifo_control_cs_FFd2,
      ADR2 => rx_input_fifo_control_cs_FFd1,
      ADR3 => rx_input_fifo_control_d1(3),
      O => rx_input_fifo_control_CHOICE1595_GROM
    );
  rx_input_fifo_control_CHOICE1595_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1595_FROM,
      O => rx_input_fifo_control_CHOICE1595
    );
  rx_input_fifo_control_CHOICE1595_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1595_GROM,
      O => rx_input_fifo_control_CHOICE1637
    );
  rx_input_fifo_control_ldata_2_9 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd4,
      ADR1 => rx_input_fifo_control_cs_FFd3,
      ADR2 => rx_input_fifo_control_d3(2),
      ADR3 => rx_input_fifo_control_d2(2),
      O => rx_input_data_2_FROM
    );
  rx_input_fifo_control_ldata_2_10 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_fifo_control_CHOICE1644,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_control_CHOICE1647,
      O => rx_input_fifo_control_ldata(2)
    );
  rx_input_data_2_XUSED : X_BUF
    port map (
      I => rx_input_data_2_FROM,
      O => rx_input_fifo_control_CHOICE1647
    );
  rx_input_fifo_fifo_BU287 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1525,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1539_FFX_RST,
      O => rx_input_fifo_fifo_N1539
    );
  rx_input_fifo_fifo_N1539_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1539_FFX_RST
    );
  tx_output_bcnt_inst_sum_186_36 : X_XOR2
    port map (
      I0 => tx_output_bcnt_53_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_55,
      O => tx_output_bcnt_inst_sum_186
    );
  tx_output_bcnt_inst_lut3_551 : X_LUT4
    generic map(
      INIT => X"0C3F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => q2(15),
      ADR3 => tx_output_bcnt_53,
      O => tx_output_bcnt_inst_lut3_55
    );
  tx_output_n000761 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcnt_52,
      ADR1 => tx_output_bcnt_50,
      ADR2 => tx_output_bcnt_53,
      ADR3 => tx_output_bcnt_51,
      O => tx_output_bcnt_53_GROM
    );
  tx_output_bcnt_53_YUSED : X_BUF
    port map (
      I => tx_output_bcnt_53_GROM,
      O => tx_output_CHOICE1886
    );
  tx_output_bcnt_53_CYINIT_37 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_219,
      O => tx_output_bcnt_53_CYINIT
    );
  rx_input_fifo_control_ldata_3_9 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d3(3),
      ADR1 => rx_input_fifo_control_d2(3),
      ADR2 => rx_input_fifo_control_cs_FFd3,
      ADR3 => rx_input_fifo_control_cs_FFd4,
      O => rx_input_data_3_FROM
    );
  rx_input_fifo_control_ldata_3_10 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_control_CHOICE1637,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_control_CHOICE1640,
      O => rx_input_fifo_control_ldata(3)
    );
  rx_input_data_3_XUSED : X_BUF
    port map (
      I => rx_input_data_3_FROM,
      O => rx_input_fifo_control_CHOICE1640
    );
  tx_output_n000748 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcnt_46,
      ADR1 => tx_output_bcnt_49,
      ADR2 => tx_output_bcnt_47,
      ADR3 => tx_output_bcnt_48,
      O => tx_output_CHOICE1879_GROM
    );
  tx_output_CHOICE1879_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1879_GROM,
      O => tx_output_CHOICE1879
    );
  rx_input_fifo_control_ldata_7_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd1,
      ADR1 => rx_input_fifo_control_d1(7),
      ADR2 => rx_input_fifo_control_cs_FFd2,
      ADR3 => rx_input_fifo_control_d0(7),
      O => rx_input_fifo_control_CHOICE1609_FROM
    );
  rx_input_fifo_control_ldata_5_4 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d0(5),
      ADR1 => rx_input_fifo_control_d1(5),
      ADR2 => rx_input_fifo_control_cs_FFd2,
      ADR3 => rx_input_fifo_control_cs_FFd1,
      O => rx_input_fifo_control_CHOICE1609_GROM
    );
  rx_input_fifo_control_CHOICE1609_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1609_FROM,
      O => rx_input_fifo_control_CHOICE1609
    );
  rx_input_fifo_control_CHOICE1609_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1609_GROM,
      O => rx_input_fifo_control_CHOICE1616
    );
  tx_output_n000774 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => tx_output_CHOICE1879,
      ADR1 => tx_output_CHOICE1886,
      ADR2 => tx_output_N80951,
      ADR3 => tx_output_CHOICE1871,
      O => tx_output_cs_FFd4_FROM
    );
  tx_output_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => tx_output_cs_FFd5_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_n0007,
      O => tx_output_cs_FFd4_GROM
    );
  tx_output_cs_FFd4_XUSED : X_BUF
    port map (
      I => tx_output_cs_FFd4_FROM,
      O => tx_output_n0007
    );
  tx_output_cs_FFd4_YUSED : X_BUF
    port map (
      I => tx_output_cs_FFd4_GROM,
      O => tx_output_cs_FFd4_In
    );
  rx_input_fifo_control_ldata_4_9 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d2(4),
      ADR1 => rx_input_fifo_control_d3(4),
      ADR2 => rx_input_fifo_control_cs_FFd3,
      ADR3 => rx_input_fifo_control_cs_FFd4,
      O => rx_input_data_4_FROM
    );
  rx_input_fifo_control_ldata_4_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1630,
      ADR3 => rx_input_fifo_control_CHOICE1633,
      O => rx_input_fifo_control_ldata(4)
    );
  rx_input_data_4_XUSED : X_BUF
    port map (
      I => rx_input_data_4_FROM,
      O => rx_input_fifo_control_CHOICE1633
    );
  rx_input_fifo_control_ldata_5_9 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_fifo_control_d2(5),
      ADR1 => rx_input_fifo_control_cs_FFd4,
      ADR2 => rx_input_fifo_control_cs_FFd3,
      ADR3 => rx_input_fifo_control_d3(5),
      O => rx_input_data_5_FROM
    );
  rx_input_fifo_control_ldata_5_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1616,
      ADR3 => rx_input_fifo_control_CHOICE1619,
      O => rx_input_fifo_control_ldata(5)
    );
  rx_input_data_5_XUSED : X_BUF
    port map (
      I => rx_input_data_5_FROM,
      O => rx_input_fifo_control_CHOICE1619
    );
  rx_input_fifo_control_ldata_6_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_d3(6),
      ADR1 => rx_input_fifo_control_cs_FFd4,
      ADR2 => rx_input_fifo_control_cs_FFd3,
      ADR3 => rx_input_fifo_control_d2(6),
      O => rx_input_data_6_FROM
    );
  rx_input_fifo_control_ldata_6_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1623,
      ADR3 => rx_input_fifo_control_CHOICE1626,
      O => rx_input_fifo_control_ldata(6)
    );
  rx_input_data_6_XUSED : X_BUF
    port map (
      I => rx_input_data_6_FROM,
      O => rx_input_fifo_control_CHOICE1626
    );
  rx_input_fifo_control_ldata_7_9 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd4,
      ADR1 => rx_input_fifo_control_d2(7),
      ADR2 => rx_input_fifo_control_cs_FFd3,
      ADR3 => rx_input_fifo_control_d3(7),
      O => rx_input_data_7_FROM
    );
  rx_input_fifo_control_ldata_7_10 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_CHOICE1609,
      ADR3 => rx_input_fifo_control_CHOICE1612,
      O => rx_input_fifo_control_ldata(7)
    );
  rx_input_data_7_XUSED : X_BUF
    port map (
      I => rx_input_data_7_FROM,
      O => rx_input_fifo_control_CHOICE1612
    );
  rx_input_fifo_control_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_ce,
      ADR2 => rx_input_fifo_control_cs_FFd4,
      ADR3 => VCC,
      O => rx_input_fifo_control_cs_FFd3_In
    );
  rx_input_fifo_control_ldata_8_9 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => rx_input_fifo_control_d2(8),
      ADR1 => rx_input_fifo_control_cs_FFd3,
      ADR2 => rx_input_fifo_control_d3(8),
      ADR3 => rx_input_fifo_control_cs_FFd4,
      O => rx_input_fifo_control_cs_FFd3_GROM
    );
  rx_input_fifo_control_cs_FFd3_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_cs_FFd3_GROM,
      O => rx_input_fifo_control_CHOICE1605
    );
  rx_input_fifo_control_ldata_9_9 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd4,
      ADR1 => rx_input_fifo_control_d2(9),
      ADR2 => rx_input_fifo_control_cs_FFd3,
      ADR3 => rx_input_fifo_control_d3(9),
      O => rx_input_fifo_control_CHOICE1598_FROM
    );
  rx_input_fifo_control_ldata_9_10 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_control_CHOICE1595,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_control_CHOICE1598,
      O => rx_input_fifo_control_CHOICE1598_GROM
    );
  rx_input_fifo_control_CHOICE1598_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1598_FROM,
      O => rx_input_fifo_control_CHOICE1598
    );
  rx_input_fifo_control_CHOICE1598_YUSED : X_BUF
    port map (
      I => rx_input_fifo_control_CHOICE1598_GROM,
      O => rx_input_fifo_control_ldata(9)
    );
  rx_output_Ker344841 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_cs_FFd11,
      ADR2 => rx_output_cs_FFd1,
      ADR3 => VCC,
      O => rx_output_cs_FFd9_FROM
    );
  rx_output_cs_FFd9_In1 : X_LUT4
    generic map(
      INIT => X"AA08"
    )
    port map (
      ADR0 => rx_output_nf,
      ADR1 => rx_output_cs_FFd5,
      ADR2 => rx_output_n0018,
      ADR3 => rx_output_N34486,
      O => rx_output_cs_FFd9_In
    );
  rx_output_cs_FFd9_XUSED : X_BUF
    port map (
      I => rx_output_cs_FFd9_FROM,
      O => rx_output_N34486
    );
  tx_output_crc_loigc_Mxor_CO_6_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_Mxor_n0007_Xo(0),
      ADR1 => tx_output_crc_loigc_Mxor_CO_18_Xo(0),
      ADR2 => tx_output_crc_loigc_n0115(0),
      ADR3 => tx_output_crc_loigc_n0124(0),
      O => tx_output_crcl_6_FROM
    );
  tx_output_n0034_6_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_6_Q,
      O => tx_output_n0034_6_1_O
    );
  tx_output_crcl_6_XUSED : X_BUF
    port map (
      I => tx_output_crcl_6_FROM,
      O => tx_output_crc_6_Q
    );
  mac_control_Ker53107 : X_LUT4
    generic map(
      INIT => X"0080"
    )
    port map (
      ADR0 => mac_control_addr(3),
      ADR1 => mac_control_sclkdeltal,
      ADR2 => mac_control_addr(4),
      ADR3 => mac_control_N69572,
      O => mac_control_N53109_FROM
    );
  mac_control_n00281 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => mac_control_addr_0_1,
      ADR1 => mac_control_addr(2),
      ADR2 => mac_control_addr(1),
      ADR3 => mac_control_N53109,
      O => mac_control_N53109_GROM
    );
  mac_control_N53109_XUSED : X_BUF
    port map (
      I => mac_control_N53109_FROM,
      O => mac_control_N53109
    );
  mac_control_N53109_YUSED : X_BUF
    port map (
      I => mac_control_N53109_GROM,
      O => mac_control_n0028
    );
  mac_control_Ker53142 : X_LUT4
    generic map(
      INIT => X"0008"
    )
    port map (
      ADR0 => mac_control_N53132,
      ADR1 => mac_control_addr(0),
      ADR2 => mac_control_addr(3),
      ADR3 => mac_control_N69759,
      O => mac_control_N53144_FROM
    );
  mac_control_n00331 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_N53144,
      O => mac_control_N53144_GROM
    );
  mac_control_N53144_XUSED : X_BUF
    port map (
      I => mac_control_N53144_FROM,
      O => mac_control_N53144
    );
  mac_control_N53144_YUSED : X_BUF
    port map (
      I => mac_control_N53144_GROM,
      O => mac_control_n0033
    );
  mac_control_PHY_status_MII_Interface_n0004_38 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(1),
      ADR1 => mac_control_PHY_status_MII_Interface_N70497,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(2),
      O => mac_control_PHY_status_MII_Interface_cs_FFd2_FROM
    );
  mac_control_PHY_status_MII_Interface_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_n0004,
      O => mac_control_PHY_status_MII_Interface_cs_FFd2_In
    );
  mac_control_PHY_status_MII_Interface_cs_FFd2_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd2_FROM,
      O => mac_control_PHY_status_MII_Interface_n0004
    );
  macaddr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_3_FFY_RST
    );
  mac_control_MACADDR_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_3_FFY_RST,
      O => macaddr(2)
    );
  macaddr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_5_FFY_RST
    );
  mac_control_MACADDR_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_5_FFY_RST,
      O => macaddr(4)
    );
  macaddr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_9_FFY_RST
    );
  mac_control_MACADDR_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_9_FFY_RST,
      O => macaddr(8)
    );
  tx_output_crc_loigc_Mxor_n0001_Result1 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_crcl(24),
      ADR2 => VCC,
      ADR3 => tx_output_data(7),
      O => tx_output_crc_loigc_n0122_1_FROM
    );
  tx_output_crc_loigc_Mxor_CO_7_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(7),
      ADR1 => tx_output_data(4),
      ADR2 => tx_output_crcl(27),
      ADR3 => tx_output_crcl(24),
      O => tx_output_crc_loigc_n0122_1_GROM
    );
  tx_output_crc_loigc_n0122_1_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0122_1_FROM,
      O => tx_output_crc_loigc_n0122(1)
    );
  tx_output_crc_loigc_n0122_1_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0122_1_GROM,
      O => tx_output_crc_loigc_Mxor_CO_7_Xo(1)
    );
  rx_input_fifo_fifo_BU309 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1540,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1547_FFX_RST,
      O => rx_input_fifo_fifo_N1547
    );
  rx_input_fifo_fifo_N1547_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1547_FFX_RST
    );
  tx_output_crc_loigc_Mxor_CO_7_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0118(0),
      ADR1 => tx_output_crc_loigc_n0118(1),
      ADR2 => tx_output_crc_loigc_Mxor_CO_7_Xo(1),
      ADR3 => tx_output_crc_loigc_n0124(0),
      O => tx_output_crcl_7_FROM
    );
  tx_output_n0034_7_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16_1,
      ADR3 => tx_output_crc_7_Q,
      O => tx_output_n0034_7_Q
    );
  tx_output_crcl_7_XUSED : X_BUF
    port map (
      I => tx_output_crcl_7_FROM,
      O => tx_output_crc_7_Q
    );
  tx_input_Ker35859120_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_input_CNT(1),
      ADR1 => tx_input_CNT(2),
      ADR2 => tx_input_CNT(0),
      ADR3 => tx_input_CNT(3),
      O => tx_input_N80947_FROM
    );
  tx_input_Ker358594 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => tx_input_CNT(1),
      ADR1 => tx_input_CNT(3),
      ADR2 => tx_input_CNT(0),
      ADR3 => tx_input_CNT(2),
      O => tx_input_N80947_GROM
    );
  tx_input_N80947_XUSED : X_BUF
    port map (
      I => tx_input_N80947_FROM,
      O => tx_input_N80947
    );
  tx_input_N80947_YUSED : X_BUF
    port map (
      I => tx_input_N80947_GROM,
      O => tx_input_CHOICE1988
    );
  tx_input_Ker3585970 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_input_CNT(5),
      ADR1 => tx_input_CNT(7),
      ADR2 => tx_input_CNT(6),
      ADR3 => tx_input_CNT(4),
      O => tx_input_CHOICE2014_FROM
    );
  tx_input_Ker358599 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => tx_input_CNT(7),
      ADR1 => tx_input_CNT(5),
      ADR2 => tx_input_CNT(4),
      ADR3 => tx_input_CNT(6),
      O => tx_input_CHOICE2014_GROM
    );
  tx_input_CHOICE2014_XUSED : X_BUF
    port map (
      I => tx_input_CHOICE2014_FROM,
      O => tx_input_CHOICE2014
    );
  tx_input_CHOICE2014_YUSED : X_BUF
    port map (
      I => tx_input_CHOICE2014_GROM,
      O => tx_input_CHOICE1991
    );
  mac_control_Mmux_n0016_Result_1_97_SW1 : X_LUT4
    generic map(
      INIT => X"FF15"
    )
    port map (
      ADR0 => mac_control_CHOICE2625,
      ADR1 => mac_control_phydo(1),
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_addr(5),
      O => mac_control_dout_1_FROM
    );
  mac_control_Mmux_n0016_Result_1_97 : X_LUT4
    generic map(
      INIT => X"70F8"
    )
    port map (
      ADR0 => mac_control_sclkdeltall,
      ADR1 => mac_control_n0086,
      ADR2 => mac_control_dout(0),
      ADR3 => mac_control_N81427,
      O => mac_control_n0016(1)
    );
  mac_control_dout_1_XUSED : X_BUF
    port map (
      I => mac_control_dout_1_FROM,
      O => mac_control_N81427
    );
  mac_control_PHY_status_din_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_1_FFY_RST
    );
  mac_control_PHY_status_din_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(0),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_1_FFY_RST,
      O => mac_control_PHY_status_din(0)
    );
  mac_control_PHY_status_din_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_5_FFY_RST
    );
  mac_control_PHY_status_din_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(4),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_5_FFY_RST,
      O => mac_control_PHY_status_din(4)
    );
  rx_input_fifo_fifo_BU352 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1525,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1553_FFX_RST,
      O => rx_input_fifo_fifo_N1553
    );
  rx_input_fifo_fifo_N1553_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1553_FFX_RST
    );
  mac_control_PHY_status_din_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_7_FFY_RST
    );
  mac_control_PHY_status_din_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(6),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_7_FFY_RST,
      O => mac_control_PHY_status_din(6)
    );
  mac_control_rxfifowerr_cntl_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_10_FFY_RST
    );
  mac_control_rxfifowerr_cntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(10),
      CE => mac_control_rxfifowerr_cntl_10_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_10_FFY_RST,
      O => mac_control_rxfifowerr_cntl(10)
    );
  mac_control_rxfifowerr_cntl_10_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_10_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_11_FFY_RST
    );
  mac_control_rxfifowerr_cntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(11),
      CE => mac_control_rxfifowerr_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_11_FFY_RST,
      O => mac_control_rxfifowerr_cntl(11)
    );
  mac_control_rxfifowerr_cntl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_11_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_21_FFY_RST
    );
  mac_control_rxfifowerr_cntl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(20),
      CE => mac_control_rxfifowerr_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_21_FFY_RST,
      O => mac_control_rxfifowerr_cntl(20)
    );
  mac_control_rxfifowerr_cntl_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_21_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_13_FFY_RST
    );
  mac_control_rxfifowerr_cntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(12),
      CE => mac_control_rxfifowerr_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_13_FFY_RST,
      O => mac_control_rxfifowerr_cntl(12)
    );
  mac_control_rxfifowerr_cntl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_13_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_31_FFY_RST
    );
  mac_control_rxfifowerr_cntl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(30),
      CE => mac_control_rxfifowerr_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_31_FFY_RST,
      O => mac_control_rxfifowerr_cntl(30)
    );
  mac_control_rxfifowerr_cntl_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_31_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_23_FFY_RST
    );
  mac_control_rxfifowerr_cntl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(22),
      CE => mac_control_rxfifowerr_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_23_FFY_RST,
      O => mac_control_rxfifowerr_cntl(22)
    );
  mac_control_rxfifowerr_cntl_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_23_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_15_FFY_RST
    );
  mac_control_rxfifowerr_cntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(14),
      CE => mac_control_rxfifowerr_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_15_FFY_RST,
      O => mac_control_rxfifowerr_cntl(14)
    );
  mac_control_rxfifowerr_cntl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_15_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_25_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_17_FFY_RST
    );
  mac_control_rxfifowerr_cntl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(16),
      CE => mac_control_rxfifowerr_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_17_FFY_RST,
      O => mac_control_rxfifowerr_cntl(16)
    );
  mac_control_rxfifowerr_cntl_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_17_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_27_FFY_RST
    );
  mac_control_rxfifowerr_cntl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(26),
      CE => mac_control_rxfifowerr_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_27_FFY_RST,
      O => mac_control_rxfifowerr_cntl(26)
    );
  mac_control_rxfifowerr_cntl_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_27_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_19_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_29_FFY_RST
    );
  mac_control_rxfifowerr_cntl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(28),
      CE => mac_control_rxfifowerr_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_29_FFY_RST,
      O => mac_control_rxfifowerr_cntl(28)
    );
  mac_control_rxfifowerr_cntl_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_29_CEMUXNOT
    );
  mac_control_dout_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_2_FFY_RST
    );
  mac_control_dout_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(2),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_2_FFY_RST,
      O => mac_control_dout(2)
    );
  mac_control_Mmux_n0016_Result_2_97_SW1 : X_LUT4
    generic map(
      INIT => X"FF07"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_phydo(2),
      ADR2 => mac_control_CHOICE2651,
      ADR3 => mac_control_addr(5),
      O => mac_control_dout_2_FROM
    );
  mac_control_Mmux_n0016_Result_2_97 : X_LUT4
    generic map(
      INIT => X"2AEA"
    )
    port map (
      ADR0 => mac_control_dout(1),
      ADR1 => mac_control_n0086,
      ADR2 => mac_control_sclkdeltall,
      ADR3 => mac_control_N81431,
      O => mac_control_n0016(2)
    );
  mac_control_dout_2_XUSED : X_BUF
    port map (
      I => mac_control_dout_2_FROM,
      O => mac_control_N81431
    );
  rx_input_memio_crccomb_Mxor_CO_18_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_datal(1),
      ADR1 => rx_input_memio_crcl(26),
      ADR2 => rx_input_memio_crcl(30),
      ADR3 => rx_input_memio_datal(5),
      O => rx_input_memio_crccomb_Mxor_CO_18_Xo_0_FROM
    );
  rx_input_memio_crccomb_Mxor_n0000_Result1 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_input_memio_datal(1),
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcl(30),
      ADR3 => VCC,
      O => rx_input_memio_crccomb_Mxor_CO_18_Xo_0_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_18_Xo_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_18_Xo_0_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_18_Xo(0)
    );
  rx_input_memio_crccomb_Mxor_CO_18_Xo_0_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_18_Xo_0_GROM,
      O => rx_input_memio_crccomb_n0104(0)
    );
  tx_input_fifofulll_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_fifofulll_CEMUXNOT
    );
  rx_input_fifo_fifo_BU336 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1574_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1574
    );
  rx_input_fifo_fifo_N1574_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1574_FFX_SET
    );
  mac_control_dout_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_3_FFY_RST
    );
  mac_control_dout_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(3),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_3_FFY_RST,
      O => mac_control_dout(3)
    );
  mac_control_Mmux_n0016_Result_3_93_SW1 : X_LUT4
    generic map(
      INIT => X"CDDD"
    )
    port map (
      ADR0 => mac_control_CHOICE2449,
      ADR1 => mac_control_addr(5),
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_phydo(3),
      O => mac_control_dout_3_FROM
    );
  mac_control_Mmux_n0016_Result_3_93 : X_LUT4
    generic map(
      INIT => X"70F8"
    )
    port map (
      ADR0 => mac_control_n0086,
      ADR1 => mac_control_sclkdeltall,
      ADR2 => mac_control_dout(2),
      ADR3 => mac_control_N81435,
      O => mac_control_n0016(3)
    );
  mac_control_dout_3_XUSED : X_BUF
    port map (
      I => mac_control_dout_3_FROM,
      O => mac_control_N81435
    );
  tx_output_crc_loigc_Mxor_CO_8_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0122(0),
      ADR1 => tx_output_crc_loigc_Mxor_CO_7_Xo(1),
      ADR2 => tx_output_crcl(0),
      ADR3 => tx_output_crc_loigc_n0115(0),
      O => tx_output_crcl_8_FROM
    );
  tx_output_n0034_8_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16_1,
      ADR3 => tx_output_crc_8_Q,
      O => tx_output_n0034_8_1_O
    );
  tx_output_crcl_8_XUSED : X_BUF
    port map (
      I => tx_output_crcl_8_FROM,
      O => tx_output_crc_8_Q
    );
  mac_control_CLKSL_5_39 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => clksl,
      O => mac_control_CLKSL_5_FROM
    );
  mac_control_CLKSL_1_40 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => clksl,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_CLKSL_5_GROM
    );
  mac_control_CLKSL_5_XUSED : X_BUF
    port map (
      I => mac_control_CLKSL_5_FROM,
      O => mac_control_CLKSL_5
    );
  mac_control_CLKSL_5_YUSED : X_BUF
    port map (
      I => mac_control_CLKSL_5_GROM,
      O => mac_control_CLKSL_1
    );
  mac_control_CLKSL_4_41 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => clksl,
      ADR3 => VCC,
      O => mac_control_CLKSL_4_FROM
    );
  mac_control_CLKSL_2_42 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => clksl,
      ADR3 => VCC,
      O => mac_control_CLKSL_4_GROM
    );
  mac_control_CLKSL_4_XUSED : X_BUF
    port map (
      I => mac_control_CLKSL_4_FROM,
      O => mac_control_CLKSL_4
    );
  mac_control_CLKSL_4_YUSED : X_BUF
    port map (
      I => mac_control_CLKSL_4_GROM,
      O => mac_control_CLKSL_2
    );
  mac_control_CLKSL_3_43 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => clksl,
      ADR3 => VCC,
      O => mac_control_CLKSL_3_GROM
    );
  mac_control_CLKSL_3_YUSED : X_BUF
    port map (
      I => mac_control_CLKSL_3_GROM,
      O => mac_control_CLKSL_3
    );
  rx_input_memio_n0059100 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => rx_input_memio_crcll(18),
      ADR1 => rx_input_memio_crcll(17),
      ADR2 => rx_input_memio_crcll(19),
      ADR3 => rx_input_memio_crcll(16),
      O => rx_input_memio_CHOICE1839_GROM
    );
  rx_input_memio_CHOICE1839_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1839_GROM,
      O => rx_input_memio_CHOICE1839
    );
  rx_input_memio_n0059113 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_input_memio_crcll(20),
      ADR1 => rx_input_memio_crcll(21),
      ADR2 => rx_input_memio_crcll(22),
      ADR3 => rx_input_memio_crcll(23),
      O => rx_input_memio_CHOICE1846_GROM
    );
  rx_input_memio_CHOICE1846_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1846_GROM,
      O => rx_input_memio_CHOICE1846
    );
  rx_input_memio_n0059126 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => rx_input_memio_CHOICE1839,
      ADR1 => rx_input_memio_CHOICE1846,
      ADR2 => rx_input_memio_N80955,
      ADR3 => rx_input_memio_CHOICE1832,
      O => rx_input_memio_crcequal_FROM
    );
  rx_input_memio_n0059141 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_CHOICE1812,
      ADR1 => rx_input_memio_CHOICE1808,
      ADR2 => rx_input_memio_CHOICE1822,
      ADR3 => rx_input_memio_CHOICE1848,
      O => rx_input_memio_n0059
    );
  rx_input_memio_crcequal_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcequal_CEMUXNOT
    );
  rx_input_memio_crcequal_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcequal_FROM,
      O => rx_input_memio_CHOICE1848
    );
  rx_input_fifo_fifo_BU408 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3688,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1560_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1561
    );
  rx_input_fifo_fifo_N1560_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1560_FFY_SET
    );
  rx_input_memio_n00331 : X_LUT4
    generic map(
      INIT => X"000C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_men,
      ADR2 => rx_input_memio_RESET_1,
      ADR3 => rx_input_memio_menl,
      O => rx_input_memio_n0033_FROM
    );
  rx_input_memio_n00331_1_44 : X_LUT4
    generic map(
      INIT => X"0404"
    )
    port map (
      ADR0 => rx_input_memio_menl,
      ADR1 => rx_input_memio_men,
      ADR2 => rx_input_RESET_1,
      ADR3 => VCC,
      O => rx_input_memio_n0033_GROM
    );
  rx_input_memio_n0033_XUSED : X_BUF
    port map (
      I => rx_input_memio_n0033_FROM,
      O => rx_input_memio_n0033
    );
  rx_input_memio_n0033_YUSED : X_BUF
    port map (
      I => rx_input_memio_n0033_GROM,
      O => rx_input_memio_n00331_1
    );
  mac_control_Mmux_n0016_Result_4_93_SW1 : X_LUT4
    generic map(
      INIT => X"CDCF"
    )
    port map (
      ADR0 => mac_control_phydo(4),
      ADR1 => mac_control_addr(5),
      ADR2 => mac_control_CHOICE2424,
      ADR3 => mac_control_n0060,
      O => mac_control_dout_4_FROM
    );
  mac_control_Mmux_n0016_Result_4_93 : X_LUT4
    generic map(
      INIT => X"4CEC"
    )
    port map (
      ADR0 => mac_control_n0086,
      ADR1 => mac_control_dout(3),
      ADR2 => mac_control_sclkdeltall,
      ADR3 => mac_control_N81439,
      O => mac_control_n0016(4)
    );
  mac_control_dout_4_XUSED : X_BUF
    port map (
      I => mac_control_dout_4_FROM,
      O => mac_control_N81439
    );
  rx_input_memio_crccomb_Mxor_CO_23_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_datal(6),
      ADR1 => rx_input_memio_datal(7),
      ADR2 => rx_input_memio_crcl(25),
      ADR3 => rx_input_memio_crcl(24),
      O => rx_input_memio_crccomb_Mxor_CO_23_Xo_0_FROM
    );
  rx_input_memio_crccomb_Mxor_n0001_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcl(24),
      ADR3 => rx_input_memio_datal(7),
      O => rx_input_memio_crccomb_Mxor_CO_23_Xo_0_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_23_Xo_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_23_Xo_0_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_23_Xo(0)
    );
  rx_input_memio_crccomb_Mxor_CO_23_Xo_0_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_23_Xo_0_GROM,
      O => rx_input_memio_crccomb_n0122(1)
    );
  tx_output_crc_loigc_Mxor_CO_18_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(5),
      ADR1 => tx_output_crcl(26),
      ADR2 => tx_output_data(1),
      ADR3 => tx_output_crcl(30),
      O => tx_output_crc_loigc_Mxor_CO_18_Xo_0_FROM
    );
  tx_output_crc_loigc_Mxor_n0000_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_crcl(30),
      ADR3 => tx_output_data(1),
      O => tx_output_crc_loigc_Mxor_CO_18_Xo_0_GROM
    );
  tx_output_crc_loigc_Mxor_CO_18_Xo_0_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_18_Xo_0_FROM,
      O => tx_output_crc_loigc_Mxor_CO_18_Xo(0)
    );
  tx_output_crc_loigc_Mxor_CO_18_Xo_0_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_18_Xo_0_GROM,
      O => tx_output_crc_loigc_n0104(0)
    );
  tx_output_crc_loigc_Mxor_n0012_Result1 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => tx_output_data(6),
      ADR1 => VCC,
      ADR2 => tx_output_crcl(25),
      ADR3 => VCC,
      O => tx_output_crc_loigc_n0122_0_FROM
    );
  tx_output_crc_loigc_Mxor_CO_9_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(28),
      ADR1 => tx_output_data(6),
      ADR2 => tx_output_data(3),
      ADR3 => tx_output_crcl(25),
      O => tx_output_crc_loigc_n0122_0_GROM
    );
  tx_output_crc_loigc_n0122_0_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0122_0_FROM,
      O => tx_output_crc_loigc_n0122(0)
    );
  tx_output_crc_loigc_n0122_0_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0122_0_GROM,
      O => tx_output_crc_loigc_Mxor_CO_9_Xo(0)
    );
  rx_output_fifo_nearfull_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifo_nearfull_CEMUXNOT
    );
  tx_output_crcl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_9_FFY_RST
    );
  tx_output_crcl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_9_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_9_FFY_RST,
      O => tx_output_crcl(9)
    );
  tx_output_crc_loigc_Mxor_CO_9_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0118(0),
      ADR1 => tx_output_crc_loigc_Mxor_CO_9_Xo(0),
      ADR2 => tx_output_crcl(1),
      ADR3 => tx_output_crc_loigc_n0118(1),
      O => tx_output_crcl_9_FROM
    );
  tx_output_n0034_9_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_9_Q,
      O => tx_output_n0034_9_Q
    );
  tx_output_crcl_9_XUSED : X_BUF
    port map (
      I => tx_output_crcl_9_FROM,
      O => tx_output_crc_9_Q
    );
  mac_control_Mmux_n0016_Result_5_97_SW1 : X_LUT4
    generic map(
      INIT => X"ABBB"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_CHOICE2677,
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_phydo(5),
      O => mac_control_dout_5_FROM
    );
  mac_control_Mmux_n0016_Result_5_97 : X_LUT4
    generic map(
      INIT => X"2AEA"
    )
    port map (
      ADR0 => mac_control_dout(4),
      ADR1 => mac_control_n0086,
      ADR2 => mac_control_sclkdeltall,
      ADR3 => mac_control_N81443,
      O => mac_control_n0016(5)
    );
  mac_control_dout_5_XUSED : X_BUF
    port map (
      I => mac_control_dout_5_FROM,
      O => mac_control_N81443
    );
  addr4ext_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_5_FFY_RST
    );
  tx_input_MA_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_20,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_5_FFY_RST,
      O => addr4ext(4)
    );
  addr4ext_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_7_FFY_RST
    );
  tx_input_MA_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_22,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_7_FFY_RST,
      O => addr4ext(6)
    );
  addr4ext_9_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_9_FFY_RST
    );
  tx_input_MA_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_24,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_9_FFY_RST,
      O => addr4ext(8)
    );
  d4_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_3_FFY_RST
    );
  tx_input_MD_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(2),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_3_FFY_RST,
      O => d4(2)
    );
  d4_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_5_FFY_RST
    );
  tx_input_MD_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(4),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_5_FFY_RST,
      O => d4(4)
    );
  d4_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_7_FFY_RST
    );
  tx_input_MD_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(6),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_7_FFY_RST,
      O => d4(6)
    );
  rx_input_fifo_fifo_BU410 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3689,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1560_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1560
    );
  rx_input_fifo_fifo_N1560_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1560_FFX_SET
    );
  tx_fifocheck_fbbpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_11_FFY_RST
    );
  tx_fifocheck_fbbpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_11_FFY_RST,
      O => tx_fifocheck_fbbpl(10)
    );
  rx_input_fifo_fifo_BU281 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1528,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1541_FFY_RST,
      O => rx_input_fifo_fifo_N1542
    );
  rx_input_fifo_fifo_N1541_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1541_FFY_RST
    );
  tx_fifocheck_fbbpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_13_FFY_RST
    );
  tx_fifocheck_fbbpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_13_FFY_RST,
      O => tx_fifocheck_fbbpl(12)
    );
  tx_fifocheck_fbbpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_15_FFY_RST
    );
  tx_fifocheck_fbbpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_15_FFY_RST,
      O => tx_fifocheck_fbbpl(14)
    );
  rx_output_cs_FFd12_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd12_FFY_RST
    );
  rx_output_cs_FFd11_45 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd12,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd12_FFY_RST,
      O => rx_output_cs_FFd11
    );
  rx_output_cs_FFd14_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd14_FFY_RST
    );
  rx_output_cs_FFd13_46 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd14,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd14_FFY_RST,
      O => rx_output_cs_FFd13
    );
  rx_input_fifo_fifo_BU251 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3119,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1584_FFY_RST,
      O => rx_input_fifo_fifo_N1583
    );
  rx_input_fifo_fifo_N1584_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1584_FFY_RST
    );
  rx_output_cs_FFd16_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd16_FFY_RST
    );
  rx_output_cs_FFd15_47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd16,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd16_FFY_RST,
      O => rx_output_cs_FFd15
    );
  rx_output_cs_Out41 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_cs_FFd7,
      ADR2 => rx_output_cs_FFd12,
      ADR3 => rx_output_cs_FFd8,
      O => rx_output_cein
    );
  rx_output_n00331 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_cs_FFd12,
      ADR3 => RESET_IBUF,
      O => rx_output_ceinl_GROM
    );
  rx_output_ceinl_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_ceinl_CEMUXNOT
    );
  rx_output_ceinl_YUSED : X_BUF
    port map (
      I => rx_output_ceinl_GROM,
      O => rx_output_n0033
    );
  rx_output_cs_Out51 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_cs_FFd19,
      ADR2 => rx_output_cs_FFd10,
      ADR3 => VCC,
      O => rx_output_fifo_reset_FROM
    );
  rx_output_n00341 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => rx_output_cs_FFd10,
      O => rx_output_fifo_reset_GROM
    );
  rx_output_fifo_reset_XUSED : X_BUF
    port map (
      I => rx_output_fifo_reset_FROM,
      O => rx_output_fifo_reset
    );
  rx_output_fifo_reset_YUSED : X_BUF
    port map (
      I => rx_output_fifo_reset_GROM,
      O => rx_output_n0034
    );
  mac_control_Mmux_n0016_Result_6_97_SW1 : X_LUT4
    generic map(
      INIT => X"ABAF"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_phydo(6),
      ADR2 => mac_control_CHOICE2703,
      ADR3 => mac_control_n0060,
      O => mac_control_dout_6_FROM
    );
  mac_control_Mmux_n0016_Result_6_97 : X_LUT4
    generic map(
      INIT => X"4CEC"
    )
    port map (
      ADR0 => mac_control_sclkdeltall,
      ADR1 => mac_control_dout(5),
      ADR2 => mac_control_n0086,
      ADR3 => mac_control_N81447,
      O => mac_control_n0016(6)
    );
  mac_control_dout_6_XUSED : X_BUF
    port map (
      I => mac_control_dout_6_FROM,
      O => mac_control_N81447
    );
  tx_input_n00231 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => RESET_IBUF_1,
      ADR3 => tx_input_cs_FFd2,
      O => tx_input_n0023_FROM
    );
  tx_input_n00211 : X_LUT4
    generic map(
      INIT => X"00C8"
    )
    port map (
      ADR0 => tx_input_cs_FFd6,
      ADR1 => tx_input_den,
      ADR2 => tx_input_cs_FFd7,
      ADR3 => RESET_IBUF_1,
      O => tx_input_n0023_GROM
    );
  tx_input_n0023_XUSED : X_BUF
    port map (
      I => tx_input_n0023_FROM,
      O => tx_input_n0023
    );
  tx_input_n0023_YUSED : X_BUF
    port map (
      I => tx_input_n0023_GROM,
      O => tx_input_n0021
    );
  mac_control_Mmux_n0016_Result_7_93_SW1 : X_LUT4
    generic map(
      INIT => X"CDCF"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_addr(5),
      ADR2 => mac_control_CHOICE2474,
      ADR3 => mac_control_phydo(7),
      O => mac_control_dout_7_FROM
    );
  mac_control_Mmux_n0016_Result_7_93 : X_LUT4
    generic map(
      INIT => X"70F8"
    )
    port map (
      ADR0 => mac_control_n0086,
      ADR1 => mac_control_sclkdeltall,
      ADR2 => mac_control_dout(6),
      ADR3 => mac_control_N81451,
      O => mac_control_n0016(7)
    );
  mac_control_dout_7_XUSED : X_BUF
    port map (
      I => mac_control_dout_7_FROM,
      O => mac_control_N81451
    );
  mac_control_rxphyerr_cntl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_1_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_2_FFY_RST
    );
  mac_control_rxphyerr_cntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(2),
      CE => mac_control_rxphyerr_cntl_2_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_2_FFY_RST,
      O => mac_control_rxphyerr_cntl(2)
    );
  mac_control_rxphyerr_cntl_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_2_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_3_FFY_RST
    );
  mac_control_rxphyerr_cntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(3),
      CE => mac_control_rxphyerr_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_3_FFY_RST,
      O => mac_control_rxphyerr_cntl(3)
    );
  mac_control_rxphyerr_cntl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_3_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_5_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_7_FFY_RST
    );
  mac_control_rxphyerr_cntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(6),
      CE => mac_control_rxphyerr_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_7_FFY_RST,
      O => mac_control_rxphyerr_cntl(6)
    );
  mac_control_rxphyerr_cntl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_7_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_9_FFY_RST
    );
  mac_control_rxphyerr_cntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(8),
      CE => mac_control_rxphyerr_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_9_FFY_RST,
      O => mac_control_rxphyerr_cntl(8)
    );
  mac_control_rxphyerr_cntl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_9_CEMUXNOT
    );
  mac_control_n004014 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_159,
      ADR1 => mac_control_ledrx_cnt_158,
      ADR2 => mac_control_ledrx_cnt_157,
      ADR3 => mac_control_ledrx_cnt_156,
      O => mac_control_CHOICE1272_FROM
    );
  mac_control_n004023 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => mac_control_CHOICE1266,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE1269,
      ADR3 => mac_control_CHOICE1272,
      O => mac_control_CHOICE1272_GROM
    );
  mac_control_CHOICE1272_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1272_FROM,
      O => mac_control_CHOICE1272
    );
  mac_control_CHOICE1272_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1272_GROM,
      O => mac_control_n0040
    );
  rx_input_fifo_fifo_BU244 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3079,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1584_FFX_RST,
      O => rx_input_fifo_fifo_N1584
    );
  rx_input_fifo_fifo_N1584_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1584_FFX_RST
    );
  mac_control_n003223 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_130,
      ADR1 => mac_control_phyrstcnt_128,
      ADR2 => mac_control_phyrstcnt_111,
      ADR3 => mac_control_phyrstcnt_129,
      O => mac_control_CHOICE1387_FROM
    );
  mac_control_n003224 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE1384,
      ADR3 => mac_control_CHOICE1387,
      O => mac_control_CHOICE1387_GROM
    );
  mac_control_CHOICE1387_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1387_FROM,
      O => mac_control_CHOICE1387
    );
  mac_control_CHOICE1387_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1387_GROM,
      O => mac_control_CHOICE1388
    );
  mac_control_n0034161_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_117,
      ADR1 => mac_control_phyrstcnt_126,
      ADR2 => mac_control_phyrstcnt_125,
      ADR3 => mac_control_phyrstcnt_118,
      O => mac_control_N80971_FROM
    );
  mac_control_n003218 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_127,
      ADR1 => mac_control_phyrstcnt_125,
      ADR2 => mac_control_phyrstcnt_126,
      ADR3 => mac_control_phyrstcnt_124,
      O => mac_control_N80971_GROM
    );
  mac_control_N80971_XUSED : X_BUF
    port map (
      I => mac_control_N80971_FROM,
      O => mac_control_N80971
    );
  mac_control_N80971_YUSED : X_BUF
    port map (
      I => mac_control_N80971_GROM,
      O => mac_control_CHOICE1384
    );
  mac_control_n003444 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_139,
      ADR1 => mac_control_phyrstcnt_112,
      ADR2 => mac_control_phyrstcnt_138,
      ADR3 => mac_control_phyrstcnt_140,
      O => mac_control_CHOICE1333_FROM
    );
  mac_control_n003251 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_138,
      ADR1 => mac_control_phyrstcnt_136,
      ADR2 => mac_control_phyrstcnt_137,
      ADR3 => mac_control_phyrstcnt_135,
      O => mac_control_CHOICE1333_GROM
    );
  mac_control_CHOICE1333_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1333_FROM,
      O => mac_control_CHOICE1333
    );
  mac_control_CHOICE1333_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1333_GROM,
      O => mac_control_CHOICE1395
    );
  mac_control_n003421 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_137,
      ADR1 => mac_control_phyrstcnt_134,
      ADR2 => mac_control_phyrstcnt_136,
      ADR3 => mac_control_phyrstcnt_135,
      O => mac_control_CHOICE1325_FROM
    );
  mac_control_n003426 : X_LUT4
    generic map(
      INIT => X"0100"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_133,
      ADR1 => mac_control_phyrstcnt_132,
      ADR2 => mac_control_phyrstcnt_120,
      ADR3 => mac_control_CHOICE1325,
      O => mac_control_CHOICE1325_GROM
    );
  mac_control_CHOICE1325_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1325_FROM,
      O => mac_control_CHOICE1325
    );
  mac_control_CHOICE1325_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1325_GROM,
      O => mac_control_CHOICE1326
    );
  rx_input_fifo_fifo_BU204 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2687,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N6_FFY_RST,
      O => rx_input_fifo_fifo_N5
    );
  rx_input_fifo_fifo_N6_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N6_FFY_RST
    );
  mac_control_n003263 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_112,
      ADR1 => mac_control_phyrstcnt_139,
      ADR2 => mac_control_phyrstcnt_113,
      ADR3 => mac_control_phyrstcnt_140,
      O => mac_control_CHOICE1399_GROM
    );
  mac_control_CHOICE1399_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1399_GROM,
      O => mac_control_CHOICE1399
    );
  mac_control_n003268 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_114,
      ADR1 => mac_control_phyrstcnt_117,
      ADR2 => mac_control_phyrstcnt_116,
      ADR3 => mac_control_phyrstcnt_115,
      O => mac_control_CHOICE1402_GROM
    );
  mac_control_CHOICE1402_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1402_GROM,
      O => mac_control_CHOICE1402
    );
  mac_control_n003457 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_113,
      ADR1 => mac_control_phyrstcnt_114,
      ADR2 => mac_control_phyrstcnt_116,
      ADR3 => mac_control_phyrstcnt_115,
      O => mac_control_CHOICE1340_FROM
    );
  mac_control_n003458 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_CHOICE1333,
      ADR3 => mac_control_CHOICE1340,
      O => mac_control_CHOICE1340_GROM
    );
  mac_control_CHOICE1340_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1340_FROM,
      O => mac_control_CHOICE1340
    );
  mac_control_CHOICE1340_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1340_GROM,
      O => mac_control_CHOICE1341
    );
  mac_control_n00389 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_142,
      ADR1 => mac_control_ledtx_cnt_143,
      ADR2 => mac_control_ledtx_cnt_152,
      ADR3 => mac_control_ledtx_cnt_153,
      O => mac_control_CHOICE1280_FROM
    );
  mac_control_n003714 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_143,
      ADR1 => mac_control_ledtx_cnt_153,
      ADR2 => mac_control_ledtx_cnt_142,
      ADR3 => mac_control_ledtx_cnt_152,
      O => mac_control_CHOICE1280_GROM
    );
  mac_control_CHOICE1280_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1280_FROM,
      O => mac_control_CHOICE1280
    );
  mac_control_CHOICE1280_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1280_GROM,
      O => mac_control_CHOICE1308
    );
  rx_input_memio_addrchk_macaddrl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_7_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(6),
      CE => rx_input_memio_addrchk_macaddrl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_7_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(6)
    );
  rx_input_memio_addrchk_macaddrl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_7_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(7),
      CE => rx_input_memio_addrchk_macaddrl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_7_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(7)
    );
  rx_input_memio_addrchk_macaddrl_7_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_7_CEMUXNOT
    );
  rx_input_fifo_fifo_BU283 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1527,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1541_FFX_RST,
      O => rx_input_fifo_fifo_N1541
    );
  rx_input_fifo_fifo_N1541_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1541_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_9_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(8),
      CE => rx_input_memio_addrchk_macaddrl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_9_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(8)
    );
  rx_input_memio_addrchk_macaddrl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_9_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(9),
      CE => rx_input_memio_addrchk_macaddrl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_9_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(9)
    );
  rx_input_memio_addrchk_macaddrl_9_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_9_CEMUXNOT
    );
  memcontroller_n00061_1_48 : X_LUT4
    generic map(
      INIT => X"0500"
    )
    port map (
      ADR0 => memcontroller_clknum(0),
      ADR1 => VCC,
      ADR2 => RESET_IBUF,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_n00061_1_FROM
    );
  memcontroller_n00051_1_49 : X_LUT4
    generic map(
      INIT => X"0022"
    )
    port map (
      ADR0 => memcontroller_clknum(0),
      ADR1 => memcontroller_clknum(1),
      ADR2 => VCC,
      ADR3 => RESET_IBUF,
      O => memcontroller_n00061_1_GROM
    );
  memcontroller_n00061_1_XUSED : X_BUF
    port map (
      I => memcontroller_n00061_1_FROM,
      O => memcontroller_n00061_1
    );
  memcontroller_n00061_1_YUSED : X_BUF
    port map (
      I => memcontroller_n00061_1_GROM,
      O => memcontroller_n00051_1
    );
  mac_control_Mmux_n0016_Result_2_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cntl(2),
      ADR1 => mac_control_rxphyerr_cntl(2),
      ADR2 => mac_control_n0064,
      ADR3 => mac_control_n0065,
      O => mac_control_CHOICE2634_FROM
    );
  mac_control_Mmux_n0016_Result_10_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0065,
      ADR1 => mac_control_n0064,
      ADR2 => mac_control_rxfifowerr_cntl(10),
      ADR3 => mac_control_rxphyerr_cntl(10),
      O => mac_control_CHOICE2634_GROM
    );
  mac_control_CHOICE2634_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2634_FROM,
      O => mac_control_CHOICE2634
    );
  mac_control_CHOICE2634_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2634_GROM,
      O => mac_control_CHOICE2738
    );
  mac_control_Mmux_n0016_Result_9_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxf_cntl(9),
      ADR1 => mac_control_n0067,
      ADR2 => mac_control_rxcrcerr_cntl(9),
      ADR3 => mac_control_n0062,
      O => mac_control_CHOICE2508_FROM
    );
  mac_control_Mmux_n0016_Result_11_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cntl(11),
      ADR1 => mac_control_n0067,
      ADR2 => mac_control_n0062,
      ADR3 => mac_control_rxf_cntl(11),
      O => mac_control_CHOICE2508_GROM
    );
  mac_control_CHOICE2508_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2508_FROM,
      O => mac_control_CHOICE2508
    );
  mac_control_CHOICE2508_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2508_GROM,
      O => mac_control_CHOICE2483
    );
  mac_control_Mmux_n0016_Result_22_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cntl(22),
      ADR1 => mac_control_n0067,
      ADR2 => mac_control_rxf_cntl(22),
      ADR3 => mac_control_n0062,
      O => mac_control_CHOICE2105_FROM
    );
  mac_control_Mmux_n0016_Result_20_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cntl(20),
      ADR1 => mac_control_n0067,
      ADR2 => mac_control_rxf_cntl(20),
      ADR3 => mac_control_n0062,
      O => mac_control_CHOICE2105_GROM
    );
  mac_control_CHOICE2105_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2105_FROM,
      O => mac_control_CHOICE2105
    );
  mac_control_CHOICE2105_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2105_GROM,
      O => mac_control_CHOICE2128
    );
  mac_control_Mmux_n0016_Result_28_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxf_cntl(28),
      ADR1 => mac_control_n0062,
      ADR2 => mac_control_rxcrcerr_cntl(28),
      ADR3 => mac_control_n0067,
      O => mac_control_CHOICE2243_FROM
    );
  mac_control_Mmux_n0016_Result_12_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0067,
      ADR1 => mac_control_rxcrcerr_cntl(12),
      ADR2 => mac_control_rxf_cntl(12),
      ADR3 => mac_control_n0062,
      O => mac_control_CHOICE2243_GROM
    );
  mac_control_CHOICE2243_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2243_FROM,
      O => mac_control_CHOICE2243
    );
  mac_control_CHOICE2243_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2243_GROM,
      O => mac_control_CHOICE2533
    );
  mac_control_Mmux_n0016_Result_15_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cntl(15),
      ADR1 => mac_control_rxf_cntl(15),
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_n0062,
      O => mac_control_CHOICE2583_FROM
    );
  mac_control_Mmux_n0016_Result_13_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0067,
      ADR1 => mac_control_n0062,
      ADR2 => mac_control_rxcrcerr_cntl(13),
      ADR3 => mac_control_rxf_cntl(13),
      O => mac_control_CHOICE2583_GROM
    );
  mac_control_CHOICE2583_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2583_FROM,
      O => mac_control_CHOICE2583
    );
  mac_control_CHOICE2583_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2583_GROM,
      O => mac_control_CHOICE2558
    );
  mac_control_Mmux_n0016_Result_8_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cntl(8),
      ADR1 => mac_control_rxfifowerr_cntl(8),
      ADR2 => mac_control_n0064,
      ADR3 => mac_control_n0065,
      O => mac_control_CHOICE2712_FROM
    );
  mac_control_Mmux_n0016_Result_21_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cntl(21),
      ADR1 => mac_control_n0065,
      ADR2 => mac_control_rxphyerr_cntl(21),
      ADR3 => mac_control_n0064,
      O => mac_control_CHOICE2712_GROM
    );
  mac_control_CHOICE2712_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2712_FROM,
      O => mac_control_CHOICE2712
    );
  mac_control_CHOICE2712_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2712_GROM,
      O => mac_control_CHOICE2360
    );
  mac_control_Mmux_n0016_Result_26_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0062,
      ADR1 => mac_control_rxcrcerr_cntl(26),
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_rxf_cntl(26),
      O => mac_control_CHOICE2174_FROM
    );
  mac_control_Mmux_n0016_Result_30_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0062,
      ADR1 => mac_control_rxcrcerr_cntl(30),
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_rxf_cntl(30),
      O => mac_control_CHOICE2174_GROM
    );
  mac_control_CHOICE2174_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2174_FROM,
      O => mac_control_CHOICE2174
    );
  mac_control_CHOICE2174_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2174_GROM,
      O => mac_control_CHOICE2289
    );
  mac_control_Mmux_n0016_Result_24_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_rxphyerr_cntl(24),
      ADR2 => mac_control_rxfifowerr_cntl(24),
      ADR3 => mac_control_n0065,
      O => mac_control_CHOICE2384_FROM
    );
  mac_control_Mmux_n0016_Result_14_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cntl(14),
      ADR1 => mac_control_n0065,
      ADR2 => mac_control_n0064,
      ADR3 => mac_control_rxphyerr_cntl(14),
      O => mac_control_CHOICE2384_GROM
    );
  mac_control_CHOICE2384_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2384_FROM,
      O => mac_control_CHOICE2384
    );
  mac_control_CHOICE2384_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2384_GROM,
      O => mac_control_CHOICE2764
    );
  mac_control_Mmux_n0016_Result_24_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0066,
      ADR1 => mac_control_n0059,
      ADR2 => mac_control_rxoferr_cntl(24),
      ADR3 => mac_control_phydi(24),
      O => mac_control_CHOICE2387_FROM
    );
  mac_control_Mmux_n0016_Result_0_10 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxoferr_cntl(0),
      ADR1 => mac_control_phydi(0),
      ADR2 => mac_control_n0059,
      ADR3 => mac_control_n0066,
      O => mac_control_CHOICE2387_GROM
    );
  mac_control_CHOICE2387_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2387_FROM,
      O => mac_control_CHOICE2387
    );
  mac_control_CHOICE2387_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2387_GROM,
      O => mac_control_CHOICE1895
    );
  mac_control_Mmux_n0016_Result_19_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cntl(19),
      ADR1 => mac_control_rxf_cntl(19),
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_n0062,
      O => mac_control_CHOICE2082_FROM
    );
  mac_control_Mmux_n0016_Result_23_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0067,
      ADR1 => mac_control_n0062,
      ADR2 => mac_control_rxcrcerr_cntl(23),
      ADR3 => mac_control_rxf_cntl(23),
      O => mac_control_CHOICE2082_GROM
    );
  mac_control_CHOICE2082_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2082_FROM,
      O => mac_control_CHOICE2082
    );
  mac_control_CHOICE2082_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2082_GROM,
      O => mac_control_CHOICE2151
    );
  mac_control_Mmux_n0016_Result_6_30 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cntl(6),
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_n00851_1,
      ADR3 => mac_control_phyaddr(6),
      O => mac_control_CHOICE2698_FROM
    );
  mac_control_Mmux_n0016_Result_0_30 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_phyaddr(0),
      ADR2 => mac_control_txfifowerr_cntl(0),
      ADR3 => mac_control_n0063,
      O => mac_control_CHOICE2698_GROM
    );
  mac_control_CHOICE2698_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2698_FROM,
      O => mac_control_CHOICE2698
    );
  mac_control_CHOICE2698_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2698_GROM,
      O => mac_control_CHOICE1904
    );
  mac_control_Mmux_n0016_Result_0_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0061,
      ADR1 => mac_control_rxf_cntl(0),
      ADR2 => mac_control_n0062,
      ADR3 => mac_control_txf_cntl(0),
      O => mac_control_CHOICE1899_FROM
    );
  mac_control_Mmux_n0016_Result_0_48_SW0 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_n0056,
      ADR1 => mac_control_rxcrcerr_cntl(0),
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_CHOICE1899,
      O => mac_control_CHOICE1899_GROM
    );
  mac_control_CHOICE1899_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1899_FROM,
      O => mac_control_CHOICE1899
    );
  mac_control_CHOICE1899_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1899_GROM,
      O => mac_control_N81050
    );
  mac_control_Mmux_n0016_Result_5_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cntl(5),
      ADR1 => mac_control_n0065,
      ADR2 => mac_control_n0064,
      ADR3 => mac_control_rxfifowerr_cntl(5),
      O => mac_control_CHOICE2660_FROM
    );
  mac_control_Mmux_n0016_Result_16_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_rxphyerr_cntl(16),
      ADR2 => mac_control_rxfifowerr_cntl(16),
      ADR3 => mac_control_n0065,
      O => mac_control_CHOICE2660_GROM
    );
  mac_control_CHOICE2660_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2660_FROM,
      O => mac_control_CHOICE2660
    );
  mac_control_CHOICE2660_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2660_GROM,
      O => mac_control_CHOICE2312
    );
  mac_control_Mmux_n0016_Result_2_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0066,
      ADR1 => mac_control_rxoferr_cntl(2),
      ADR2 => mac_control_n0059,
      ADR3 => mac_control_phydi(2),
      O => mac_control_CHOICE2637_FROM
    );
  mac_control_Mmux_n0016_Result_1_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0066,
      ADR1 => mac_control_rxoferr_cntl(1),
      ADR2 => mac_control_n0059,
      ADR3 => mac_control_phydi(1),
      O => mac_control_CHOICE2637_GROM
    );
  mac_control_CHOICE2637_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2637_FROM,
      O => mac_control_CHOICE2637
    );
  mac_control_CHOICE2637_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2637_GROM,
      O => mac_control_CHOICE2611
    );
  mac_control_Mmux_n0016_Result_31_22 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cntl(31),
      ADR1 => mac_control_rxfifowerr_cntl(31),
      ADR2 => mac_control_n0065,
      ADR3 => mac_control_n0064,
      O => mac_control_CHOICE2043_FROM
    );
  mac_control_Mmux_n0016_Result_17_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cntl(17),
      ADR1 => mac_control_n0064,
      ADR2 => mac_control_n0065,
      ADR3 => mac_control_rxfifowerr_cntl(17),
      O => mac_control_CHOICE2043_GROM
    );
  mac_control_CHOICE2043_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2043_FROM,
      O => mac_control_CHOICE2043
    );
  mac_control_CHOICE2043_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2043_GROM,
      O => mac_control_CHOICE2336
    );
  mac_control_Mmux_n0016_Result_4_5 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0067,
      ADR1 => mac_control_rxcrcerr_cntl(4),
      ADR2 => mac_control_n0062,
      ADR3 => mac_control_rxf_cntl(4),
      O => mac_control_CHOICE2408_FROM
    );
  mac_control_Mmux_n0016_Result_25_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0062,
      ADR1 => mac_control_n0067,
      ADR2 => mac_control_rxf_cntl(25),
      ADR3 => mac_control_rxcrcerr_cntl(25),
      O => mac_control_CHOICE2408_GROM
    );
  mac_control_CHOICE2408_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2408_FROM,
      O => mac_control_CHOICE2408
    );
  mac_control_CHOICE2408_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2408_GROM,
      O => mac_control_CHOICE2197
    );
  mac_control_Mmux_n0016_Result_1_22 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxf_cntl(1),
      ADR1 => mac_control_n0061,
      ADR2 => mac_control_n0062,
      ADR3 => mac_control_txf_cntl(1),
      O => mac_control_CHOICE2615_FROM
    );
  mac_control_Mmux_n0016_Result_1_48_SW0 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_n0056,
      ADR1 => mac_control_rxcrcerr_cntl(1),
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_CHOICE2615,
      O => mac_control_CHOICE2615_GROM
    );
  mac_control_CHOICE2615_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2615_FROM,
      O => mac_control_CHOICE2615
    );
  mac_control_CHOICE2615_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2615_GROM,
      O => mac_control_N81034
    );
  mac_control_Mmux_n0016_Result_0_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_N81050,
      ADR1 => mac_control_CHOICE1892,
      ADR2 => mac_control_CHOICE1904,
      ADR3 => mac_control_CHOICE1895,
      O => mac_control_dout_0_FROM
    );
  mac_control_Mmux_n0016_Result_0_82 : X_LUT4
    generic map(
      INIT => X"4404"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_n0044,
      ADR2 => mac_control_N81030,
      ADR3 => mac_control_CHOICE1907,
      O => mac_control_n0016(0)
    );
  mac_control_dout_0_XUSED : X_BUF
    port map (
      I => mac_control_dout_0_FROM,
      O => mac_control_CHOICE1907
    );
  mac_control_Mmux_n0016_Result_27_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0062,
      ADR1 => mac_control_rxcrcerr_cntl(27),
      ADR2 => mac_control_rxf_cntl(27),
      ADR3 => mac_control_n0067,
      O => mac_control_CHOICE2220_FROM
    );
  mac_control_Mmux_n0016_Result_18_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0062,
      ADR1 => mac_control_rxcrcerr_cntl(18),
      ADR2 => mac_control_rxf_cntl(18),
      ADR3 => mac_control_n0067,
      O => mac_control_CHOICE2220_GROM
    );
  mac_control_CHOICE2220_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2220_FROM,
      O => mac_control_CHOICE2220
    );
  mac_control_CHOICE2220_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2220_GROM,
      O => mac_control_CHOICE2059
    );
  rx_input_fifo_fifo_BU404 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3686,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1562_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1563
    );
  rx_input_fifo_fifo_N1562_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1562_FFY_SET
    );
  mac_control_Mmux_n0016_Result_2_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cntl(2),
      ADR1 => mac_control_n0061,
      ADR2 => mac_control_rxf_cntl(2),
      ADR3 => mac_control_n0062,
      O => mac_control_CHOICE2641_FROM
    );
  mac_control_Mmux_n0016_Result_2_48_SW0 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_n0056,
      ADR1 => mac_control_rxcrcerr_cntl(2),
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_CHOICE2641,
      O => mac_control_CHOICE2641_GROM
    );
  mac_control_CHOICE2641_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2641_FROM,
      O => mac_control_CHOICE2641
    );
  mac_control_CHOICE2641_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2641_GROM,
      O => mac_control_N81062
    );
  mac_control_Mmux_n0016_Result_21_30 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0063,
      ADR1 => mac_control_txfifowerr_cntl(21),
      ADR2 => mac_control_phyaddr(21),
      ADR3 => mac_control_n00851_1,
      O => mac_control_CHOICE2372_FROM
    );
  mac_control_Mmux_n0016_Result_2_30 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_phyaddr(2),
      ADR2 => mac_control_n0063,
      ADR3 => mac_control_txfifowerr_cntl(2),
      O => mac_control_CHOICE2372_GROM
    );
  mac_control_CHOICE2372_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2372_FROM,
      O => mac_control_CHOICE2372
    );
  mac_control_CHOICE2372_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2372_GROM,
      O => mac_control_CHOICE2646
    );
  mac_control_Mmux_n0016_Result_1_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2620,
      ADR1 => mac_control_N81034,
      ADR2 => mac_control_CHOICE2611,
      ADR3 => mac_control_CHOICE2608,
      O => mac_control_CHOICE2623_FROM
    );
  mac_control_Mmux_n0016_Result_1_60 : X_LUT4
    generic map(
      INIT => X"FFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0057,
      ADR2 => mac_control_phystat(1),
      ADR3 => mac_control_CHOICE2623,
      O => mac_control_CHOICE2623_GROM
    );
  mac_control_CHOICE2623_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2623_FROM,
      O => mac_control_CHOICE2623
    );
  mac_control_CHOICE2623_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2623_GROM,
      O => mac_control_CHOICE2625
    );
  mac_control_Mmux_n0016_Result_22_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cntl(22),
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_n0064,
      ADR3 => mac_control_txfifowerr_cntl(22),
      O => mac_control_CHOICE2108_FROM
    );
  mac_control_Mmux_n0016_Result_3_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0063,
      ADR1 => mac_control_txfifowerr_cntl(3),
      ADR2 => mac_control_rxfifowerr_cntl(3),
      ADR3 => mac_control_n0064,
      O => mac_control_CHOICE2108_GROM
    );
  mac_control_CHOICE2108_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2108_FROM,
      O => mac_control_CHOICE2108
    );
  mac_control_CHOICE2108_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2108_GROM,
      O => mac_control_CHOICE2436
    );
  mac_control_Mmux_n0016_Result_3_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0067,
      ADR1 => mac_control_rxf_cntl(3),
      ADR2 => mac_control_n0062,
      ADR3 => mac_control_rxcrcerr_cntl(3),
      O => mac_control_CHOICE2433_FROM
    );
  mac_control_Mmux_n0016_Result_29_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cntl(29),
      ADR1 => mac_control_rxf_cntl(29),
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_n0062,
      O => mac_control_CHOICE2433_GROM
    );
  mac_control_CHOICE2433_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2433_FROM,
      O => mac_control_CHOICE2433
    );
  mac_control_CHOICE2433_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2433_GROM,
      O => mac_control_CHOICE2266
    );
  mac_control_Mmux_n0016_Result_30_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phyaddr(30),
      ADR1 => mac_control_n00851_1,
      ADR2 => mac_control_n0065,
      ADR3 => mac_control_rxphyerr_cntl(30),
      O => mac_control_CHOICE2296_FROM
    );
  mac_control_Mmux_n0016_Result_3_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0065,
      ADR1 => mac_control_n00851_1,
      ADR2 => mac_control_phyaddr(3),
      ADR3 => mac_control_rxphyerr_cntl(3),
      O => mac_control_CHOICE2296_GROM
    );
  mac_control_CHOICE2296_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2296_FROM,
      O => mac_control_CHOICE2296
    );
  mac_control_CHOICE2296_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2296_GROM,
      O => mac_control_CHOICE2440
    );
  mac_control_Mmux_n0016_Result_2_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2634,
      ADR1 => mac_control_CHOICE2646,
      ADR2 => mac_control_CHOICE2637,
      ADR3 => mac_control_N81062,
      O => mac_control_CHOICE2649_FROM
    );
  mac_control_Mmux_n0016_Result_2_60 : X_LUT4
    generic map(
      INIT => X"FFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phystat(2),
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_CHOICE2649,
      O => mac_control_CHOICE2649_GROM
    );
  mac_control_CHOICE2649_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2649_FROM,
      O => mac_control_CHOICE2649
    );
  mac_control_CHOICE2649_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2649_GROM,
      O => mac_control_CHOICE2651
    );
  rx_input_fifo_fifo_BU348 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1527,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1555_FFX_RST,
      O => rx_input_fifo_fifo_N1555
    );
  rx_input_fifo_fifo_N1555_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1555_FFX_RST
    );
  mac_control_Mmux_n0016_Result_28_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_rxfifowerr_cntl(28),
      ADR2 => mac_control_txfifowerr_cntl(28),
      ADR3 => mac_control_n0063,
      O => mac_control_CHOICE2246_FROM
    );
  mac_control_Mmux_n0016_Result_4_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_rxfifowerr_cntl(4),
      ADR2 => mac_control_n0063,
      ADR3 => mac_control_txfifowerr_cntl(4),
      O => mac_control_CHOICE2246_GROM
    );
  mac_control_CHOICE2246_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2246_FROM,
      O => mac_control_CHOICE2246
    );
  mac_control_CHOICE2246_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2246_GROM,
      O => mac_control_CHOICE2411
    );
  mac_control_Mmux_n0016_Result_3_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0066,
      ADR1 => mac_control_rxoferr_cntl(3),
      ADR2 => mac_control_n0061,
      ADR3 => mac_control_txf_cntl(3),
      O => mac_control_CHOICE2444_FROM
    );
  mac_control_Mmux_n0016_Result_3_45_SW0 : X_LUT4
    generic map(
      INIT => X"FF88"
    )
    port map (
      ADR0 => mac_control_phydi(3),
      ADR1 => mac_control_n0059,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2444,
      O => mac_control_CHOICE2444_GROM
    );
  mac_control_CHOICE2444_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2444_FROM,
      O => mac_control_CHOICE2444
    );
  mac_control_CHOICE2444_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2444_GROM,
      O => mac_control_N81106
    );
  mac_control_Mmux_n0016_Result_3_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2436,
      ADR1 => mac_control_CHOICE2440,
      ADR2 => mac_control_N81106,
      ADR3 => mac_control_CHOICE2433,
      O => mac_control_CHOICE2447_FROM
    );
  mac_control_Mmux_n0016_Result_3_56 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_phystat(3),
      ADR1 => VCC,
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_CHOICE2447,
      O => mac_control_CHOICE2447_GROM
    );
  mac_control_CHOICE2447_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2447_FROM,
      O => mac_control_CHOICE2447
    );
  mac_control_CHOICE2447_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2447_GROM,
      O => mac_control_CHOICE2449
    );
  mac_control_Mmux_n0016_Result_8_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxoferr_cntl(8),
      ADR1 => mac_control_phydi(8),
      ADR2 => mac_control_n0066,
      ADR3 => mac_control_n0059,
      O => mac_control_CHOICE2715_FROM
    );
  mac_control_Mmux_n0016_Result_5_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0059,
      ADR1 => mac_control_phydi(5),
      ADR2 => mac_control_rxoferr_cntl(5),
      ADR3 => mac_control_n0066,
      O => mac_control_CHOICE2715_GROM
    );
  mac_control_CHOICE2715_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2715_FROM,
      O => mac_control_CHOICE2715
    );
  mac_control_CHOICE2715_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2715_GROM,
      O => mac_control_CHOICE2663
    );
  mac_control_Mmux_n0016_Result_4_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0066,
      ADR1 => mac_control_rxoferr_cntl(4),
      ADR2 => mac_control_txf_cntl(4),
      ADR3 => mac_control_n0061,
      O => mac_control_CHOICE2419_FROM
    );
  mac_control_Mmux_n0016_Result_4_45_SW0 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_phydi(4),
      ADR1 => VCC,
      ADR2 => mac_control_n0059,
      ADR3 => mac_control_CHOICE2419,
      O => mac_control_CHOICE2419_GROM
    );
  mac_control_CHOICE2419_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2419_FROM,
      O => mac_control_CHOICE2419
    );
  mac_control_CHOICE2419_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2419_GROM,
      O => mac_control_N81122
    );
  mac_control_Mmux_n0016_Result_4_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_N81122,
      ADR1 => mac_control_CHOICE2408,
      ADR2 => mac_control_CHOICE2415,
      ADR3 => mac_control_CHOICE2411,
      O => mac_control_CHOICE2422_FROM
    );
  mac_control_Mmux_n0016_Result_4_56 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_phystat(4),
      ADR1 => VCC,
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_CHOICE2422,
      O => mac_control_CHOICE2422_GROM
    );
  mac_control_CHOICE2422_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2422_FROM,
      O => mac_control_CHOICE2422
    );
  mac_control_CHOICE2422_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2422_GROM,
      O => mac_control_CHOICE2424
    );
  mac_control_Mmux_n0016_Result_5_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxf_cntl(5),
      ADR1 => mac_control_txf_cntl(5),
      ADR2 => mac_control_n0061,
      ADR3 => mac_control_n0062,
      O => mac_control_CHOICE2667_FROM
    );
  mac_control_Mmux_n0016_Result_5_48_SW0 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_n0056,
      ADR1 => mac_control_n0067,
      ADR2 => mac_control_rxcrcerr_cntl(5),
      ADR3 => mac_control_CHOICE2667,
      O => mac_control_CHOICE2667_GROM
    );
  mac_control_CHOICE2667_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2667_FROM,
      O => mac_control_CHOICE2667
    );
  mac_control_CHOICE2667_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2667_GROM,
      O => mac_control_N81054
    );
  mac_control_Mmux_n0016_Result_16_30 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phyaddr(16),
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_txfifowerr_cntl(16),
      ADR3 => mac_control_n00851_1,
      O => mac_control_CHOICE2324_FROM
    );
  mac_control_Mmux_n0016_Result_5_30 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_phyaddr(5),
      ADR3 => mac_control_txfifowerr_cntl(5),
      O => mac_control_CHOICE2324_GROM
    );
  mac_control_CHOICE2324_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2324_FROM,
      O => mac_control_CHOICE2324
    );
  mac_control_CHOICE2324_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2324_GROM,
      O => mac_control_CHOICE2672
    );
  mac_control_Mmux_n0016_Result_10_10 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0059,
      ADR1 => mac_control_n0066,
      ADR2 => mac_control_rxoferr_cntl(10),
      ADR3 => mac_control_phydi(10),
      O => mac_control_CHOICE2741_FROM
    );
  mac_control_Mmux_n0016_Result_6_10 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0059,
      ADR1 => mac_control_n0066,
      ADR2 => mac_control_rxoferr_cntl(6),
      ADR3 => mac_control_phydi(6),
      O => mac_control_CHOICE2741_GROM
    );
  mac_control_CHOICE2741_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2741_FROM,
      O => mac_control_CHOICE2741
    );
  mac_control_CHOICE2741_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2741_GROM,
      O => mac_control_CHOICE2689
    );
  mac_control_Mmux_n0016_Result_6_22 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0062,
      ADR1 => mac_control_n0061,
      ADR2 => mac_control_rxf_cntl(6),
      ADR3 => mac_control_txf_cntl(6),
      O => mac_control_CHOICE2693_FROM
    );
  mac_control_Mmux_n0016_Result_6_48_SW0 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => mac_control_n0067,
      ADR1 => mac_control_n0056,
      ADR2 => mac_control_rxcrcerr_cntl(6),
      ADR3 => mac_control_CHOICE2693,
      O => mac_control_CHOICE2693_GROM
    );
  mac_control_CHOICE2693_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2693_FROM,
      O => mac_control_CHOICE2693
    );
  mac_control_CHOICE2693_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2693_GROM,
      O => mac_control_N81078
    );
  mac_control_Mmux_n0016_Result_5_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2663,
      ADR1 => mac_control_CHOICE2672,
      ADR2 => mac_control_CHOICE2660,
      ADR3 => mac_control_N81054,
      O => mac_control_CHOICE2675_FROM
    );
  mac_control_Mmux_n0016_Result_5_60 : X_LUT4
    generic map(
      INIT => X"FF88"
    )
    port map (
      ADR0 => mac_control_n0057,
      ADR1 => mac_control_phystat(5),
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2675,
      O => mac_control_CHOICE2675_GROM
    );
  mac_control_CHOICE2675_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2675_FROM,
      O => mac_control_CHOICE2675
    );
  mac_control_CHOICE2675_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2675_GROM,
      O => mac_control_CHOICE2677
    );
  rx_input_memio_crccomb_Mxor_CO_7_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(24),
      ADR1 => rx_input_memio_crcl(27),
      ADR2 => rx_input_memio_datal(4),
      ADR3 => rx_input_memio_datal(7),
      O => rx_input_memio_crccomb_Mxor_CO_7_Xo_1_FROM
    );
  rx_input_memio_crccomb_Mxor_n0004_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcl(27),
      ADR3 => rx_input_memio_datal(4),
      O => rx_input_memio_crccomb_Mxor_CO_7_Xo_1_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_7_Xo_1_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_7_Xo_1_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_7_Xo(1)
    );
  rx_input_memio_crccomb_Mxor_CO_7_Xo_1_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_7_Xo_1_GROM,
      O => rx_input_memio_crccomb_n0124(1)
    );
  rx_input_memio_crccomb_Mxor_CO_9_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_datal(6),
      ADR1 => rx_input_memio_crcl(28),
      ADR2 => rx_input_memio_datal(3),
      ADR3 => rx_input_memio_crcl(25),
      O => rx_input_memio_crccomb_Mxor_CO_9_Xo_0_FROM
    );
  rx_input_memio_crccomb_Mxor_n0012_Result1 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_input_memio_datal(6),
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcl(25),
      ADR3 => VCC,
      O => rx_input_memio_crccomb_Mxor_CO_9_Xo_0_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_9_Xo_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_9_Xo_0_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_9_Xo(0)
    );
  rx_input_memio_crccomb_Mxor_CO_9_Xo_0_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_9_Xo_0_GROM,
      O => rx_input_memio_crccomb_n0122(0)
    );
  mac_control_Mmux_n0016_Result_30_10 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cntl(30),
      ADR1 => mac_control_txfifowerr_cntl(30),
      ADR2 => mac_control_n0063,
      ADR3 => mac_control_n0064,
      O => mac_control_CHOICE2292_FROM
    );
  mac_control_Mmux_n0016_Result_7_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0063,
      ADR1 => mac_control_rxfifowerr_cntl(7),
      ADR2 => mac_control_txfifowerr_cntl(7),
      ADR3 => mac_control_n0064,
      O => mac_control_CHOICE2292_GROM
    );
  mac_control_CHOICE2292_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2292_FROM,
      O => mac_control_CHOICE2292
    );
  mac_control_CHOICE2292_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2292_GROM,
      O => mac_control_CHOICE2461
    );
  mac_control_PHY_status_MII_Interface_dreg_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_6_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(4),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_6_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(5)
    );
  mac_control_n003814 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_146,
      ADR1 => mac_control_ledtx_cnt_147,
      ADR2 => mac_control_ledtx_cnt_144,
      ADR3 => mac_control_ledtx_cnt_145,
      O => mac_control_CHOICE1283_FROM
    );
  mac_control_n003823 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_CHOICE1280,
      ADR2 => mac_control_CHOICE1277,
      ADR3 => mac_control_CHOICE1283,
      O => mac_control_CHOICE1283_GROM
    );
  mac_control_CHOICE1283_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1283_FROM,
      O => mac_control_CHOICE1283
    );
  mac_control_CHOICE1283_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1283_GROM,
      O => mac_control_n0038
    );
  mac_control_n003735 : X_LUT4
    generic map(
      INIT => X"F8F0"
    )
    port map (
      ADR0 => mac_control_CHOICE1302,
      ADR1 => mac_control_CHOICE1305,
      ADR2 => mac_control_ledtx_rst,
      ADR3 => mac_control_CHOICE1308,
      O => mac_control_CHOICE1311_FROM
    );
  mac_control_n003746 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE1311,
      O => mac_control_CHOICE1311_GROM
    );
  mac_control_CHOICE1311_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1311_FROM,
      O => mac_control_CHOICE1311
    );
  mac_control_CHOICE1311_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1311_GROM,
      O => mac_control_n0037
    );
  mac_control_PHY_status_MII_Interface_dreg_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_10_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(8),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_10_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(9)
    );
  mac_control_n00409 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_164,
      ADR1 => mac_control_ledrx_cnt_155,
      ADR2 => mac_control_ledrx_cnt_165,
      ADR3 => mac_control_ledrx_cnt_154,
      O => mac_control_CHOICE1269_FROM
    );
  mac_control_n003914 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_154,
      ADR1 => mac_control_ledrx_cnt_164,
      ADR2 => mac_control_ledrx_cnt_155,
      ADR3 => mac_control_ledrx_cnt_165,
      O => mac_control_CHOICE1269_GROM
    );
  mac_control_CHOICE1269_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1269_FROM,
      O => mac_control_CHOICE1269
    );
  mac_control_CHOICE1269_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1269_GROM,
      O => mac_control_CHOICE1294
    );
  mac_control_n003935 : X_LUT4
    generic map(
      INIT => X"ECCC"
    )
    port map (
      ADR0 => mac_control_CHOICE1288,
      ADR1 => mac_control_ledrx_rst,
      ADR2 => mac_control_CHOICE1291,
      ADR3 => mac_control_CHOICE1294,
      O => mac_control_CHOICE1297_FROM
    );
  mac_control_n003946 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE1297,
      O => mac_control_CHOICE1297_GROM
    );
  mac_control_CHOICE1297_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1297_FROM,
      O => mac_control_CHOICE1297
    );
  mac_control_CHOICE1297_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1297_GROM,
      O => mac_control_n0039
    );
  mac_control_Mmux_n0016_Result_8_97_SW1 : X_LUT4
    generic map(
      INIT => X"F1F5"
    )
    port map (
      ADR0 => mac_control_CHOICE2729,
      ADR1 => mac_control_n0060,
      ADR2 => mac_control_addr(5),
      ADR3 => mac_control_phydo(8),
      O => mac_control_dout_8_FROM
    );
  mac_control_Mmux_n0016_Result_8_97 : X_LUT4
    generic map(
      INIT => X"70F8"
    )
    port map (
      ADR0 => mac_control_n0086,
      ADR1 => mac_control_sclkdeltall,
      ADR2 => mac_control_dout(7),
      ADR3 => mac_control_N81455,
      O => mac_control_n0016(8)
    );
  mac_control_dout_8_XUSED : X_BUF
    port map (
      I => mac_control_dout_8_FROM,
      O => mac_control_N81455
    );
  tx_input_dh_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_3_FFY_RST
    );
  tx_input_dh_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(2),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_3_FFY_RST,
      O => tx_input_dh(2)
    );
  tx_input_dh_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_5_FFY_RST
    );
  tx_input_dh_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(4),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_5_FFY_RST,
      O => tx_input_dh(4)
    );
  rx_input_memio_crccomb_Mxor_CO_14_Xo_3_1_SW0 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_datal(3),
      ADR1 => rx_input_memio_datal(5),
      ADR2 => rx_input_memio_crcl(6),
      ADR3 => rx_input_memio_crcl(28),
      O => rx_input_memio_crccomb_N81261_FROM
    );
  rx_input_memio_crccomb_Mxor_n0003_Result1 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_datal(5),
      ADR2 => VCC,
      ADR3 => rx_input_memio_crcl(26),
      O => rx_input_memio_crccomb_N81261_GROM
    );
  rx_input_memio_crccomb_N81261_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_N81261_FROM,
      O => rx_input_memio_crccomb_N81261
    );
  rx_input_memio_crccomb_N81261_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_N81261_GROM,
      O => rx_input_memio_crccomb_n0118(1)
    );
  rx_input_memio_crccomb_Mxor_n0011_Result1 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_datal(0),
      ADR2 => rx_input_memio_crcl(31),
      ADR3 => VCC,
      O => rx_input_memio_crccomb_n0124_0_GROM
    );
  rx_input_memio_crccomb_n0124_0_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_n0124_0_GROM,
      O => rx_input_memio_crccomb_n0124(0)
    );
  tx_input_dh_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_9_FFY_RST
    );
  tx_input_dh_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(8),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_9_FFY_RST,
      O => tx_input_dh(8)
    );
  txbp_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_1_FFY_RST
    );
  tx_input_bp_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_16,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_1_FFY_RST,
      O => txbp(0)
    );
  tx_input_dl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_3_FFY_RST
    );
  tx_input_dl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(2),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_3_FFY_RST,
      O => tx_input_dl(2)
    );
  tx_input_dl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_5_FFY_RST
    );
  tx_input_dl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(4),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_5_FFY_RST,
      O => tx_input_dl(4)
    );
  rx_input_fifo_fifo_BU198 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2686,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N6_FFX_RST,
      O => rx_input_fifo_fifo_N6
    );
  rx_input_fifo_fifo_N6_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N6_FFX_RST
    );
  tx_input_dl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_7_FFY_RST
    );
  tx_input_dl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(6),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_7_FFY_RST,
      O => tx_input_dl(6)
    );
  tx_input_dl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_9_FFY_RST
    );
  tx_input_dl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(8),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_9_FFY_RST,
      O => tx_input_dl(8)
    );
  MDC_OBUF_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MDC_OBUF_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_mdcint : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_37,
      CE => MDC_OBUF_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MDC_OBUF_FFY_RST,
      O => MDC_OBUF
    );
  MDC_OBUF_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => MDC_OBUF_CEMUXNOT
    );
  mac_control_dout_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_9_FFY_RST
    );
  mac_control_dout_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(9),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_9_FFY_RST,
      O => mac_control_dout(9)
    );
  mac_control_Mmux_n0016_Result_9_93_SW1 : X_LUT4
    generic map(
      INIT => X"ABAF"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_n0060,
      ADR2 => mac_control_CHOICE2524,
      ADR3 => mac_control_phydo(9),
      O => mac_control_dout_9_FROM
    );
  mac_control_Mmux_n0016_Result_9_93 : X_LUT4
    generic map(
      INIT => X"2AEA"
    )
    port map (
      ADR0 => mac_control_dout(8),
      ADR1 => mac_control_sclkdeltall,
      ADR2 => mac_control_n0086,
      ADR3 => mac_control_N81459,
      O => mac_control_n0016(9)
    );
  mac_control_dout_9_XUSED : X_BUF
    port map (
      I => mac_control_dout_9_FROM,
      O => mac_control_N81459
    );
  mac_control_lmacaddr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_3_FFY_RST
    );
  mac_control_lmacaddr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_3_FFY_RST,
      O => mac_control_lmacaddr(2)
    );
  mac_control_lmacaddr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_5_FFY_RST
    );
  mac_control_lmacaddr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_5_FFY_RST,
      O => mac_control_lmacaddr(4)
    );
  mac_control_lmacaddr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_7_FFY_RST
    );
  mac_control_lmacaddr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_7_FFY_RST,
      O => mac_control_lmacaddr(6)
    );
  mac_control_lmacaddr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_9_FFY_RST
    );
  mac_control_lmacaddr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_9_FFY_RST,
      O => mac_control_lmacaddr(8)
    );
  rxbp_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_1_FFX_RST
    );
  rx_input_memio_BPOUT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_1_68,
      CE => rxbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_1_FFX_RST,
      O => rxbp(1)
    );
  rxbp_1_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxbp_1_CEMUXNOT
    );
  rx_input_fifo_fifo_BU303 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1542,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1549_FFY_RST,
      O => rx_input_fifo_fifo_N1549
    );
  rx_input_fifo_fifo_N1549_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1549_FFY_RST
    );
  rxbp_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_3_FFY_RST
    );
  rx_input_memio_BPOUT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_2_67,
      CE => rxbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_3_FFY_RST,
      O => rxbp(2)
    );
  rxbp_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_3_FFX_RST
    );
  rx_input_memio_BPOUT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_3_66,
      CE => rxbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_3_FFX_RST,
      O => rxbp(3)
    );
  rxbp_3_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxbp_3_CEMUXNOT
    );
  rxbp_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_5_FFY_RST
    );
  rx_input_memio_BPOUT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_4_65,
      CE => rxbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_5_FFY_RST,
      O => rxbp(4)
    );
  rxbp_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_5_FFX_RST
    );
  rx_input_memio_BPOUT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_5_64,
      CE => rxbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_5_FFX_RST,
      O => rxbp(5)
    );
  rxbp_5_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxbp_5_CEMUXNOT
    );
  rxbp_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_7_FFY_RST
    );
  rx_input_memio_BPOUT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_6_63,
      CE => rxbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_7_FFY_RST,
      O => rxbp(6)
    );
  rxbp_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_7_FFX_RST
    );
  rx_input_memio_BPOUT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_7_62,
      CE => rxbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_7_FFX_RST,
      O => rxbp(7)
    );
  rxbp_7_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxbp_7_CEMUXNOT
    );
  rxbp_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_9_FFY_RST
    );
  rx_input_memio_BPOUT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_8_61,
      CE => rxbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_9_FFY_RST,
      O => rxbp(8)
    );
  rxbp_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_9_FFX_RST
    );
  rx_input_memio_BPOUT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_9_60,
      CE => rxbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_9_FFX_RST,
      O => rxbp(9)
    );
  rxbp_9_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxbp_9_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_1_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(0),
      CE => rx_input_memio_addrchk_macaddrl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_1_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(0)
    );
  rx_input_memio_addrchk_macaddrl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_1_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(1),
      CE => rx_input_memio_addrchk_macaddrl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_1_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(1)
    );
  rx_input_memio_addrchk_macaddrl_1_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_1_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_3_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(2),
      CE => rx_input_memio_addrchk_macaddrl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_3_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(2)
    );
  rx_input_memio_addrchk_macaddrl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_3_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(3),
      CE => rx_input_memio_addrchk_macaddrl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_3_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(3)
    );
  rx_input_memio_addrchk_macaddrl_3_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_3_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_5_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(4),
      CE => rx_input_memio_addrchk_macaddrl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_5_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(4)
    );
  rx_input_memio_addrchk_macaddrl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_5_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(5),
      CE => rx_input_memio_addrchk_macaddrl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_5_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(5)
    );
  rx_input_memio_addrchk_macaddrl_5_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_5_CEMUXNOT
    );
  mac_control_Mmux_n0016_Result_28_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cntl(28),
      ADR1 => mac_control_n0065,
      ADR2 => mac_control_n00851_1,
      ADR3 => mac_control_phyaddr(28),
      O => mac_control_CHOICE2250_FROM
    );
  mac_control_Mmux_n0016_Result_7_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_n0065,
      ADR2 => mac_control_rxphyerr_cntl(7),
      ADR3 => mac_control_phyaddr(7),
      O => mac_control_CHOICE2250_GROM
    );
  mac_control_CHOICE2250_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2250_FROM,
      O => mac_control_CHOICE2250
    );
  mac_control_CHOICE2250_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2250_GROM,
      O => mac_control_CHOICE2465
    );
  rx_input_fifo_fifo_BU332 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N5,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1576_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1576
    );
  rx_input_fifo_fifo_N1576_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1576_FFX_SET
    );
  mac_control_Mmux_n0016_Result_6_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_N81078,
      ADR1 => mac_control_CHOICE2698,
      ADR2 => mac_control_CHOICE2689,
      ADR3 => mac_control_CHOICE2686,
      O => mac_control_CHOICE2701_FROM
    );
  mac_control_Mmux_n0016_Result_6_60 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_phystat(6),
      ADR1 => VCC,
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_CHOICE2701,
      O => mac_control_CHOICE2701_GROM
    );
  mac_control_CHOICE2701_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2701_FROM,
      O => mac_control_CHOICE2701
    );
  mac_control_CHOICE2701_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2701_GROM,
      O => mac_control_CHOICE2703
    );
  tx_output_crc_loigc_Mxor_CO_14_Xo_3_1_SW0 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(6),
      ADR1 => tx_output_crcl(28),
      ADR2 => tx_output_data(3),
      ADR3 => tx_output_data(5),
      O => tx_output_crc_loigc_N81257_FROM
    );
  tx_output_crc_loigc_Mxor_n0003_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_data(5),
      ADR3 => tx_output_crcl(26),
      O => tx_output_crc_loigc_N81257_GROM
    );
  tx_output_crc_loigc_N81257_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_N81257_FROM,
      O => tx_output_crc_loigc_N81257
    );
  tx_output_crc_loigc_N81257_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_N81257_GROM,
      O => tx_output_crc_loigc_n0118(1)
    );
  tx_output_ncrcbyte_7_10 : X_LUT4
    generic map(
      INIT => X"30BA"
    )
    port map (
      ADR0 => tx_output_crcsell(2),
      ADR1 => tx_output_crcl(31),
      ADR2 => tx_output_crcsell(3),
      ADR3 => tx_output_crcl(23),
      O => tx_output_CHOICE1439_FROM
    );
  tx_output_crc_loigc_Mxor_n0011_Result1 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => tx_output_data(0),
      ADR1 => VCC,
      ADR2 => tx_output_crcl(31),
      ADR3 => VCC,
      O => tx_output_CHOICE1439_GROM
    );
  tx_output_CHOICE1439_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1439_FROM,
      O => tx_output_CHOICE1439
    );
  tx_output_CHOICE1439_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1439_GROM,
      O => tx_output_crc_loigc_n0124(0)
    );
  mac_control_Mmux_n0016_Result_7_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cntl(7),
      ADR1 => mac_control_n0061,
      ADR2 => mac_control_rxoferr_cntl(7),
      ADR3 => mac_control_n0066,
      O => mac_control_CHOICE2469_FROM
    );
  mac_control_Mmux_n0016_Result_7_45_SW0 : X_LUT4
    generic map(
      INIT => X"FFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0059,
      ADR2 => mac_control_phydi(7),
      ADR3 => mac_control_CHOICE2469,
      O => mac_control_CHOICE2469_GROM
    );
  mac_control_CHOICE2469_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2469_FROM,
      O => mac_control_CHOICE2469
    );
  mac_control_CHOICE2469_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2469_GROM,
      O => mac_control_N81150
    );
  mac_control_Mmux_n0016_Result_7_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2465,
      ADR1 => mac_control_N81150,
      ADR2 => mac_control_CHOICE2461,
      ADR3 => mac_control_CHOICE2458,
      O => mac_control_CHOICE2472_FROM
    );
  mac_control_Mmux_n0016_Result_7_56 : X_LUT4
    generic map(
      INIT => X"FF88"
    )
    port map (
      ADR0 => mac_control_phystat(7),
      ADR1 => mac_control_n0057,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2472,
      O => mac_control_CHOICE2472_GROM
    );
  mac_control_CHOICE2472_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2472_FROM,
      O => mac_control_CHOICE2472
    );
  mac_control_CHOICE2472_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2472_GROM,
      O => mac_control_CHOICE2474
    );
  mac_control_Mmux_n0016_Result_8_22 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxf_cntl(8),
      ADR1 => mac_control_txf_cntl(8),
      ADR2 => mac_control_n0062,
      ADR3 => mac_control_n0061,
      O => mac_control_CHOICE2719_FROM
    );
  mac_control_Mmux_n0016_Result_8_48_SW0 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_n0067,
      ADR1 => mac_control_rxcrcerr_cntl(8),
      ADR2 => mac_control_n0056,
      ADR3 => mac_control_CHOICE2719,
      O => mac_control_CHOICE2719_GROM
    );
  mac_control_CHOICE2719_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2719_FROM,
      O => mac_control_CHOICE2719
    );
  mac_control_CHOICE2719_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2719_GROM,
      O => mac_control_N81066
    );
  mac_control_Mmux_n0016_Result_24_30 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cntl(24),
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_phyaddr(24),
      ADR3 => mac_control_n00851_1,
      O => mac_control_CHOICE2396_FROM
    );
  mac_control_Mmux_n0016_Result_8_30 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_txfifowerr_cntl(8),
      ADR2 => mac_control_phyaddr(8),
      ADR3 => mac_control_n0063,
      O => mac_control_CHOICE2396_GROM
    );
  mac_control_CHOICE2396_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2396_FROM,
      O => mac_control_CHOICE2396
    );
  mac_control_CHOICE2396_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2396_GROM,
      O => mac_control_CHOICE2724
    );
  mac_control_Mmux_n0016_Result_26_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cntl(26),
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_n0064,
      ADR3 => mac_control_rxfifowerr_cntl(26),
      O => mac_control_CHOICE2177_FROM
    );
  mac_control_Mmux_n0016_Result_9_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_txfifowerr_cntl(9),
      ADR2 => mac_control_rxfifowerr_cntl(9),
      ADR3 => mac_control_n0063,
      O => mac_control_CHOICE2177_GROM
    );
  mac_control_CHOICE2177_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2177_FROM,
      O => mac_control_CHOICE2177
    );
  mac_control_CHOICE2177_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2177_GROM,
      O => mac_control_CHOICE2511
    );
  mac_control_Mmux_n0016_Result_12_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0065,
      ADR1 => mac_control_n00851_1,
      ADR2 => mac_control_phyaddr(12),
      ADR3 => mac_control_rxphyerr_cntl(12),
      O => mac_control_CHOICE2540_FROM
    );
  mac_control_Mmux_n0016_Result_9_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_n0065,
      ADR2 => mac_control_rxphyerr_cntl(9),
      ADR3 => mac_control_phyaddr(9),
      O => mac_control_CHOICE2540_GROM
    );
  mac_control_CHOICE2540_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2540_FROM,
      O => mac_control_CHOICE2540
    );
  mac_control_CHOICE2540_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2540_GROM,
      O => mac_control_CHOICE2515
    );
  mac_control_Mmux_n0016_Result_8_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2712,
      ADR1 => mac_control_CHOICE2715,
      ADR2 => mac_control_CHOICE2724,
      ADR3 => mac_control_N81066,
      O => mac_control_CHOICE2727_FROM
    );
  mac_control_Mmux_n0016_Result_8_60 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_phystat(8),
      ADR1 => VCC,
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_CHOICE2727,
      O => mac_control_CHOICE2727_GROM
    );
  mac_control_CHOICE2727_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2727_FROM,
      O => mac_control_CHOICE2727
    );
  mac_control_CHOICE2727_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2727_GROM,
      O => mac_control_CHOICE2729
    );
  mac_control_Mmux_n0016_Result_9_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cntl(9),
      ADR1 => mac_control_n0061,
      ADR2 => mac_control_n0066,
      ADR3 => mac_control_rxoferr_cntl(9),
      O => mac_control_CHOICE2519_FROM
    );
  mac_control_Mmux_n0016_Result_9_45_SW0 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_n0059,
      ADR1 => VCC,
      ADR2 => mac_control_phydi(9),
      ADR3 => mac_control_CHOICE2519,
      O => mac_control_CHOICE2519_GROM
    );
  mac_control_CHOICE2519_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2519_FROM,
      O => mac_control_CHOICE2519
    );
  mac_control_CHOICE2519_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2519_GROM,
      O => mac_control_N81114
    );
  mac_control_Mmux_n0016_Result_9_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2511,
      ADR1 => mac_control_N81114,
      ADR2 => mac_control_CHOICE2515,
      ADR3 => mac_control_CHOICE2508,
      O => mac_control_CHOICE2522_FROM
    );
  mac_control_Mmux_n0016_Result_9_56 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_n0057,
      ADR1 => VCC,
      ADR2 => mac_control_phystat(9),
      ADR3 => mac_control_CHOICE2522,
      O => mac_control_CHOICE2522_GROM
    );
  mac_control_CHOICE2522_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2522_FROM,
      O => mac_control_CHOICE2522
    );
  mac_control_CHOICE2522_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2522_GROM,
      O => mac_control_CHOICE2524
    );
  rx_output_cs_FFd10_In9 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_output_cs_FFd7,
      ADR1 => rx_output_cs_FFd9,
      ADR2 => rx_output_cs_FFd6,
      ADR3 => rx_output_cs_FFd8,
      O => rx_output_CHOICE1800_FROM
    );
  rx_output_cs_Out64 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_output_cs_FFd1,
      ADR1 => rx_output_cs_FFd2,
      ADR2 => rx_output_cs_FFd6,
      ADR3 => rx_output_cs_FFd3,
      O => rx_output_CHOICE1800_GROM
    );
  rx_output_CHOICE1800_XUSED : X_BUF
    port map (
      I => rx_output_CHOICE1800_FROM,
      O => rx_output_CHOICE1800
    );
  rx_output_CHOICE1800_YUSED : X_BUF
    port map (
      I => rx_output_CHOICE1800_GROM,
      O => rx_output_CHOICE876
    );
  rx_output_denl_LOGIC_ZERO_50 : X_ZERO
    port map (
      O => rx_output_denl_LOGIC_ZERO
    );
  rx_output_cs_Out68 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_cs_FFd8,
      ADR2 => rx_output_cs_FFd7,
      ADR3 => rx_output_cs_FFd5,
      O => rx_output_denl_FROM
    );
  rx_output_cs_Out610 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_cs_FFd4,
      ADR2 => rx_output_cs_FFd9,
      ADR3 => rx_output_CHOICE879,
      O => rx_output_CHOICE880
    );
  rx_output_denl_XUSED : X_BUF
    port map (
      I => rx_output_denl_FROM,
      O => rx_output_CHOICE879
    );
  rxbcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbcast_FFY_RST
    );
  mac_control_RXBCAST : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lrxbcast,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbcast_FFY_RST,
      O => rxbcast
    );
  mac_control_PHY_status_MII_Interface_sts28_SW0 : X_LUT4
    generic map(
      INIT => X"77FF"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(1),
      O => mac_control_PHY_status_MII_Interface_N81159_FROM
    );
  mac_control_PHY_status_MII_Interface_sout12 : X_LUT4
    generic map(
      INIT => X"C840"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR2 => mac_control_PHY_status_din(11),
      ADR3 => mac_control_PHY_status_din(3),
      O => mac_control_PHY_status_MII_Interface_N81159_GROM
    );
  mac_control_PHY_status_MII_Interface_N81159_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81159_FROM,
      O => mac_control_PHY_status_MII_Interface_N81159
    );
  mac_control_PHY_status_MII_Interface_N81159_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81159_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE886
    );
  mac_control_PHY_status_MII_Interface_sout27 : X_LUT4
    generic map(
      INIT => X"4450"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR1 => mac_control_PHY_status_din(7),
      ADR2 => mac_control_PHY_status_din(15),
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(3),
      O => mac_control_PHY_status_MII_Interface_CHOICE892_FROM
    );
  mac_control_PHY_status_MII_Interface_sout73 : X_LUT4
    generic map(
      INIT => X"CFCE"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_CHOICE886,
      ADR1 => mac_control_PHY_status_MII_Interface_CHOICE901,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE892,
      O => mac_control_PHY_status_MII_Interface_CHOICE892_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE892_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE892_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE892
    );
  mac_control_PHY_status_MII_Interface_CHOICE892_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE892_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE902
    );
  mac_control_PHY_status_MII_Interface_sout63 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(2),
      O => mac_control_PHY_status_MII_Interface_CHOICE900_FROM
    );
  mac_control_PHY_status_MII_Interface_sout68 : X_LUT4
    generic map(
      INIT => X"D800"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_din(2),
      ADR2 => mac_control_PHY_status_din(10),
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE900,
      O => mac_control_PHY_status_MII_Interface_CHOICE900_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE900_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE900_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE900
    );
  mac_control_PHY_status_MII_Interface_CHOICE900_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE900_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE901
    );
  tx_input_cs_Out51 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_cs_FFd6,
      ADR2 => tx_input_cs_FFd11,
      ADR3 => tx_input_cs_FFd4,
      O => tx_input_mrw_GROM
    );
  tx_input_mrw_YUSED : X_BUF
    port map (
      I => tx_input_mrw_GROM,
      O => tx_input_mrw
    );
  rx_input_memio_addrchk_n00504 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(40),
      ADR1 => rx_input_memio_addrchk_datal(41),
      ADR2 => rx_input_memio_addrchk_datal(42),
      ADR3 => rx_input_memio_addrchk_datal(43),
      O => rx_input_memio_addrchk_CHOICE1525_FROM
    );
  rx_input_memio_addrchk_n004911 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(40),
      ADR1 => rx_input_memio_addrchk_datal(41),
      ADR2 => rx_input_memio_addrchk_datal(42),
      ADR3 => rx_input_memio_addrchk_datal(43),
      O => rx_input_memio_addrchk_CHOICE1525_GROM
    );
  rx_input_memio_addrchk_CHOICE1525_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1525_FROM,
      O => rx_input_memio_addrchk_CHOICE1525
    );
  rx_input_memio_addrchk_CHOICE1525_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1525_GROM,
      O => rx_input_memio_addrchk_CHOICE1535
    );
  rx_input_memio_addrchk_n004924 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(44),
      ADR1 => rx_input_memio_addrchk_datal(45),
      ADR2 => rx_input_memio_addrchk_datal(47),
      ADR3 => rx_input_memio_addrchk_datal(46),
      O => rx_input_memio_addrchk_mcast_0_FROM
    );
  rx_input_memio_addrchk_n004925 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_CHOICE1535,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1542,
      O => rx_input_memio_addrchk_lmcast(0)
    );
  rx_input_memio_addrchk_mcast_0_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_mcast_0_CEMUXNOT
    );
  rx_input_memio_addrchk_mcast_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_mcast_0_FROM,
      O => rx_input_memio_addrchk_CHOICE1542
    );
  tx_output_ncrcbyte_2_10 : X_LUT4
    generic map(
      INIT => X"0CAE"
    )
    port map (
      ADR0 => tx_output_crcsell(3),
      ADR1 => tx_output_crcsell(2),
      ADR2 => tx_output_crcl(18),
      ADR3 => tx_output_crcl(26),
      O => tx_output_CHOICE1505_FROM
    );
  tx_output_ncrcbyte_0_10 : X_LUT4
    generic map(
      INIT => X"2F22"
    )
    port map (
      ADR0 => tx_output_crcsell(2),
      ADR1 => tx_output_crcl(16),
      ADR2 => tx_output_crcl(24),
      ADR3 => tx_output_crcsell(3),
      O => tx_output_CHOICE1505_GROM
    );
  tx_output_CHOICE1505_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1505_FROM,
      O => tx_output_CHOICE1505
    );
  tx_output_CHOICE1505_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1505_GROM,
      O => tx_output_CHOICE1516
    );
  tx_output_ncrcbyte_0_21 : X_LUT4
    generic map(
      INIT => X"30BA"
    )
    port map (
      ADR0 => tx_output_crcsell(1),
      ADR1 => tx_output_crcl(0),
      ADR2 => tx_output_crcsell(0),
      ADR3 => tx_output_crcl(8),
      O => tx_output_ncrcbytel_0_FROM
    );
  tx_output_ncrcbyte_0_22 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_CHOICE1516,
      ADR3 => tx_output_CHOICE1521,
      O => tx_output_ncrcbyte(0)
    );
  tx_output_ncrcbytel_0_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_ncrcbytel_0_CEMUXNOT
    );
  tx_output_ncrcbytel_0_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_0_FROM,
      O => tx_output_CHOICE1521
    );
  mac_control_PHY_status_dout_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_13_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(12),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_13_FFY_RST,
      O => mac_control_PHY_status_dout(12)
    );
  mac_control_PHY_status_dout_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_15_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(14),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_15_FFY_RST,
      O => mac_control_PHY_status_dout(14)
    );
  tx_output_ncrcbyte_3_10 : X_LUT4
    generic map(
      INIT => X"4F44"
    )
    port map (
      ADR0 => tx_output_crcl(19),
      ADR1 => tx_output_crcsell(2),
      ADR2 => tx_output_crcl(27),
      ADR3 => tx_output_crcsell(3),
      O => tx_output_CHOICE1483_FROM
    );
  tx_output_ncrcbyte_1_10 : X_LUT4
    generic map(
      INIT => X"2F22"
    )
    port map (
      ADR0 => tx_output_crcsell(3),
      ADR1 => tx_output_crcl(25),
      ADR2 => tx_output_crcl(17),
      ADR3 => tx_output_crcsell(2),
      O => tx_output_CHOICE1483_GROM
    );
  tx_output_CHOICE1483_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1483_FROM,
      O => tx_output_CHOICE1483
    );
  tx_output_CHOICE1483_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1483_GROM,
      O => tx_output_CHOICE1494
    );
  tx_output_ncrcbyte_1_21 : X_LUT4
    generic map(
      INIT => X"0ACE"
    )
    port map (
      ADR0 => tx_output_crcsell(0),
      ADR1 => tx_output_crcsell(1),
      ADR2 => tx_output_crcl(1),
      ADR3 => tx_output_crcl(9),
      O => tx_output_ncrcbytel_1_FROM
    );
  tx_output_ncrcbyte_1_22 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_CHOICE1494,
      ADR3 => tx_output_CHOICE1499,
      O => tx_output_ncrcbyte(1)
    );
  tx_output_ncrcbytel_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_ncrcbytel_1_CEMUXNOT
    );
  tx_output_ncrcbytel_1_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_1_FROM,
      O => tx_output_CHOICE1499
    );
  tx_output_ncrcbyte_2_21 : X_LUT4
    generic map(
      INIT => X"50DC"
    )
    port map (
      ADR0 => tx_output_crcl(10),
      ADR1 => tx_output_crcsell(0),
      ADR2 => tx_output_crcsell(1),
      ADR3 => tx_output_crcl(2),
      O => tx_output_ncrcbytel_2_FROM
    );
  tx_output_ncrcbyte_2_22 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_CHOICE1505,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1510,
      O => tx_output_ncrcbyte(2)
    );
  tx_output_ncrcbytel_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_ncrcbytel_2_CEMUXNOT
    );
  tx_output_ncrcbytel_2_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_2_FROM,
      O => tx_output_CHOICE1510
    );
  tx_output_ncrcbyte_3_21 : X_LUT4
    generic map(
      INIT => X"4F44"
    )
    port map (
      ADR0 => tx_output_crcl(3),
      ADR1 => tx_output_crcsell(0),
      ADR2 => tx_output_crcl(11),
      ADR3 => tx_output_crcsell(1),
      O => tx_output_ncrcbytel_3_FROM
    );
  tx_output_ncrcbyte_3_22 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_CHOICE1483,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1488,
      O => tx_output_ncrcbyte(3)
    );
  tx_output_ncrcbytel_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_ncrcbytel_3_CEMUXNOT
    );
  tx_output_ncrcbytel_3_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_3_FROM,
      O => tx_output_CHOICE1488
    );
  rx_input_fifo_fifo_BU406 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N1562_FROM,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1562_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1562
    );
  rx_input_fifo_fifo_N1562_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1562_FFX_SET
    );
  tx_output_ncrcbyte_6_10 : X_LUT4
    generic map(
      INIT => X"7350"
    )
    port map (
      ADR0 => tx_output_crcl(30),
      ADR1 => tx_output_crcl(22),
      ADR2 => tx_output_crcsell(3),
      ADR3 => tx_output_crcsell(2),
      O => tx_output_CHOICE1450_FROM
    );
  tx_output_ncrcbyte_4_10 : X_LUT4
    generic map(
      INIT => X"3B0A"
    )
    port map (
      ADR0 => tx_output_crcsell(2),
      ADR1 => tx_output_crcl(28),
      ADR2 => tx_output_crcl(20),
      ADR3 => tx_output_crcsell(3),
      O => tx_output_CHOICE1450_GROM
    );
  tx_output_CHOICE1450_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1450_FROM,
      O => tx_output_CHOICE1450
    );
  tx_output_CHOICE1450_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1450_GROM,
      O => tx_output_CHOICE1461
    );
  rx_input_memio_crccomb_Mxor_n0007_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(29),
      ADR1 => rx_input_memio_datal(6),
      ADR2 => rx_input_memio_datal(2),
      ADR3 => rx_input_memio_crcl(25),
      O => rx_input_memio_crccomb_Mxor_n0007_Xo_0_FROM
    );
  rx_input_memio_crccomb_Mxor_n0021_Result1 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_input_memio_crcl(29),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_datal(2),
      O => rx_input_memio_crccomb_Mxor_n0007_Xo_0_GROM
    );
  rx_input_memio_crccomb_Mxor_n0007_Xo_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_n0007_Xo_0_FROM,
      O => rx_input_memio_crccomb_Mxor_n0007_Xo(0)
    );
  rx_input_memio_crccomb_Mxor_n0007_Xo_0_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_n0007_Xo_0_GROM,
      O => rx_input_memio_crccomb_n0118(0)
    );
  tx_output_ncrcbyte_4_21 : X_LUT4
    generic map(
      INIT => X"2F22"
    )
    port map (
      ADR0 => tx_output_crcsell(1),
      ADR1 => tx_output_crcl(12),
      ADR2 => tx_output_crcl(4),
      ADR3 => tx_output_crcsell(0),
      O => tx_output_ncrcbytel_4_FROM
    );
  tx_output_ncrcbyte_4_22 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_CHOICE1461,
      ADR3 => tx_output_CHOICE1466,
      O => tx_output_ncrcbyte(4)
    );
  tx_output_ncrcbytel_4_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_ncrcbytel_4_CEMUXNOT
    );
  tx_output_ncrcbytel_4_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_4_FROM,
      O => tx_output_CHOICE1466
    );
  tx_output_crc_loigc_Mxor_n0021_Result1 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_data(2),
      ADR2 => VCC,
      ADR3 => tx_output_crcl(29),
      O => tx_output_crc_loigc_n0118_0_FROM
    );
  tx_output_ncrcbyte_5_10 : X_LUT4
    generic map(
      INIT => X"2F22"
    )
    port map (
      ADR0 => tx_output_crcsell(2),
      ADR1 => tx_output_crcl(21),
      ADR2 => tx_output_crcl(29),
      ADR3 => tx_output_crcsell(3),
      O => tx_output_crc_loigc_n0118_0_GROM
    );
  tx_output_crc_loigc_n0118_0_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0118_0_FROM,
      O => tx_output_crc_loigc_n0118(0)
    );
  tx_output_crc_loigc_n0118_0_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0118_0_GROM,
      O => tx_output_CHOICE1472
    );
  rx_input_fifo_fifo_BU237 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N3039,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1586_FFY_RST,
      O => rx_input_fifo_fifo_N1585
    );
  rx_input_fifo_fifo_N1586_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1586_FFY_RST
    );
  tx_output_crc_loigc_Mxor_n0004_Result1 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => tx_output_crcl(27),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_data(4),
      O => tx_output_crc_loigc_n0124_1_GROM
    );
  tx_output_crc_loigc_n0124_1_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0124_1_GROM,
      O => tx_output_crc_loigc_n0124(1)
    );
  tx_output_ncrcbyte_5_21 : X_LUT4
    generic map(
      INIT => X"7350"
    )
    port map (
      ADR0 => tx_output_crcl(13),
      ADR1 => tx_output_crcl(5),
      ADR2 => tx_output_crcsell(1),
      ADR3 => tx_output_crcsell(0),
      O => tx_output_ncrcbytel_5_FROM
    );
  tx_output_ncrcbyte_5_22 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_CHOICE1472,
      ADR2 => VCC,
      ADR3 => tx_output_CHOICE1477,
      O => tx_output_ncrcbyte(5)
    );
  tx_output_ncrcbytel_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_ncrcbytel_5_CEMUXNOT
    );
  tx_output_ncrcbytel_5_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_5_FROM,
      O => tx_output_CHOICE1477
    );
  tx_output_ncrcbyte_6_21 : X_LUT4
    generic map(
      INIT => X"2F22"
    )
    port map (
      ADR0 => tx_output_crcsell(0),
      ADR1 => tx_output_crcl(6),
      ADR2 => tx_output_crcl(14),
      ADR3 => tx_output_crcsell(1),
      O => tx_output_ncrcbytel_6_FROM
    );
  tx_output_ncrcbyte_6_22 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_CHOICE1450,
      ADR3 => tx_output_CHOICE1455,
      O => tx_output_ncrcbyte(6)
    );
  tx_output_ncrcbytel_6_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_ncrcbytel_6_CEMUXNOT
    );
  tx_output_ncrcbytel_6_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_6_FROM,
      O => tx_output_CHOICE1455
    );
  tx_output_ncrcbyte_7_21 : X_LUT4
    generic map(
      INIT => X"5D0C"
    )
    port map (
      ADR0 => tx_output_crcl(15),
      ADR1 => tx_output_crcsell(0),
      ADR2 => tx_output_crcl(7),
      ADR3 => tx_output_crcsell(1),
      O => tx_output_ncrcbytel_7_FROM
    );
  tx_output_ncrcbyte_7_22 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_CHOICE1439,
      ADR3 => tx_output_CHOICE1444,
      O => tx_output_ncrcbyte(7)
    );
  tx_output_ncrcbytel_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_ncrcbytel_7_CEMUXNOT
    );
  tx_output_ncrcbytel_7_XUSED : X_BUF
    port map (
      I => tx_output_ncrcbytel_7_FROM,
      O => tx_output_CHOICE1444
    );
  mac_control_rxf_cntl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_11_FFY_RST
    );
  mac_control_rxf_cntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(10),
      CE => mac_control_rxf_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_11_FFY_RST,
      O => mac_control_rxf_cntl(10)
    );
  mac_control_rxf_cntl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_11_CEMUXNOT
    );
  rx_input_fifo_fifo_BU192 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2685,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N8_FFY_RST,
      O => rx_input_fifo_fifo_N7
    );
  rx_input_fifo_fifo_N8_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N8_FFY_RST
    );
  mac_control_rxf_cntl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_21_FFY_RST
    );
  mac_control_rxf_cntl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(20),
      CE => mac_control_rxf_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_21_FFY_RST,
      O => mac_control_rxf_cntl(20)
    );
  mac_control_rxf_cntl_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_21_CEMUXNOT
    );
  mac_control_rxf_cntl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_13_FFY_RST
    );
  mac_control_rxf_cntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(12),
      CE => mac_control_rxf_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_13_FFY_RST,
      O => mac_control_rxf_cntl(12)
    );
  mac_control_rxf_cntl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_13_CEMUXNOT
    );
  rx_input_fifo_fifo_BU230 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2999,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1586_FFX_RST,
      O => rx_input_fifo_fifo_N1586
    );
  rx_input_fifo_fifo_N1586_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1586_FFX_RST
    );
  mac_control_rxf_cntl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_31_FFY_RST
    );
  mac_control_rxf_cntl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(30),
      CE => mac_control_rxf_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_31_FFY_RST,
      O => mac_control_rxf_cntl(30)
    );
  mac_control_rxf_cntl_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_31_CEMUXNOT
    );
  mac_control_rxf_cntl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_23_FFY_RST
    );
  mac_control_rxf_cntl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(22),
      CE => mac_control_rxf_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_23_FFY_RST,
      O => mac_control_rxf_cntl(22)
    );
  mac_control_rxf_cntl_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_23_CEMUXNOT
    );
  mac_control_rxf_cntl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_15_FFY_RST
    );
  mac_control_rxf_cntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(14),
      CE => mac_control_rxf_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_15_FFY_RST,
      O => mac_control_rxf_cntl(14)
    );
  mac_control_rxf_cntl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_15_CEMUXNOT
    );
  mac_control_rxf_cntl_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_25_CEMUXNOT
    );
  mac_control_rxf_cntl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_17_FFY_RST
    );
  mac_control_rxf_cntl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(16),
      CE => mac_control_rxf_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_17_FFY_RST,
      O => mac_control_rxf_cntl(16)
    );
  mac_control_rxf_cntl_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_17_CEMUXNOT
    );
  mac_control_rxf_cntl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_27_FFY_RST
    );
  mac_control_rxf_cntl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(26),
      CE => mac_control_rxf_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_27_FFY_RST,
      O => mac_control_rxf_cntl(26)
    );
  mac_control_rxf_cntl_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_27_CEMUXNOT
    );
  mac_control_rxf_cntl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_19_FFY_RST
    );
  mac_control_rxf_cntl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(18),
      CE => mac_control_rxf_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_19_FFY_RST,
      O => mac_control_rxf_cntl(18)
    );
  mac_control_rxf_cntl_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_19_CEMUXNOT
    );
  mac_control_rxf_cntl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_29_FFY_RST
    );
  mac_control_rxf_cntl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(28),
      CE => mac_control_rxf_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_29_FFY_RST,
      O => mac_control_rxf_cntl(28)
    );
  mac_control_rxf_cntl_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_29_CEMUXNOT
    );
  rx_fifocheck_n000212 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(0),
      ADR1 => rx_fifocheck_diff(2),
      ADR2 => rx_fifocheck_diff(1),
      ADR3 => rx_fifocheck_diff(3),
      O => rx_fifocheck_CHOICE1950_GROM
    );
  rx_fifocheck_CHOICE1950_YUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1950_GROM,
      O => rx_fifocheck_CHOICE1950
    );
  rx_fifocheck_n000225 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(4),
      ADR1 => rx_fifocheck_diff(5),
      ADR2 => rx_fifocheck_diff(7),
      ADR3 => rx_fifocheck_diff(6),
      O => rx_fifocheck_CHOICE1957_GROM
    );
  rx_fifocheck_CHOICE1957_YUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1957_GROM,
      O => rx_fifocheck_CHOICE1957
    );
  mac_control_Mmux_n0016_Result_10_97_SW1 : X_LUT4
    generic map(
      INIT => X"AABF"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_phydo(10),
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_CHOICE2755,
      O => mac_control_dout_10_FROM
    );
  mac_control_Mmux_n0016_Result_10_97 : X_LUT4
    generic map(
      INIT => X"2AEA"
    )
    port map (
      ADR0 => mac_control_dout(9),
      ADR1 => mac_control_sclkdeltall,
      ADR2 => mac_control_n0086,
      ADR3 => mac_control_N81463,
      O => mac_control_n0016(10)
    );
  mac_control_dout_10_XUSED : X_BUF
    port map (
      I => mac_control_dout_10_FROM,
      O => mac_control_N81463
    );
  rx_fifocheck_n000262 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(13),
      ADR1 => rx_fifocheck_diff(12),
      ADR2 => rx_fifocheck_diff(15),
      ADR3 => rx_fifocheck_diff(14),
      O => rx_fifocheck_CHOICE1972_GROM
    );
  rx_fifocheck_CHOICE1972_YUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1972_GROM,
      O => rx_fifocheck_CHOICE1972
    );
  rx_fifocheck_n000263 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_fifocheck_CHOICE1972,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_CHOICE1965,
      O => rx_fifocheck_CHOICE1973_FROM
    );
  rx_fifocheck_n000292 : X_LUT4
    generic map(
      INIT => X"F8F0"
    )
    port map (
      ADR0 => rx_fifocheck_CHOICE1950,
      ADR1 => rx_fifocheck_CHOICE1957,
      ADR2 => rx_fifocheck_n0003,
      ADR3 => rx_fifocheck_CHOICE1973,
      O => rx_fifocheck_CHOICE1973_GROM
    );
  rx_fifocheck_CHOICE1973_XUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1973_FROM,
      O => rx_fifocheck_CHOICE1973
    );
  rx_fifocheck_CHOICE1973_YUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1973_GROM,
      O => rx_fifocheck_n0002
    );
  rx_fifocheck_n000249 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(9),
      ADR1 => rx_fifocheck_diff(8),
      ADR2 => rx_fifocheck_diff(11),
      ADR3 => rx_fifocheck_diff(10),
      O => rx_fifocheck_CHOICE1965_GROM
    );
  rx_fifocheck_CHOICE1965_YUSED : X_BUF
    port map (
      I => rx_fifocheck_CHOICE1965_GROM,
      O => rx_fifocheck_CHOICE1965
    );
  mac_control_Mmux_n0016_Result_20_45_SW0 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_phydi(20),
      ADR1 => VCC,
      ADR2 => mac_control_n0059,
      ADR3 => mac_control_CHOICE2139,
      O => mac_control_N81102_FROM
    );
  mac_control_Mmux_n0016_Result_20_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2135,
      ADR1 => mac_control_CHOICE2128,
      ADR2 => mac_control_CHOICE2131,
      ADR3 => mac_control_N81102,
      O => mac_control_N81102_GROM
    );
  mac_control_N81102_XUSED : X_BUF
    port map (
      I => mac_control_N81102_FROM,
      O => mac_control_N81102
    );
  mac_control_N81102_YUSED : X_BUF
    port map (
      I => mac_control_N81102_GROM,
      O => mac_control_CHOICE2142
    );
  mac_control_Mmux_n0016_Result_11_93_SW1 : X_LUT4
    generic map(
      INIT => X"ABBB"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_CHOICE2499,
      ADR2 => mac_control_phydo(11),
      ADR3 => mac_control_n0060,
      O => mac_control_dout_11_FROM
    );
  mac_control_Mmux_n0016_Result_11_93 : X_LUT4
    generic map(
      INIT => X"4CEC"
    )
    port map (
      ADR0 => mac_control_sclkdeltall,
      ADR1 => mac_control_dout(10),
      ADR2 => mac_control_n0086,
      ADR3 => mac_control_N81467,
      O => mac_control_n0016(11)
    );
  mac_control_dout_11_XUSED : X_BUF
    port map (
      I => mac_control_dout_11_FROM,
      O => mac_control_N81467
    );
  rx_input_memio_RESET_1_51 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_RESET_1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_RESET_1_FROM
    );
  rx_input_memio_addrchk_n00321 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_RESET_1,
      O => rx_input_memio_RESET_1_GROM
    );
  rx_input_memio_RESET_1_XUSED : X_BUF
    port map (
      I => rx_input_memio_RESET_1_FROM,
      O => rx_input_memio_RESET_1
    );
  rx_input_memio_RESET_1_YUSED : X_BUF
    port map (
      I => rx_input_memio_RESET_1_GROM,
      O => rx_input_memio_addrchk_n0032
    );
  tx_output_n0034_12_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_crc_12_Q,
      ADR2 => VCC,
      ADR3 => tx_output_cs_FFd16,
      O => tx_output_n0034_12_1_O
    );
  tx_output_n00251 : X_LUT4
    generic map(
      INIT => X"0F0A"
    )
    port map (
      ADR0 => tx_output_crcenl,
      ADR1 => VCC,
      ADR2 => RESET_IBUF_2,
      ADR3 => tx_output_cs_FFd16,
      O => tx_output_crcl_12_GROM
    );
  tx_output_crcl_12_YUSED : X_BUF
    port map (
      I => tx_output_crcl_12_GROM,
      O => tx_output_n0025
    );
  tx_output_cs_Out149 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd9,
      ADR1 => tx_output_cs_FFd10,
      ADR2 => tx_output_cs_FFd6_1,
      ADR3 => tx_output_cs_FFd8,
      O => tx_output_CHOICE1775_FROM
    );
  tx_output_cs_Out1132 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_cs_FFd5_1,
      ADR1 => tx_output_cs_FFd13,
      ADR2 => tx_output_cs_FFd10,
      ADR3 => tx_output_cs_FFd11,
      O => tx_output_CHOICE1775_GROM
    );
  tx_output_CHOICE1775_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1775_FROM,
      O => tx_output_CHOICE1775
    );
  tx_output_CHOICE1775_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1775_GROM,
      O => tx_output_CHOICE1760
    );
  tx_output_ldata_4_17 : X_LUT4
    generic map(
      INIT => X"0004"
    )
    port map (
      ADR0 => tx_output_cs_FFd5_1,
      ADR1 => q2(4),
      ADR2 => tx_output_cs_FFd4_1,
      ADR3 => tx_output_cs_FFd6_1,
      O => tx_output_CHOICE1682_FROM
    );
  tx_output_cs_Out1421 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd7,
      ADR1 => tx_output_cs_FFd3,
      ADR2 => tx_output_cs_FFd4_1,
      ADR3 => tx_output_cs_FFd5_1,
      O => tx_output_CHOICE1682_GROM
    );
  tx_output_CHOICE1682_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1682_FROM,
      O => tx_output_CHOICE1682
    );
  tx_output_CHOICE1682_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1682_GROM,
      O => tx_output_CHOICE1779
    );
  tx_output_cs_Out101 : X_LUT4
    generic map(
      INIT => X"0101"
    )
    port map (
      ADR0 => tx_output_cs_FFd3,
      ADR1 => tx_output_cs_FFd2,
      ADR2 => tx_output_cs_FFd7,
      ADR3 => VCC,
      O => tx_output_crcsel(0)
    );
  tx_output_cs_Out1426 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd2,
      ADR1 => tx_output_cs_FFd1,
      ADR2 => tx_output_cs_FFd15,
      ADR3 => tx_output_cs_FFd16,
      O => tx_output_crcsell_0_GROM
    );
  tx_output_crcsell_0_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_crcsell_0_CEMUXNOT
    );
  tx_output_crcsell_0_YUSED : X_BUF
    port map (
      I => tx_output_crcsell_0_GROM,
      O => tx_output_CHOICE1782
    );
  mac_control_rxoferr_cntl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_1_CEMUXNOT
    );
  mac_control_rxoferr_cntl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_3_FFY_RST
    );
  mac_control_rxoferr_cntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(2),
      CE => mac_control_rxoferr_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_3_FFY_RST,
      O => mac_control_rxoferr_cntl(2)
    );
  mac_control_rxoferr_cntl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_3_CEMUXNOT
    );
  mac_control_rxoferr_cntl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_5_FFY_RST
    );
  mac_control_rxoferr_cntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(4),
      CE => mac_control_rxoferr_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_5_FFY_RST,
      O => mac_control_rxoferr_cntl(4)
    );
  mac_control_rxoferr_cntl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_5_CEMUXNOT
    );
  mac_control_rxoferr_cntl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_7_FFY_RST
    );
  mac_control_rxoferr_cntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(6),
      CE => mac_control_rxoferr_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_7_FFY_RST,
      O => mac_control_rxoferr_cntl(6)
    );
  mac_control_rxoferr_cntl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_7_CEMUXNOT
    );
  mac_control_rxoferr_cntl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_9_FFY_RST
    );
  mac_control_rxoferr_cntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(8),
      CE => mac_control_rxoferr_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_9_FFY_RST,
      O => mac_control_rxoferr_cntl(8)
    );
  mac_control_rxoferr_cntl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_9_CEMUXNOT
    );
  mac_control_dout_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_12_FFY_RST
    );
  mac_control_dout_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(12),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_12_FFY_RST,
      O => mac_control_dout(12)
    );
  mac_control_Mmux_n0016_Result_12_93_SW1 : X_LUT4
    generic map(
      INIT => X"AABF"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_phydo(12),
      ADR2 => mac_control_n0060,
      ADR3 => mac_control_CHOICE2549,
      O => mac_control_dout_12_FROM
    );
  mac_control_Mmux_n0016_Result_12_93 : X_LUT4
    generic map(
      INIT => X"2AEA"
    )
    port map (
      ADR0 => mac_control_dout(11),
      ADR1 => mac_control_n0086,
      ADR2 => mac_control_sclkdeltall,
      ADR3 => mac_control_N81471,
      O => mac_control_n0016(12)
    );
  mac_control_dout_12_XUSED : X_BUF
    port map (
      I => mac_control_dout_12_FROM,
      O => mac_control_N81471
    );
  mac_control_Mmux_n0016_Result_21_48_SW0 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cntl(21),
      ADR1 => mac_control_n0067,
      ADR2 => mac_control_n0056,
      ADR3 => mac_control_CHOICE2367,
      O => mac_control_N81038_FROM
    );
  mac_control_Mmux_n0016_Result_21_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2363,
      ADR1 => mac_control_CHOICE2372,
      ADR2 => mac_control_CHOICE2360,
      ADR3 => mac_control_N81038,
      O => mac_control_N81038_GROM
    );
  mac_control_N81038_XUSED : X_BUF
    port map (
      I => mac_control_N81038_FROM,
      O => mac_control_N81038
    );
  mac_control_N81038_YUSED : X_BUF
    port map (
      I => mac_control_N81038_GROM,
      O => mac_control_CHOICE2375
    );
  rx_input_fifo_fifo_BU294 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N1544,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N1550_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1551
    );
  rx_input_fifo_fifo_N1550_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1550_FFY_SET
    );
  tx_output_crc_loigc_Mxor_CO_2_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0118(1),
      ADR1 => tx_output_crc_loigc_n0124(0),
      ADR2 => tx_output_crc_loigc_n0122(0),
      ADR3 => tx_output_crc_0_Q,
      O => tx_output_crcl_2_FROM
    );
  tx_output_n0034_2_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_2_Q,
      O => tx_output_n0034_2_Q
    );
  tx_output_crcl_2_XUSED : X_BUF
    port map (
      I => tx_output_crcl_2_FROM,
      O => tx_output_crc_2_Q
    );
  mac_control_Mmux_n0016_Result_22_45_SW0 : X_LUT4
    generic map(
      INIT => X"EECC"
    )
    port map (
      ADR0 => mac_control_n0059,
      ADR1 => mac_control_CHOICE2116,
      ADR2 => VCC,
      ADR3 => mac_control_phydi(22),
      O => mac_control_N81090_FROM
    );
  mac_control_Mmux_n0016_Result_22_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2108,
      ADR1 => mac_control_CHOICE2105,
      ADR2 => mac_control_CHOICE2112,
      ADR3 => mac_control_N81090,
      O => mac_control_N81090_GROM
    );
  mac_control_N81090_XUSED : X_BUF
    port map (
      I => mac_control_N81090_FROM,
      O => mac_control_N81090
    );
  mac_control_N81090_YUSED : X_BUF
    port map (
      I => mac_control_N81090_GROM,
      O => mac_control_CHOICE2119
    );
  mac_control_Mmux_n0016_Result_30_45_SW0 : X_LUT4
    generic map(
      INIT => X"EAEA"
    )
    port map (
      ADR0 => mac_control_CHOICE2300,
      ADR1 => mac_control_phydi(30),
      ADR2 => mac_control_n0059,
      ADR3 => VCC,
      O => mac_control_N81094_FROM
    );
  mac_control_Mmux_n0016_Result_30_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2292,
      ADR1 => mac_control_CHOICE2296,
      ADR2 => mac_control_CHOICE2289,
      ADR3 => mac_control_N81094,
      O => mac_control_N81094_GROM
    );
  mac_control_N81094_XUSED : X_BUF
    port map (
      I => mac_control_N81094_FROM,
      O => mac_control_N81094
    );
  mac_control_N81094_YUSED : X_BUF
    port map (
      I => mac_control_N81094_GROM,
      O => mac_control_CHOICE2303
    );
  mac_control_Mmux_n0016_Result_13_93_SW1 : X_LUT4
    generic map(
      INIT => X"FF07"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_phydo(13),
      ADR2 => mac_control_CHOICE2574,
      ADR3 => mac_control_addr(5),
      O => mac_control_dout_13_FROM
    );
  mac_control_Mmux_n0016_Result_13_93 : X_LUT4
    generic map(
      INIT => X"70F8"
    )
    port map (
      ADR0 => mac_control_n0086,
      ADR1 => mac_control_sclkdeltall,
      ADR2 => mac_control_dout(12),
      ADR3 => mac_control_N81475,
      O => mac_control_n0016(13)
    );
  mac_control_dout_13_XUSED : X_BUF
    port map (
      I => mac_control_dout_13_FROM,
      O => mac_control_N81475
    );
  rx_input_fifo_fifo_BU186 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2684,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N8_FFX_RST,
      O => rx_input_fifo_fifo_N8
    );
  rx_input_fifo_fifo_N8_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N8_FFX_RST
    );
  mac_control_Mshreg_scslll_103_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_Mshreg_scslll_103_CEMUXNOT
    );
  rx_input_GMII_rx_of_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_GMII_rx_of_FFY_RST
    );
  rx_input_GMII_rx_of_52 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_rx_nearf,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_GMII_rx_of_FFY_RST,
      O => rx_input_GMII_rx_of
    );
  mac_control_Mmux_n0016_Result_26_28 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxoferr_cntl(26),
      ADR1 => mac_control_txf_cntl(26),
      ADR2 => mac_control_n0061,
      ADR3 => mac_control_n0066,
      O => mac_control_CHOICE2185_FROM
    );
  mac_control_Mmux_n0016_Result_31_36_SW0 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0059,
      ADR1 => mac_control_txf_cntl(31),
      ADR2 => mac_control_n0061,
      ADR3 => mac_control_phydi(31),
      O => mac_control_CHOICE2185_GROM
    );
  mac_control_CHOICE2185_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2185_FROM,
      O => mac_control_CHOICE2185
    );
  mac_control_CHOICE2185_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2185_GROM,
      O => mac_control_N80963
    );
  rx_input_fifo_fifo_BU277 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N1530,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N1543_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1544
    );
  rx_input_fifo_fifo_N1543_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1543_FFY_SET
    );
  rx_input_memio_n005915 : X_LUT4
    generic map(
      INIT => X"0080"
    )
    port map (
      ADR0 => rx_input_memio_crcll(4),
      ADR1 => rx_input_memio_crcll(6),
      ADR2 => rx_input_memio_crcll(5),
      ADR3 => rx_input_memio_crcll(7),
      O => rx_input_memio_CHOICE1812_GROM
    );
  rx_input_memio_CHOICE1812_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1812_GROM,
      O => rx_input_memio_CHOICE1812
    );
  mac_control_Mmux_n0016_Result_23_45_SW0 : X_LUT4
    generic map(
      INIT => X"ECEC"
    )
    port map (
      ADR0 => mac_control_phydi(23),
      ADR1 => mac_control_CHOICE2162,
      ADR2 => mac_control_n0059,
      ADR3 => VCC,
      O => mac_control_N81134_FROM
    );
  mac_control_Mmux_n0016_Result_23_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2154,
      ADR1 => mac_control_CHOICE2151,
      ADR2 => mac_control_CHOICE2158,
      ADR3 => mac_control_N81134,
      O => mac_control_N81134_GROM
    );
  mac_control_N81134_XUSED : X_BUF
    port map (
      I => mac_control_N81134_FROM,
      O => mac_control_N81134
    );
  mac_control_N81134_YUSED : X_BUF
    port map (
      I => mac_control_N81134_GROM,
      O => mac_control_CHOICE2165
    );
  rx_input_memio_n005940 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => rx_input_memio_crcll(13),
      ADR1 => rx_input_memio_crcll(12),
      ADR2 => rx_input_memio_crcll(15),
      ADR3 => rx_input_memio_crcll(14),
      O => rx_input_memio_CHOICE1821_FROM
    );
  rx_input_memio_n005941 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_CHOICE1817,
      ADR2 => VCC,
      ADR3 => rx_input_memio_CHOICE1821,
      O => rx_input_memio_CHOICE1821_GROM
    );
  rx_input_memio_CHOICE1821_XUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1821_FROM,
      O => rx_input_memio_CHOICE1821
    );
  rx_input_memio_CHOICE1821_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1821_GROM,
      O => rx_input_memio_CHOICE1822
    );
  rx_input_memio_n005932 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => rx_input_memio_crcll(9),
      ADR1 => rx_input_memio_crcll(8),
      ADR2 => rx_input_memio_crcll(11),
      ADR3 => rx_input_memio_crcll(10),
      O => rx_input_memio_CHOICE1817_GROM
    );
  rx_input_memio_CHOICE1817_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1817_GROM,
      O => rx_input_memio_CHOICE1817
    );
  rx_input_memio_n005979 : X_LUT4
    generic map(
      INIT => X"0040"
    )
    port map (
      ADR0 => rx_input_memio_crcll(28),
      ADR1 => rx_input_memio_crcll(31),
      ADR2 => rx_input_memio_crcll(30),
      ADR3 => rx_input_memio_crcll(29),
      O => rx_input_memio_CHOICE1832_GROM
    );
  rx_input_memio_CHOICE1832_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1832_GROM,
      O => rx_input_memio_CHOICE1832
    );
  mac_control_txfifowerr_cntl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_11_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_21_FFY_RST
    );
  mac_control_txfifowerr_cntl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(20),
      CE => mac_control_txfifowerr_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_21_FFY_RST,
      O => mac_control_txfifowerr_cntl(20)
    );
  mac_control_txfifowerr_cntl_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_21_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_13_FFY_RST
    );
  mac_control_txfifowerr_cntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(12),
      CE => mac_control_txfifowerr_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_13_FFY_RST,
      O => mac_control_txfifowerr_cntl(12)
    );
  mac_control_txfifowerr_cntl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_13_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_31_FFY_RST
    );
  mac_control_txfifowerr_cntl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(30),
      CE => mac_control_txfifowerr_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_31_FFY_RST,
      O => mac_control_txfifowerr_cntl(30)
    );
  mac_control_txfifowerr_cntl_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_31_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_23_FFY_RST
    );
  mac_control_txfifowerr_cntl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(22),
      CE => mac_control_txfifowerr_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_23_FFY_RST,
      O => mac_control_txfifowerr_cntl(22)
    );
  mac_control_txfifowerr_cntl_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_23_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_15_FFY_RST
    );
  mac_control_txfifowerr_cntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(14),
      CE => mac_control_txfifowerr_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_15_FFY_RST,
      O => mac_control_txfifowerr_cntl(14)
    );
  mac_control_txfifowerr_cntl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_15_CEMUXNOT
    );
  mac_control_dout_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_14_FFY_RST
    );
  mac_control_dout_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(14),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_14_FFY_RST,
      O => mac_control_dout(14)
    );
  mac_control_Mmux_n0016_Result_14_97_SW1 : X_LUT4
    generic map(
      INIT => X"F0F7"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_phydo(14),
      ADR2 => mac_control_addr(5),
      ADR3 => mac_control_CHOICE2781,
      O => mac_control_dout_14_FROM
    );
  mac_control_Mmux_n0016_Result_14_97 : X_LUT4
    generic map(
      INIT => X"2AEA"
    )
    port map (
      ADR0 => mac_control_dout(13),
      ADR1 => mac_control_n0086,
      ADR2 => mac_control_sclkdeltall,
      ADR3 => mac_control_N81479,
      O => mac_control_n0016(14)
    );
  mac_control_dout_14_XUSED : X_BUF
    port map (
      I => mac_control_dout_14_FROM,
      O => mac_control_N81479
    );
  mac_control_txfifowerr_cntl_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_25_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_17_FFY_RST
    );
  mac_control_txfifowerr_cntl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(16),
      CE => mac_control_txfifowerr_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_17_FFY_RST,
      O => mac_control_txfifowerr_cntl(16)
    );
  mac_control_txfifowerr_cntl_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_17_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_27_FFY_RST
    );
  mac_control_txfifowerr_cntl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(26),
      CE => mac_control_txfifowerr_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_27_FFY_RST,
      O => mac_control_txfifowerr_cntl(26)
    );
  mac_control_txfifowerr_cntl_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_27_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_19_FFY_RST
    );
  mac_control_txfifowerr_cntl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(18),
      CE => mac_control_txfifowerr_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_19_FFY_RST,
      O => mac_control_txfifowerr_cntl(18)
    );
  mac_control_txfifowerr_cntl_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_19_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_29_FFY_RST
    );
  mac_control_txfifowerr_cntl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(28),
      CE => mac_control_txfifowerr_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_29_FFY_RST,
      O => mac_control_txfifowerr_cntl(28)
    );
  mac_control_txfifowerr_cntl_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_29_CEMUXNOT
    );
  mac_control_dout_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_15_FFY_RST
    );
  mac_control_dout_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(15),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_15_FFY_RST,
      O => mac_control_dout(15)
    );
  mac_control_Mmux_n0016_Result_15_93_SW1 : X_LUT4
    generic map(
      INIT => X"F1F3"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_CHOICE2599,
      ADR2 => mac_control_addr(5),
      ADR3 => mac_control_phydo(15),
      O => mac_control_dout_15_FROM
    );
  mac_control_Mmux_n0016_Result_15_93 : X_LUT4
    generic map(
      INIT => X"4CEC"
    )
    port map (
      ADR0 => mac_control_sclkdeltall,
      ADR1 => mac_control_dout(14),
      ADR2 => mac_control_n0086,
      ADR3 => mac_control_N81483,
      O => mac_control_n0016(15)
    );
  mac_control_dout_15_XUSED : X_BUF
    port map (
      I => mac_control_dout_15_FROM,
      O => mac_control_N81483
    );
  tx_output_ldata_6_17 : X_LUT4
    generic map(
      INIT => X"0004"
    )
    port map (
      ADR0 => tx_output_cs_FFd5_1,
      ADR1 => q2(6),
      ADR2 => tx_output_cs_FFd6_1,
      ADR3 => tx_output_cs_FFd4_1,
      O => tx_output_CHOICE1670_FROM
    );
  tx_output_cs_Out1157_SW1 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd4_1,
      ADR1 => tx_output_cs_FFd6_1,
      ADR2 => tx_output_cs_FFd9,
      ADR3 => tx_output_cs_FFd8,
      O => tx_output_CHOICE1670_GROM
    );
  tx_output_CHOICE1670_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1670_FROM,
      O => tx_output_CHOICE1670
    );
  tx_output_CHOICE1670_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1670_GROM,
      O => tx_output_N81401
    );
  rx_input_fifo_fifo_BU279 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1529,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1543_FFX_RST,
      O => rx_input_fifo_fifo_N1543
    );
  rx_input_fifo_fifo_N1543_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1543_FFX_RST
    );
  tx_fifocheck_fbbpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_3_FFY_RST
    );
  tx_fifocheck_fbbpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_3_FFY_RST,
      O => tx_fifocheck_fbbpl(2)
    );
  tx_fifocheck_fbbpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_5_FFY_RST
    );
  tx_fifocheck_fbbpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_5_FFY_RST,
      O => tx_fifocheck_fbbpl(4)
    );
  mac_control_Mmux_n0016_Result_24_48_SW0 : X_LUT4
    generic map(
      INIT => X"FEFC"
    )
    port map (
      ADR0 => mac_control_n0067,
      ADR1 => mac_control_CHOICE2391,
      ADR2 => mac_control_n0056,
      ADR3 => mac_control_rxcrcerr_cntl(24),
      O => mac_control_N81046_FROM
    );
  mac_control_Mmux_n0016_Result_24_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2387,
      ADR1 => mac_control_CHOICE2396,
      ADR2 => mac_control_CHOICE2384,
      ADR3 => mac_control_N81046,
      O => mac_control_N81046_GROM
    );
  mac_control_N81046_XUSED : X_BUF
    port map (
      I => mac_control_N81046_FROM,
      O => mac_control_N81046
    );
  mac_control_N81046_YUSED : X_BUF
    port map (
      I => mac_control_N81046_GROM,
      O => mac_control_CHOICE2399
    );
  mac_control_Mmux_n0016_Result_16_48_SW0 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_CHOICE2319,
      ADR1 => mac_control_rxcrcerr_cntl(16),
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_n0056,
      O => mac_control_N81074_FROM
    );
  mac_control_Mmux_n0016_Result_16_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2312,
      ADR1 => mac_control_CHOICE2324,
      ADR2 => mac_control_CHOICE2315,
      ADR3 => mac_control_N81074,
      O => mac_control_N81074_GROM
    );
  mac_control_N81074_XUSED : X_BUF
    port map (
      I => mac_control_N81074_FROM,
      O => mac_control_N81074
    );
  mac_control_N81074_YUSED : X_BUF
    port map (
      I => mac_control_N81074_GROM,
      O => mac_control_CHOICE2327
    );
  tx_fifocheck_fbbpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_9_FFY_RST
    );
  tx_fifocheck_fbbpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_9_FFY_RST,
      O => tx_fifocheck_fbbpl(8)
    );
  mac_control_phydo_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_11_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(10),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_11_FFY_RST,
      O => mac_control_phydo(10)
    );
  mac_control_n00151 : X_LUT4
    generic map(
      INIT => X"3330"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => mac_control_sclkdelta,
      ADR3 => mac_control_Mshreg_scslll_103,
      O => mac_control_n0015_FROM
    );
  mac_control_n00101 : X_LUT4
    generic map(
      INIT => X"00A0"
    )
    port map (
      ADR0 => mac_control_N53154,
      ADR1 => VCC,
      ADR2 => mac_control_sclkdelta,
      ADR3 => RESET_IBUF,
      O => mac_control_n0015_GROM
    );
  mac_control_n0015_XUSED : X_BUF
    port map (
      I => mac_control_n0015_FROM,
      O => mac_control_n0015
    );
  mac_control_n0015_YUSED : X_BUF
    port map (
      I => mac_control_n0015_GROM,
      O => mac_control_n0010
    );
  tx_output_cs_Out1435_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd11,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_cs_FFd14,
      ADR3 => tx_output_cs_FFd13,
      O => tx_output_ltxen3_FROM
    );
  tx_output_cs_Out1435 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_N80959,
      ADR1 => tx_output_CHOICE1779,
      ADR2 => tx_output_CHOICE1775,
      ADR3 => tx_output_CHOICE1782,
      O => tx_output_ltxen
    );
  tx_output_ltxen3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_ltxen3_CEMUXNOT
    );
  tx_output_ltxen3_XUSED : X_BUF
    port map (
      I => tx_output_ltxen3_FROM,
      O => tx_output_N80959
    );
  mac_control_n00241 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => RESET_IBUF,
      ADR2 => mac_control_addr(7),
      ADR3 => mac_control_sclkdeltal,
      O => mac_control_n0024_FROM
    );
  mac_control_n00131 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => mac_control_addr(7),
      ADR1 => mac_control_sclkdeltal,
      ADR2 => RESET_IBUF,
      ADR3 => mac_control_n0059,
      O => mac_control_n0024_GROM
    );
  mac_control_n0024_XUSED : X_BUF
    port map (
      I => mac_control_n0024_FROM,
      O => mac_control_n0024
    );
  mac_control_n0024_YUSED : X_BUF
    port map (
      I => mac_control_n0024_GROM,
      O => mac_control_n0013
    );
  mac_control_n00251 : X_LUT4
    generic map(
      INIT => X"0008"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_N53109,
      ADR2 => mac_control_addr(2),
      ADR3 => mac_control_addr_0_1,
      O => mac_control_n0025_FROM
    );
  mac_control_n00301 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_N53109,
      ADR2 => mac_control_addr_0_1,
      ADR3 => mac_control_addr(2),
      O => mac_control_n0025_GROM
    );
  mac_control_n0025_XUSED : X_BUF
    port map (
      I => mac_control_n0025_FROM,
      O => mac_control_n0025
    );
  mac_control_n0025_YUSED : X_BUF
    port map (
      I => mac_control_n0025_GROM,
      O => mac_control_n0030
    );
  rx_input_fifo_fifo_BU342 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1530,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1557_FFY_RST,
      O => rx_input_fifo_fifo_N1558
    );
  rx_input_fifo_fifo_N1557_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1557_FFY_RST
    );
  mac_control_n00399 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_161,
      ADR1 => mac_control_ledrx_cnt_163,
      ADR2 => mac_control_ledrx_cnt_160,
      ADR3 => mac_control_ledrx_cnt_162,
      O => mac_control_CHOICE1291_FROM
    );
  mac_control_n00404 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_161,
      ADR1 => mac_control_ledrx_cnt_160,
      ADR2 => mac_control_ledrx_cnt_162,
      ADR3 => mac_control_ledrx_cnt_163,
      O => mac_control_CHOICE1291_GROM
    );
  mac_control_CHOICE1291_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1291_FROM,
      O => mac_control_CHOICE1291
    );
  mac_control_CHOICE1291_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1291_GROM,
      O => mac_control_CHOICE1266
    );
  rx_input_fifo_fifo_BU297 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N1543,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N1550_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1550
    );
  rx_input_fifo_fifo_N1550_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1550_FFX_SET
    );
  mac_control_n00291 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_N53109,
      ADR2 => mac_control_addr_0_1,
      ADR3 => mac_control_addr(2),
      O => mac_control_n0029_FROM
    );
  mac_control_n00261 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_N53109,
      ADR2 => mac_control_addr(2),
      ADR3 => mac_control_addr_0_1,
      O => mac_control_n0029_GROM
    );
  mac_control_n0029_XUSED : X_BUF
    port map (
      I => mac_control_n0029_FROM,
      O => mac_control_n0029
    );
  mac_control_n0029_YUSED : X_BUF
    port map (
      I => mac_control_n0029_GROM,
      O => mac_control_n0026
    );
  mac_control_n00327 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_123,
      ADR1 => mac_control_phyrstcnt_121,
      ADR2 => mac_control_phyrstcnt_122,
      ADR3 => mac_control_phyrstcnt_120,
      O => mac_control_CHOICE1380_FROM
    );
  mac_control_n003210 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_119,
      ADR1 => mac_control_phyrstcnt_118,
      ADR2 => mac_control_phyrstcnt_110,
      ADR3 => mac_control_CHOICE1380,
      O => mac_control_CHOICE1380_GROM
    );
  mac_control_CHOICE1380_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1380_FROM,
      O => mac_control_CHOICE1380
    );
  mac_control_CHOICE1380_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1380_GROM,
      O => mac_control_CHOICE1381
    );
  mac_control_n00601 : X_LUT4
    generic map(
      INIT => X"0020"
    )
    port map (
      ADR0 => mac_control_addr(3),
      ADR1 => mac_control_addr(2),
      ADR2 => mac_control_N53204,
      ADR3 => mac_control_addr(4),
      O => mac_control_n0060_FROM
    );
  mac_control_n00271 : X_LUT4
    generic map(
      INIT => X"0008"
    )
    port map (
      ADR0 => mac_control_N53109,
      ADR1 => mac_control_addr(2),
      ADR2 => mac_control_addr_0_1,
      ADR3 => mac_control_addr(1),
      O => mac_control_n0060_GROM
    );
  mac_control_n0060_XUSED : X_BUF
    port map (
      I => mac_control_n0060_FROM,
      O => mac_control_n0060
    );
  mac_control_n0060_YUSED : X_BUF
    port map (
      I => mac_control_n0060_GROM,
      O => mac_control_n0027
    );
  mac_control_n00361 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phystat(4),
      ADR2 => mac_control_phystat(3),
      ADR3 => VCC,
      O => mac_control_n0036_FROM
    );
  mac_control_n00351 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phystat(4),
      ADR2 => VCC,
      ADR3 => mac_control_phystat(3),
      O => mac_control_n0036_GROM
    );
  mac_control_n0036_XUSED : X_BUF
    port map (
      I => mac_control_n0036_FROM,
      O => mac_control_n0036
    );
  mac_control_n0036_YUSED : X_BUF
    port map (
      I => mac_control_n0036_GROM,
      O => mac_control_n0035
    );
  mac_control_Mmux_n0016_Result_25_45_SW0 : X_LUT4
    generic map(
      INIT => X"EAEA"
    )
    port map (
      ADR0 => mac_control_CHOICE2208,
      ADR1 => mac_control_phydi(25),
      ADR2 => mac_control_n0059,
      ADR3 => VCC,
      O => mac_control_N81098_FROM
    );
  mac_control_Mmux_n0016_Result_25_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2204,
      ADR1 => mac_control_CHOICE2200,
      ADR2 => mac_control_CHOICE2197,
      ADR3 => mac_control_N81098,
      O => mac_control_N81098_GROM
    );
  mac_control_N81098_XUSED : X_BUF
    port map (
      I => mac_control_N81098_FROM,
      O => mac_control_N81098
    );
  mac_control_N81098_YUSED : X_BUF
    port map (
      I => mac_control_N81098_GROM,
      O => mac_control_CHOICE2211
    );
  mac_control_n00374 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_147,
      ADR1 => mac_control_ledtx_cnt_144,
      ADR2 => mac_control_ledtx_cnt_146,
      ADR3 => mac_control_ledtx_cnt_145,
      O => mac_control_CHOICE1302_GROM
    );
  mac_control_CHOICE1302_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1302_GROM,
      O => mac_control_CHOICE1302
    );
  mac_control_n00631 : X_LUT4
    generic map(
      INIT => X"8800"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => mac_control_addr(1),
      ADR2 => VCC,
      ADR3 => mac_control_N53125,
      O => mac_control_n0063_FROM
    );
  mac_control_Mmux_n0016_Result_1_30 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cntl(1),
      ADR1 => mac_control_phyaddr(1),
      ADR2 => mac_control_n00851_1,
      ADR3 => mac_control_n0063,
      O => mac_control_n0063_GROM
    );
  mac_control_n0063_XUSED : X_BUF
    port map (
      I => mac_control_n0063_FROM,
      O => mac_control_n0063
    );
  mac_control_n0063_YUSED : X_BUF
    port map (
      I => mac_control_n0063_GROM,
      O => mac_control_CHOICE2620
    );
  mac_control_n00379 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_151,
      ADR1 => mac_control_ledtx_cnt_149,
      ADR2 => mac_control_ledtx_cnt_148,
      ADR3 => mac_control_ledtx_cnt_150,
      O => mac_control_CHOICE1305_FROM
    );
  mac_control_n00384 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_ledtx_cnt_151,
      ADR1 => mac_control_ledtx_cnt_148,
      ADR2 => mac_control_ledtx_cnt_149,
      ADR3 => mac_control_ledtx_cnt_150,
      O => mac_control_CHOICE1305_GROM
    );
  mac_control_CHOICE1305_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1305_FROM,
      O => mac_control_CHOICE1305
    );
  mac_control_CHOICE1305_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1305_GROM,
      O => mac_control_CHOICE1277
    );
  mac_control_Mmux_n0016_Result_31_85_SW0_SW0 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => mac_control_addr(3),
      ADR1 => mac_control_addr_0_1,
      ADR2 => mac_control_phyaddr(31),
      ADR3 => mac_control_N53132,
      O => mac_control_N81417_FROM
    );
  mac_control_n00561 : X_LUT4
    generic map(
      INIT => X"000C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N53132,
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_addr(3),
      O => mac_control_N81417_GROM
    );
  mac_control_N81417_XUSED : X_BUF
    port map (
      I => mac_control_N81417_FROM,
      O => mac_control_N81417
    );
  mac_control_N81417_YUSED : X_BUF
    port map (
      I => mac_control_N81417_GROM,
      O => mac_control_n0056
    );
  rx_input_fifo_fifo_BU344 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1529,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1557_FFX_RST,
      O => rx_input_fifo_fifo_N1557
    );
  rx_input_fifo_fifo_N1557_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1557_FFX_RST
    );
  mac_control_n00641 : X_LUT4
    generic map(
      INIT => X"0022"
    )
    port map (
      ADR0 => mac_control_N53118,
      ADR1 => mac_control_addr(0),
      ADR2 => VCC,
      ADR3 => mac_control_addr(1),
      O => mac_control_n0064_FROM
    );
  mac_control_Mmux_n0016_Result_12_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cntl(12),
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_rxfifowerr_cntl(12),
      ADR3 => mac_control_n0064,
      O => mac_control_n0064_GROM
    );
  mac_control_n0064_XUSED : X_BUF
    port map (
      I => mac_control_n0064_FROM,
      O => mac_control_n0064
    );
  mac_control_n0064_YUSED : X_BUF
    port map (
      I => mac_control_n0064_GROM,
      O => mac_control_CHOICE2536
    );
  mac_control_n00394 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_156,
      ADR1 => mac_control_ledrx_cnt_159,
      ADR2 => mac_control_ledrx_cnt_158,
      ADR3 => mac_control_ledrx_cnt_157,
      O => mac_control_CHOICE1288_GROM
    );
  mac_control_CHOICE1288_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1288_GROM,
      O => mac_control_CHOICE1288
    );
  mac_control_n00571 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => mac_control_N53204,
      ADR1 => mac_control_addr(3),
      ADR2 => mac_control_addr(2),
      ADR3 => mac_control_addr(4),
      O => mac_control_n0057_FROM
    );
  mac_control_Mmux_n0016_Result_0_82_SW0 : X_LUT4
    generic map(
      INIT => X"0777"
    )
    port map (
      ADR0 => mac_control_n0060,
      ADR1 => mac_control_phydo(0),
      ADR2 => mac_control_phystat(0),
      ADR3 => mac_control_n0057,
      O => mac_control_n0057_GROM
    );
  mac_control_n0057_XUSED : X_BUF
    port map (
      I => mac_control_n0057_FROM,
      O => mac_control_n0057
    );
  mac_control_n0057_YUSED : X_BUF
    port map (
      I => mac_control_n0057_GROM,
      O => mac_control_N81030
    );
  mac_control_n00651 : X_LUT4
    generic map(
      INIT => X"2200"
    )
    port map (
      ADR0 => mac_control_N53118,
      ADR1 => mac_control_addr(1),
      ADR2 => VCC,
      ADR3 => mac_control_addr(0),
      O => mac_control_n0065_FROM
    );
  mac_control_Mmux_n0016_Result_6_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_rxphyerr_cntl(6),
      ADR2 => mac_control_rxfifowerr_cntl(6),
      ADR3 => mac_control_n0065,
      O => mac_control_n0065_GROM
    );
  mac_control_n0065_XUSED : X_BUF
    port map (
      I => mac_control_n0065_FROM,
      O => mac_control_n0065
    );
  mac_control_n0065_YUSED : X_BUF
    port map (
      I => mac_control_n0065_GROM,
      O => mac_control_CHOICE2686
    );
  mac_control_n00661 : X_LUT4
    generic map(
      INIT => X"0080"
    )
    port map (
      ADR0 => mac_control_N53204,
      ADR1 => mac_control_addr(2),
      ADR2 => mac_control_addr(4),
      ADR3 => mac_control_addr(3),
      O => mac_control_n0066_FROM
    );
  mac_control_Mmux_n0016_Result_20_28 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0061,
      ADR1 => mac_control_rxoferr_cntl(20),
      ADR2 => mac_control_txf_cntl(20),
      ADR3 => mac_control_n0066,
      O => mac_control_n0066_GROM
    );
  mac_control_n0066_XUSED : X_BUF
    port map (
      I => mac_control_n0066_FROM,
      O => mac_control_n0066
    );
  mac_control_n0066_YUSED : X_BUF
    port map (
      I => mac_control_n0066_GROM,
      O => mac_control_CHOICE2139
    );
  mac_control_Mmux_n0016_Result_17_48_SW0 : X_LUT4
    generic map(
      INIT => X"FEFA"
    )
    port map (
      ADR0 => mac_control_CHOICE2343,
      ADR1 => mac_control_rxcrcerr_cntl(17),
      ADR2 => mac_control_n0056,
      ADR3 => mac_control_n0067,
      O => mac_control_N81070_FROM
    );
  mac_control_Mmux_n0016_Result_17_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2339,
      ADR1 => mac_control_CHOICE2336,
      ADR2 => mac_control_CHOICE2348,
      ADR3 => mac_control_N81070,
      O => mac_control_N81070_GROM
    );
  mac_control_N81070_XUSED : X_BUF
    port map (
      I => mac_control_N81070_FROM,
      O => mac_control_N81070
    );
  mac_control_N81070_YUSED : X_BUF
    port map (
      I => mac_control_N81070_GROM,
      O => mac_control_CHOICE2351
    );
  mac_control_Mmux_n0016_Result_26_45_SW0 : X_LUT4
    generic map(
      INIT => X"ECEC"
    )
    port map (
      ADR0 => mac_control_phydi(26),
      ADR1 => mac_control_CHOICE2185,
      ADR2 => mac_control_n0059,
      ADR3 => VCC,
      O => mac_control_N81154_FROM
    );
  mac_control_Mmux_n0016_Result_26_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2177,
      ADR1 => mac_control_CHOICE2181,
      ADR2 => mac_control_CHOICE2174,
      ADR3 => mac_control_N81154,
      O => mac_control_N81154_GROM
    );
  mac_control_N81154_XUSED : X_BUF
    port map (
      I => mac_control_N81154_FROM,
      O => mac_control_N81154
    );
  mac_control_N81154_YUSED : X_BUF
    port map (
      I => mac_control_N81154_GROM,
      O => mac_control_CHOICE2188
    );
  mac_control_Mmux_n0016_Result_18_45_SW0 : X_LUT4
    generic map(
      INIT => X"F8F8"
    )
    port map (
      ADR0 => mac_control_phydi(18),
      ADR1 => mac_control_n0059,
      ADR2 => mac_control_CHOICE2070,
      ADR3 => VCC,
      O => mac_control_N81130_FROM
    );
  mac_control_Mmux_n0016_Result_18_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2059,
      ADR1 => mac_control_CHOICE2066,
      ADR2 => mac_control_CHOICE2062,
      ADR3 => mac_control_N81130,
      O => mac_control_N81130_GROM
    );
  mac_control_N81130_XUSED : X_BUF
    port map (
      I => mac_control_N81130_FROM,
      O => mac_control_N81130
    );
  mac_control_N81130_YUSED : X_BUF
    port map (
      I => mac_control_N81130_GROM,
      O => mac_control_CHOICE2073
    );
  tx_output_ldata_0_26_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => q2(8),
      ADR1 => tx_output_cs_FFd4_1,
      ADR2 => tx_output_cs_FFd6_1,
      ADR3 => q2(24),
      O => tx_output_data_0_FROM
    );
  tx_output_ldata_0_26 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => q2(16),
      ADR1 => tx_output_cs_FFd5_1,
      ADR2 => tx_output_CHOICE1742,
      ADR3 => tx_output_N80998,
      O => tx_output_ldata(0)
    );
  tx_output_data_0_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_data_0_CEMUXNOT
    );
  tx_output_data_0_XUSED : X_BUF
    port map (
      I => tx_output_data_0_FROM,
      O => tx_output_N80998
    );
  mac_control_PHY_status_MII_Interface_sts28 : X_LUT4
    generic map(
      INIT => X"01BB"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR1 => mac_control_PHY_status_MII_Interface_N81159,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR3 => mac_control_PHY_status_miirw,
      O => mac_control_PHY_status_MII_Interface_CHOICE872_FROM
    );
  mac_control_PHY_status_MII_Interface_sts35 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(5),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE872,
      O => mac_control_PHY_status_MII_Interface_CHOICE872_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE872_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE872_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE872
    );
  mac_control_PHY_status_MII_Interface_CHOICE872_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE872_GROM,
      O => mac_control_PHY_status_MII_Interface_sts
    );
  mac_control_Mmux_n0016_Result_1_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cntl(1),
      ADR1 => mac_control_n0064,
      ADR2 => mac_control_n0065,
      ADR3 => mac_control_rxfifowerr_cntl(1),
      O => mac_control_CHOICE2608_FROM
    );
  mac_control_Mmux_n0016_Result_0_5 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_n0065,
      ADR2 => mac_control_rxfifowerr_cntl(0),
      ADR3 => mac_control_rxphyerr_cntl(0),
      O => mac_control_CHOICE2608_GROM
    );
  mac_control_CHOICE2608_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2608_FROM,
      O => mac_control_CHOICE2608
    );
  mac_control_CHOICE2608_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2608_GROM,
      O => mac_control_CHOICE1892
    );
  mac_control_Mmux_n0016_Result_16_22 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0062,
      ADR1 => mac_control_n0061,
      ADR2 => mac_control_rxf_cntl(16),
      ADR3 => mac_control_txf_cntl(16),
      O => mac_control_CHOICE2319_FROM
    );
  mac_control_Mmux_n0016_Result_7_5 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0067,
      ADR1 => mac_control_n0062,
      ADR2 => mac_control_rxf_cntl(7),
      ADR3 => mac_control_rxcrcerr_cntl(7),
      O => mac_control_CHOICE2319_GROM
    );
  mac_control_CHOICE2319_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2319_FROM,
      O => mac_control_CHOICE2319
    );
  mac_control_CHOICE2319_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2319_GROM,
      O => mac_control_CHOICE2458
    );
  mac_control_Mmux_n0016_Result_19_45_SW0 : X_LUT4
    generic map(
      INIT => X"FCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0059,
      ADR2 => mac_control_CHOICE2093,
      ADR3 => mac_control_phydi(19),
      O => mac_control_N81146_FROM
    );
  mac_control_Mmux_n0016_Result_19_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2089,
      ADR1 => mac_control_CHOICE2085,
      ADR2 => mac_control_CHOICE2082,
      ADR3 => mac_control_N81146,
      O => mac_control_N81146_GROM
    );
  mac_control_N81146_XUSED : X_BUF
    port map (
      I => mac_control_N81146_FROM,
      O => mac_control_N81146
    );
  mac_control_N81146_YUSED : X_BUF
    port map (
      I => mac_control_N81146_GROM,
      O => mac_control_CHOICE2096
    );
  rx_input_fifo_fifo_BU328 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N7,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1578_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1578
    );
  rx_input_fifo_fifo_N1578_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1578_FFX_SET
    );
  mac_control_Mmux_n0016_Result_27_45_SW0 : X_LUT4
    generic map(
      INIT => X"EECC"
    )
    port map (
      ADR0 => mac_control_phydi(27),
      ADR1 => mac_control_CHOICE2231,
      ADR2 => VCC,
      ADR3 => mac_control_n0059,
      O => mac_control_N81142_FROM
    );
  mac_control_Mmux_n0016_Result_27_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2223,
      ADR1 => mac_control_CHOICE2220,
      ADR2 => mac_control_CHOICE2227,
      ADR3 => mac_control_N81142,
      O => mac_control_N81142_GROM
    );
  mac_control_N81142_XUSED : X_BUF
    port map (
      I => mac_control_N81142_FROM,
      O => mac_control_N81142
    );
  mac_control_N81142_YUSED : X_BUF
    port map (
      I => mac_control_N81142_GROM,
      O => mac_control_CHOICE2234
    );
  rx_input_fifo_fifo_BU402 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3685,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1565_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1564
    );
  rx_input_fifo_fifo_N1565_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1565_FFY_SET
    );
  rx_input_memio_addrchk_cs_FFd6_In7 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd5,
      ADR1 => rx_input_memio_addrchk_cs_FFd6,
      ADR2 => rx_input_memio_addrchk_cs_FFd4,
      ADR3 => rx_input_memio_addrchk_cs_FFd3,
      O => rx_input_memio_addrchk_CHOICE1789_FROM
    );
  rx_input_memio_addrchk_n00301 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_RESET_1,
      ADR3 => rx_input_memio_addrchk_cs_FFd3,
      O => rx_input_memio_addrchk_CHOICE1789_GROM
    );
  rx_input_memio_addrchk_CHOICE1789_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1789_FROM,
      O => rx_input_memio_addrchk_CHOICE1789
    );
  rx_input_memio_addrchk_CHOICE1789_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1789_GROM,
      O => rx_input_memio_addrchk_n0030
    );
  rx_input_memio_addrchk_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"0B08"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd3,
      ADR1 => rx_input_memio_brdy,
      ADR2 => rx_input_memio_cs_FFd16_1,
      ADR3 => rx_input_memio_addrchk_cs_FFd2,
      O => rx_input_memio_addrchk_cs_FFd2_In
    );
  rx_input_memio_addrchk_n00311 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_cs_FFd2,
      ADR2 => VCC,
      ADR3 => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_cs_FFd2_GROM
    );
  rx_input_memio_addrchk_cs_FFd2_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_cs_FFd2_GROM,
      O => rx_input_memio_addrchk_n0031
    );
  tx_output_ldata_1_26_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => q2(9),
      ADR1 => tx_output_cs_FFd4_1,
      ADR2 => tx_output_cs_FFd6_1,
      ADR3 => q2(25),
      O => tx_output_data_1_FROM
    );
  tx_output_ldata_1_26 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => tx_output_cs_FFd5_1,
      ADR1 => tx_output_CHOICE1718,
      ADR2 => q2(17),
      ADR3 => tx_output_N81010,
      O => tx_output_ldata(1)
    );
  tx_output_data_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_data_1_CEMUXNOT
    );
  tx_output_data_1_XUSED : X_BUF
    port map (
      I => tx_output_data_1_FROM,
      O => tx_output_N81010
    );
  rx_input_memio_addrchk_n00414 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(18),
      ADR1 => rx_input_memio_addrchk_datal(16),
      ADR2 => rx_input_memio_addrchk_datal(17),
      ADR3 => rx_input_memio_addrchk_datal(19),
      O => rx_input_memio_addrchk_CHOICE1560_GROM
    );
  rx_input_memio_addrchk_CHOICE1560_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1560_GROM,
      O => rx_input_memio_addrchk_CHOICE1560
    );
  rx_input_memio_addrchk_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"00E2"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd5,
      ADR1 => rx_input_memio_brdy,
      ADR2 => rx_input_memio_addrchk_cs_FFd6,
      ADR3 => rx_input_memio_cs_FFd16_1,
      O => rx_input_memio_addrchk_cs_FFd5_In
    );
  rx_input_memio_addrchk_n00271 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_RESET_1,
      ADR3 => rx_input_memio_addrchk_cs_FFd6,
      O => rx_input_memio_addrchk_cs_FFd5_GROM
    );
  rx_input_memio_addrchk_cs_FFd5_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_cs_FFd5_GROM,
      O => rx_input_memio_addrchk_n0027
    );
  rx_input_memio_addrchk_n00281 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_cs_FFd5,
      ADR2 => rx_input_memio_RESET_1,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_n0028_GROM
    );
  rx_input_memio_addrchk_n0028_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_n0028_GROM,
      O => rx_input_memio_addrchk_n0028
    );
  rx_input_memio_addrchk_n00354 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(3),
      ADR1 => rx_input_memio_addrchk_datal(2),
      ADR2 => rx_input_memio_addrchk_datal(0),
      ADR3 => rx_input_memio_addrchk_datal(1),
      O => rx_input_memio_addrchk_CHOICE1567_GROM
    );
  rx_input_memio_addrchk_CHOICE1567_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1567_GROM,
      O => rx_input_memio_addrchk_CHOICE1567
    );
  rx_input_memio_addrchk_n00419 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(21),
      ADR1 => rx_input_memio_addrchk_datal(20),
      ADR2 => rx_input_memio_addrchk_datal(22),
      ADR3 => rx_input_memio_addrchk_datal(23),
      O => rx_input_memio_addrchk_bcast_3_FROM
    );
  rx_input_memio_addrchk_n004110 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_CHOICE1560,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1563,
      O => rx_input_memio_addrchk_lbcast(3)
    );
  rx_input_memio_addrchk_bcast_3_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_bcast_3_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_3_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_3_FROM,
      O => rx_input_memio_addrchk_CHOICE1563
    );
  rx_input_memio_addrchk_n00291 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd4,
      ADR1 => VCC,
      ADR2 => rx_input_memio_RESET_1,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_n0029_GROM
    );
  rx_input_memio_addrchk_n0029_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_n0029_GROM,
      O => rx_input_memio_addrchk_n0029
    );
  rx_input_memio_addrchk_n00444 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(27),
      ADR1 => rx_input_memio_addrchk_datal(26),
      ADR2 => rx_input_memio_addrchk_datal(24),
      ADR3 => rx_input_memio_addrchk_datal(25),
      O => rx_input_memio_addrchk_CHOICE1546_GROM
    );
  rx_input_memio_addrchk_CHOICE1546_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1546_GROM,
      O => rx_input_memio_addrchk_CHOICE1546
    );
  rx_input_memio_addrchk_n00509 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(44),
      ADR1 => rx_input_memio_addrchk_datal(45),
      ADR2 => rx_input_memio_addrchk_datal(46),
      ADR3 => rx_input_memio_addrchk_datal(47),
      O => rx_input_memio_addrchk_bcast_0_FROM
    );
  rx_input_memio_addrchk_n005010 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_addrchk_CHOICE1525,
      ADR3 => rx_input_memio_addrchk_CHOICE1528,
      O => rx_input_memio_addrchk_lbcast(0)
    );
  rx_input_memio_addrchk_bcast_0_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_bcast_0_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_0_FROM,
      O => rx_input_memio_addrchk_CHOICE1528
    );
  rx_input_memio_addrchk_n00359 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(4),
      ADR1 => rx_input_memio_addrchk_datal(5),
      ADR2 => rx_input_memio_addrchk_datal(7),
      ADR3 => rx_input_memio_addrchk_datal(6),
      O => rx_input_memio_addrchk_bcast_5_FROM
    );
  rx_input_memio_addrchk_n003510 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_CHOICE1567,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1570,
      O => rx_input_memio_addrchk_lbcast(5)
    );
  rx_input_memio_addrchk_bcast_5_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_bcast_5_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_5_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_5_FROM,
      O => rx_input_memio_addrchk_CHOICE1570
    );
  rx_input_memio_addrchk_n00384 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(8),
      ADR1 => rx_input_memio_addrchk_datal(9),
      ADR2 => rx_input_memio_addrchk_datal(10),
      ADR3 => rx_input_memio_addrchk_datal(11),
      O => rx_input_memio_addrchk_CHOICE1574_GROM
    );
  rx_input_memio_addrchk_CHOICE1574_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1574_GROM,
      O => rx_input_memio_addrchk_CHOICE1574
    );
  rx_input_memio_addrchk_n00449 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(29),
      ADR1 => rx_input_memio_addrchk_datal(28),
      ADR2 => rx_input_memio_addrchk_datal(31),
      ADR3 => rx_input_memio_addrchk_datal(30),
      O => rx_input_memio_addrchk_bcast_2_FROM
    );
  rx_input_memio_addrchk_n004410 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_addrchk_CHOICE1546,
      ADR3 => rx_input_memio_addrchk_CHOICE1549,
      O => rx_input_memio_addrchk_lbcast(2)
    );
  rx_input_memio_addrchk_bcast_2_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_bcast_2_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_2_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_2_FROM,
      O => rx_input_memio_addrchk_CHOICE1549
    );
  rx_input_memio_addrchk_n00474 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(32),
      ADR1 => rx_input_memio_addrchk_datal(33),
      ADR2 => rx_input_memio_addrchk_datal(35),
      ADR3 => rx_input_memio_addrchk_datal(34),
      O => rx_input_memio_addrchk_CHOICE1553_GROM
    );
  rx_input_memio_addrchk_CHOICE1553_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_CHOICE1553_GROM,
      O => rx_input_memio_addrchk_CHOICE1553
    );
  rx_input_memio_addrchk_n00389 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(14),
      ADR1 => rx_input_memio_addrchk_datal(15),
      ADR2 => rx_input_memio_addrchk_datal(12),
      ADR3 => rx_input_memio_addrchk_datal(13),
      O => rx_input_memio_addrchk_bcast_4_FROM
    );
  rx_input_memio_addrchk_n003810 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_CHOICE1574,
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_CHOICE1577,
      O => rx_input_memio_addrchk_lbcast(4)
    );
  rx_input_memio_addrchk_bcast_4_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_bcast_4_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_4_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_4_FROM,
      O => rx_input_memio_addrchk_CHOICE1577
    );
  rx_input_memio_addrchk_n00479 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(38),
      ADR1 => rx_input_memio_addrchk_datal(39),
      ADR2 => rx_input_memio_addrchk_datal(37),
      ADR3 => rx_input_memio_addrchk_datal(36),
      O => rx_input_memio_addrchk_bcast_1_FROM
    );
  rx_input_memio_addrchk_n004710 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_addrchk_CHOICE1553,
      ADR3 => rx_input_memio_addrchk_CHOICE1556,
      O => rx_input_memio_addrchk_lbcast(1)
    );
  rx_input_memio_addrchk_bcast_1_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_bcast_1_CEMUXNOT
    );
  rx_input_memio_addrchk_bcast_1_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_bcast_1_FROM,
      O => rx_input_memio_addrchk_CHOICE1556
    );
  mac_control_n0012_SW0 : X_LUT4
    generic map(
      INIT => X"FBFB"
    )
    port map (
      ADR0 => mac_control_N53154,
      ADR1 => mac_control_sclkdelta,
      ADR2 => mac_control_addr(7),
      ADR3 => VCC,
      O => mac_control_N69607_FROM
    );
  mac_control_n0012_53 : X_LUT4
    generic map(
      INIT => X"2033"
    )
    port map (
      ADR0 => mac_control_n0086,
      ADR1 => RESET_IBUF,
      ADR2 => mac_control_sclkdeltall,
      ADR3 => mac_control_N69607,
      O => mac_control_N69607_GROM
    );
  mac_control_N69607_XUSED : X_BUF
    port map (
      I => mac_control_N69607_FROM,
      O => mac_control_N69607
    );
  mac_control_N69607_YUSED : X_BUF
    port map (
      I => mac_control_N69607_GROM,
      O => mac_control_n0012
    );
  mac_control_Ker53142_SW0 : X_LUT4
    generic map(
      INIT => X"3FFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_sclkdeltal,
      ADR2 => mac_control_addr(7),
      ADR3 => mac_control_din(0),
      O => mac_control_N69759_FROM
    );
  mac_control_Ker53107_SW0 : X_LUT4
    generic map(
      INIT => X"CCFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => mac_control_addr(7),
      O => mac_control_N69759_GROM
    );
  mac_control_N69759_XUSED : X_BUF
    port map (
      I => mac_control_N69759_FROM,
      O => mac_control_N69759
    );
  mac_control_N69759_YUSED : X_BUF
    port map (
      I => mac_control_N69759_GROM,
      O => mac_control_N69572
    );
  mac_control_n0014_SW0 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => mac_control_addr_0_1,
      ADR1 => mac_control_addr(3),
      ADR2 => mac_control_sclkdeltal,
      ADR3 => mac_control_addr(7),
      O => mac_control_N72031_FROM
    );
  mac_control_n0014_54 : X_LUT4
    generic map(
      INIT => X"0400"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_addr(4),
      ADR2 => mac_control_addr(2),
      ADR3 => mac_control_N72031,
      O => mac_control_N72031_GROM
    );
  mac_control_N72031_XUSED : X_BUF
    port map (
      I => mac_control_N72031_FROM,
      O => mac_control_N72031
    );
  mac_control_N72031_YUSED : X_BUF
    port map (
      I => mac_control_N72031_GROM,
      O => mac_control_n0014
    );
  tx_output_cs_FFd12_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd12_FFY_RST
    );
  tx_output_cs_FFd11_55 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd12,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd12_FFY_RST,
      O => tx_output_cs_FFd11
    );
  mac_control_Mmux_n0016_Result_28_45_SW0 : X_LUT4
    generic map(
      INIT => X"EEAA"
    )
    port map (
      ADR0 => mac_control_CHOICE2254,
      ADR1 => mac_control_n0059,
      ADR2 => VCC,
      ADR3 => mac_control_phydi(28),
      O => mac_control_N81086_FROM
    );
  mac_control_Mmux_n0016_Result_28_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2250,
      ADR1 => mac_control_CHOICE2246,
      ADR2 => mac_control_CHOICE2243,
      ADR3 => mac_control_N81086,
      O => mac_control_N81086_GROM
    );
  mac_control_N81086_XUSED : X_BUF
    port map (
      I => mac_control_N81086_FROM,
      O => mac_control_N81086
    );
  mac_control_N81086_YUSED : X_BUF
    port map (
      I => mac_control_N81086_GROM,
      O => mac_control_CHOICE2257
    );
  tx_output_ldata_2_26_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => q2(10),
      ADR1 => tx_output_cs_FFd6_1,
      ADR2 => tx_output_cs_FFd4_1,
      ADR3 => q2(26),
      O => tx_output_data_2_FROM
    );
  tx_output_ldata_2_26 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => tx_output_CHOICE1730,
      ADR1 => q2(18),
      ADR2 => tx_output_cs_FFd5_1,
      ADR3 => tx_output_N81022,
      O => tx_output_ldata(2)
    );
  tx_output_data_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_data_2_CEMUXNOT
    );
  tx_output_data_2_XUSED : X_BUF
    port map (
      I => tx_output_data_2_FROM,
      O => tx_output_N81022
    );
  mac_control_Mmux_n0016_Result_29_45_SW0 : X_LUT4
    generic map(
      INIT => X"FCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_CHOICE2277,
      ADR2 => mac_control_phydi(29),
      ADR3 => mac_control_n0059,
      O => mac_control_N81126_FROM
    );
  mac_control_Mmux_n0016_Result_29_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2266,
      ADR1 => mac_control_CHOICE2269,
      ADR2 => mac_control_CHOICE2273,
      ADR3 => mac_control_N81126,
      O => mac_control_N81126_GROM
    );
  mac_control_N81126_XUSED : X_BUF
    port map (
      I => mac_control_N81126_FROM,
      O => mac_control_N81126
    );
  mac_control_N81126_YUSED : X_BUF
    port map (
      I => mac_control_N81126_GROM,
      O => mac_control_CHOICE2280
    );
  rx_input_fifo_fifo_BU400 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N3684,
      CE => VCC,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1565_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1565
    );
  rx_input_fifo_fifo_N1565_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1565_FFX_SET
    );
  tx_output_ldata_3_26_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => tx_output_cs_FFd4_1,
      ADR1 => q2(27),
      ADR2 => tx_output_cs_FFd6_1,
      ADR3 => q2(11),
      O => tx_output_data_3_FROM
    );
  tx_output_ldata_3_26 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => tx_output_cs_FFd5_1,
      ADR1 => tx_output_CHOICE1706,
      ADR2 => q2(19),
      ADR3 => tx_output_N81002,
      O => tx_output_ldata(3)
    );
  tx_output_data_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_data_3_CEMUXNOT
    );
  tx_output_data_3_XUSED : X_BUF
    port map (
      I => tx_output_data_3_FROM,
      O => tx_output_N81002
    );
  rx_input_memio_addrchk_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"5450"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16_1,
      ADR1 => rx_input_memio_addrchk_cs_FFd1,
      ADR2 => rx_input_memio_addrchk_cs_FFd7,
      ADR3 => rx_input_memio_brdy,
      O => rx_input_memio_addrchk_cs_FFd7_In
    );
  rx_input_memio_n01011 : X_LUT4
    generic map(
      INIT => X"BBAA"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16_1,
      ADR1 => rx_input_memio_menl,
      ADR2 => VCC,
      ADR3 => rx_input_memio_men,
      O => rx_input_memio_addrchk_cs_FFd7_GROM
    );
  rx_input_memio_addrchk_cs_FFd7_YUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_cs_FFd7_GROM,
      O => rx_input_memio_n0101
    );
  rx_input_memio_cs_Out917_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd1,
      ADR1 => rx_input_memio_cs_FFd3,
      ADR2 => rx_input_memio_cs_FFd2,
      ADR3 => rx_input_memio_cs_FFd5,
      O => rx_input_memio_N80990_FROM
    );
  rx_input_memio_n00301 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_memio_RESET_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd2,
      O => rx_input_memio_N80990_GROM
    );
  rx_input_memio_N80990_XUSED : X_BUF
    port map (
      I => rx_input_memio_N80990_FROM,
      O => rx_input_memio_N80990
    );
  rx_input_memio_N80990_YUSED : X_BUF
    port map (
      I => rx_input_memio_N80990_GROM,
      O => rx_input_memio_n0030
    );
  rx_input_memio_n00311 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bpen,
      ADR2 => VCC,
      ADR3 => rx_input_memio_RESET_1,
      O => rx_input_memio_n0031_GROM
    );
  rx_input_memio_n0031_YUSED : X_BUF
    port map (
      I => rx_input_memio_n0031_GROM,
      O => rx_input_memio_n0031
    );
  rx_input_memio_cs_FFd16_In1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_invalid,
      ADR2 => VCC,
      ADR3 => rx_input_endf,
      O => rx_input_memio_CHOICE1113_FROM
    );
  rx_input_memio_n00321 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_endf,
      ADR3 => rx_input_memio_RESET_1,
      O => rx_input_memio_CHOICE1113_GROM
    );
  rx_input_memio_CHOICE1113_XUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1113_FROM,
      O => rx_input_memio_CHOICE1113
    );
  rx_input_memio_CHOICE1113_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1113_GROM,
      O => rx_input_memio_n0032
    );
  rx_input_memio_n00167 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => rx_input_data(4),
      ADR1 => rx_input_data(7),
      ADR2 => rx_input_data(5),
      ADR3 => rx_input_data(6),
      O => rx_input_memio_CHOICE1979_GROM
    );
  rx_input_memio_CHOICE1979_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1979_GROM,
      O => rx_input_memio_CHOICE1979
    );
  rx_input_memio_cs_Out8_SW0 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd10,
      ADR3 => rx_input_memio_cs_FFd15,
      O => rx_input_memio_N70855_FROM
    );
  rx_input_memio_n00441 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_memio_RESET_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd15,
      O => rx_input_memio_N70855_GROM
    );
  rx_input_memio_N70855_XUSED : X_BUF
    port map (
      I => rx_input_memio_N70855_FROM,
      O => rx_input_memio_N70855
    );
  rx_input_memio_N70855_YUSED : X_BUF
    port map (
      I => rx_input_memio_N70855_GROM,
      O => rx_input_memio_n0044
    );
  rx_input_memio_n00451 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd14,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_RESET_1,
      O => rx_input_memio_n0045_GROM
    );
  rx_input_memio_n0045_YUSED : X_BUF
    port map (
      I => rx_input_memio_n0045_GROM,
      O => rx_input_memio_n0045
    );
  rx_input_fifo_fifo_BU30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1794,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_dout_9_FFY_RST,
      O => rx_input_fifo_dout(9)
    );
  rx_input_fifo_dout_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_dout_9_FFY_RST
    );
  rx_input_memio_n00461 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_memio_RESET_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd12,
      O => rx_input_memio_n0046_GROM
    );
  rx_input_memio_n0046_YUSED : X_BUF
    port map (
      I => rx_input_memio_n0046_GROM,
      O => rx_input_memio_n0046
    );
  rx_input_memio_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"AAEA"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd9,
      ADR1 => rx_input_endf,
      ADR2 => rx_input_memio_cs_FFd10,
      ADR3 => rx_input_invalid,
      O => rx_input_memio_cs_FFd8_In
    );
  rx_input_memio_n00471 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => rx_input_memio_RESET_1,
      ADR1 => rx_input_memio_cs_FFd10,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_cs_FFd8_GROM
    );
  rx_input_memio_cs_FFd8_YUSED : X_BUF
    port map (
      I => rx_input_memio_cs_FFd8_GROM,
      O => rx_input_memio_n0047
    );
  rx_input_memio_n00597 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => rx_input_memio_crcll(2),
      ADR1 => rx_input_memio_crcll(0),
      ADR2 => rx_input_memio_crcll(1),
      ADR3 => rx_input_memio_crcll(3),
      O => rx_input_memio_CHOICE1808_GROM
    );
  rx_input_memio_CHOICE1808_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1808_GROM,
      O => rx_input_memio_CHOICE1808
    );
  mac_control_bitcnt_inst_sum_256_56 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_109_CYINIT,
      I1 => mac_control_bitcnt_inst_lut3_191,
      O => mac_control_bitcnt_inst_sum_256
    );
  mac_control_bitcnt_inst_lut3_1911 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => mac_control_Mshreg_scslll_103,
      ADR1 => mac_control_bitcnt_109,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_bitcnt_inst_lut3_191
    );
  mac_control_n0086_SW0 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => mac_control_bitcnt_108,
      ADR1 => VCC,
      ADR2 => mac_control_bitcnt_105,
      ADR3 => mac_control_bitcnt_109,
      O => mac_control_bitcnt_109_GROM
    );
  mac_control_bitcnt_109_YUSED : X_BUF
    port map (
      I => mac_control_bitcnt_109_GROM,
      O => mac_control_N69675
    );
  mac_control_bitcnt_109_CYINIT_57 : X_BUF
    port map (
      I => mac_control_bitcnt_inst_cy_292,
      O => mac_control_bitcnt_109_CYINIT
    );
  tx_output_ldata_4_26_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => tx_output_cs_FFd6_1,
      ADR1 => q2(12),
      ADR2 => tx_output_cs_FFd4_1,
      ADR3 => q2(28),
      O => tx_output_data_4_FROM
    );
  tx_output_ldata_4_26 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => tx_output_cs_FFd5_1,
      ADR1 => tx_output_CHOICE1682,
      ADR2 => q2(20),
      ADR3 => tx_output_N81026,
      O => tx_output_ldata(4)
    );
  tx_output_data_4_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_data_4_CEMUXNOT
    );
  tx_output_data_4_XUSED : X_BUF
    port map (
      I => tx_output_data_4_FROM,
      O => tx_output_N81026
    );
  tx_output_bcntl_12_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bcntl_12_CEMUXNOT
    );
  tx_output_bcntl_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_14_FFY_RST
    );
  tx_output_bcntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_51,
      CE => tx_output_bcntl_14_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_14_FFY_RST,
      O => tx_output_bcntl(13)
    );
  tx_output_bcntl_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_14_FFX_RST
    );
  tx_output_bcntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_52,
      CE => tx_output_bcntl_14_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_14_FFX_RST,
      O => tx_output_bcntl(14)
    );
  tx_output_bcntl_14_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bcntl_14_CEMUXNOT
    );
  tx_output_bcntl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_15_FFY_RST
    );
  tx_output_bcntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_53,
      CE => tx_output_bcntl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_15_FFY_RST,
      O => tx_output_bcntl(15)
    );
  tx_output_bcntl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bcntl_15_CEMUXNOT
    );
  rxfbbp_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_11_FFX_RST
    );
  rx_output_bpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(11),
      CE => rxfbbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_11_FFX_RST,
      O => rxfbbp(11)
    );
  rxfbbp_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_11_FFY_RST
    );
  rx_output_bpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(10),
      CE => rxfbbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_11_FFY_RST,
      O => rxfbbp(10)
    );
  rxfbbp_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_11_CEMUXNOT
    );
  rxfbbp_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_13_FFY_RST
    );
  rx_output_bpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(12),
      CE => rxfbbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_13_FFY_RST,
      O => rxfbbp(12)
    );
  rxfbbp_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_13_FFX_RST
    );
  rx_output_bpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(13),
      CE => rxfbbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_13_FFX_RST,
      O => rxfbbp(13)
    );
  rxfbbp_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_13_CEMUXNOT
    );
  mac_control_Mshreg_scslll_srl_17 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_27,
      A1 => GLOBAL_LOGIC0_40,
      A2 => GLOBAL_LOGIC0_40,
      A3 => GLOBAL_LOGIC0_40,
      D => SCS_IBUF,
      CE => mac_control_Mshreg_scslll_net187_SRMUX_OUTPUTNOT,
      CLK => mac_control_CLKSL_4,
      Q => mac_control_Mshreg_scslll_net187_GSHIFT
    );
  mac_control_Mshreg_scslll_net187_YUSED : X_BUF
    port map (
      I => mac_control_Mshreg_scslll_net187_GSHIFT,
      O => mac_control_Mshreg_scslll_net187
    );
  mac_control_Mshreg_scslll_net187_SRMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_Mshreg_scslll_net187_SRMUX_OUTPUTNOT
    );
  rxfbbp_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_15_FFX_RST
    );
  rx_output_bpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(15),
      CE => rxfbbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_15_FFX_RST,
      O => rxfbbp(15)
    );
  rxfbbp_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_15_FFY_RST
    );
  rx_output_bpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(14),
      CE => rxfbbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_15_FFY_RST,
      O => rxfbbp(14)
    );
  rxfbbp_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_15_CEMUXNOT
    );
  rx_output_fifo_N1546_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1546_FFY_RST
    );
  rx_output_fifo_BU133 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2499,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1546_FFY_RST,
      O => rx_output_fifo_N1547
    );
  rx_output_fifo_N1546_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1546_FFX_SET
    );
  rx_output_fifo_BU140 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N10,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1546_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1546
    );
  rx_output_fifo_BU132 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N10,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N11,
      O => rx_output_fifo_N2499
    );
  rx_input_fifo_fifo_BU160 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2450,
      CE => rx_input_fifo_fifo_N2449,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_empty_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_empty
    );
  rx_input_fifo_fifo_empty_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_empty_FFY_SET
    );
  rx_output_fifo_N1610_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1610_FFY_RST
    );
  rx_output_fifo_BU294 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3427,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1610_FFY_RST,
      O => rx_output_fifo_N1611
    );
  rx_output_fifo_BU293 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_fifo_N3,
      ADR1 => rx_output_fifo_N2,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N3427
    );
  rx_output_fifo_N1563_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1563_FFY_SET
    );
  rx_output_fifo_BU320 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1546,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1563_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1562
    );
  rx_output_fifo_N1567_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1567_FFY_RST
    );
  rx_output_fifo_BU312 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1550,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1567_FFY_RST,
      O => rx_output_fifo_N1566
    );
  rx_output_fifo_BU22 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rx_output_denll,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N18_FROM
    );
  rx_output_fifo_BU144 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_output_denll,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N18_GROM
    );
  rx_output_fifo_N18_XUSED : X_BUF
    port map (
      I => rx_output_fifo_N18_FROM,
      O => rx_output_fifo_N18
    );
  rx_output_fifo_N18_YUSED : X_BUF
    port map (
      I => rx_output_fifo_N18_GROM,
      O => rx_output_fifo_N2579
    );
  rx_output_fifo_BU191 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_output_fifo_full_0,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_ceinll,
      O => rx_output_fifo_N19_FROM
    );
  rx_output_fifo_BU323 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_full_0,
      ADR2 => rx_output_ceinll,
      ADR3 => VCC,
      O => rx_output_fifo_N19_GROM
    );
  rx_output_fifo_N19_XUSED : X_BUF
    port map (
      I => rx_output_fifo_N19_FROM,
      O => rx_output_fifo_N19
    );
  rx_output_fifo_N19_YUSED : X_BUF
    port map (
      I => rx_output_fifo_N19_GROM,
      O => rx_output_fifo_N3617
    );
  rx_output_fifo_N1565_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1565_FFY_RST
    );
  rx_output_fifo_BU316 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1548,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1565_FFY_RST,
      O => rx_output_fifo_N1564
    );
  rx_input_fifo_fifo_BU127 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N2412,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_fifo_N1524_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1524
    );
  rx_input_fifo_fifo_N1524_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1524_FFY_SET
    );
  rx_output_fifo_N1569_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1569_FFX_SET
    );
  rx_output_fifo_BU306 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1553,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1569_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1569
    );
  rx_output_fifo_N1629_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1629_FFY_RST
    );
  rx_output_fifo_BU164 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1612,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1629_FFY_RST,
      O => rx_output_fifo_N1628
    );
  rx_output_fifo_N1629_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1629_FFX_RST
    );
  rx_output_fifo_BU161 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1613,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1629_FFX_RST,
      O => rx_output_fifo_N1629
    );
  rx_output_fifo_N1633_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1633_FFY_RST
    );
  rx_output_fifo_BU149 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1616,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1633_FFY_RST,
      O => rx_output_fifo_N1632
    );
  rx_output_fifo_N1633_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1633_FFX_SET
    );
  rx_output_fifo_BU146 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1617,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1633_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1633
    );
  q2_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_21_FFY_RST
    );
  memcontroller_Q2_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(20),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_21_FFY_RST,
      O => q2(20)
    );
  q2_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_21_FFX_RST
    );
  memcontroller_Q2_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(21),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_21_FFX_RST,
      O => q2(21)
    );
  q2_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_13_FFY_RST
    );
  memcontroller_Q2_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(12),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_13_FFY_RST,
      O => q2(12)
    );
  q2_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_13_FFX_RST
    );
  memcontroller_Q2_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(13),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_13_FFX_RST,
      O => q2(13)
    );
  rx_output_fifo_N1631_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1631_FFY_RST
    );
  rx_output_fifo_BU158 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1614,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1631_FFY_RST,
      O => rx_output_fifo_N1630
    );
  rx_output_fifo_N1631_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1631_FFX_RST
    );
  rx_output_fifo_BU155 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1615,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1631_FFX_RST,
      O => rx_output_fifo_N1631
    );
  rx_output_fifo_N1573_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1573_FFY_RST
    );
  rx_output_fifo_BU343 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1564,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1573_FFY_RST,
      O => rx_output_fifo_N1572
    );
  rx_output_fifo_N1573_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1573_FFX_RST
    );
  rx_output_fifo_BU340 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1565,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1573_FFX_RST,
      O => rx_output_fifo_N1573
    );
  q2_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_31_FFY_RST
    );
  memcontroller_Q2_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(30),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_31_FFY_RST,
      O => q2(30)
    );
  q2_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_31_FFX_RST
    );
  memcontroller_Q2_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(31),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_31_FFX_RST,
      O => q2(31)
    );
  q2_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_22_FFY_RST
    );
  memcontroller_Q2_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(22),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_22_FFY_RST,
      O => q2(22)
    );
  q2_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_15_FFY_RST
    );
  memcontroller_Q2_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(14),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_15_FFY_RST,
      O => q2(14)
    );
  q2_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_15_FFX_RST
    );
  memcontroller_Q2_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(15),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_15_FFX_RST,
      O => q2(15)
    );
  rx_output_fifo_N1577_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1577_FFY_SET
    );
  rx_output_fifo_BU328 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1568,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1577_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1576
    );
  rx_output_fifo_N1577_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1577_FFX_SET
    );
  rx_output_fifo_BU325 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1569,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1577_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1577
    );
  q2_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_23_FFY_RST
    );
  memcontroller_Q2_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(23),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_23_FFY_RST,
      O => q2(23)
    );
  mac_control_phystat_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_11_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(10),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_11_FFY_RST,
      O => mac_control_phystat(10)
    );
  mac_control_phystat_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_11_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(11),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_11_FFX_RST,
      O => mac_control_phystat(11)
    );
  rx_output_fifo_N1575_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1575_FFY_RST
    );
  rx_output_fifo_BU337 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1566,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1575_FFY_RST,
      O => rx_output_fifo_N1574
    );
  rx_output_fifo_N1575_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1575_FFX_RST
    );
  rx_output_fifo_BU334 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1567,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1575_FFX_RST,
      O => rx_output_fifo_N1575
    );
  rx_output_fifo_BU185 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_full_0,
      ADR2 => rx_output_ceinll,
      ADR3 => VCC,
      O => rx_output_fifo_N1517_GROM
    );
  rx_output_fifo_N1517_YUSED : X_BUF
    port map (
      I => rx_output_fifo_N1517_GROM,
      O => rx_output_fifo_N1517
    );
  q2_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_25_FFX_RST
    );
  memcontroller_Q2_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(25),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_25_FFX_RST,
      O => q2(25)
    );
  q2_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_25_FFY_RST
    );
  memcontroller_Q2_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(24),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_25_FFY_RST,
      O => q2(24)
    );
  q2_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_17_FFY_RST
    );
  memcontroller_Q2_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(16),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_17_FFY_RST,
      O => q2(16)
    );
  q2_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_17_FFX_RST
    );
  memcontroller_Q2_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(17),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_17_FFX_RST,
      O => q2(17)
    );
  rx_output_cs_FFd3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd3_FFY_RST
    );
  rx_output_cs_FFd3_58 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd3_FFY_RST,
      O => rx_output_cs_FFd3
    );
  memcontroller_n00101 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum(1),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(0),
      O => rx_output_cs_FFd3_FROM
    );
  rx_output_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => rx_output_fifo_nearfull,
      ADR1 => rx_output_cs_FFd6,
      ADR2 => rx_output_nf,
      ADR3 => clken3,
      O => rx_output_cs_FFd3_In
    );
  rx_output_cs_FFd3_XUSED : X_BUF
    port map (
      I => rx_output_cs_FFd3_FROM,
      O => clken3
    );
  rx_output_fifo_N1605_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1605_FFY_SET
    );
  rx_output_fifo_BU370 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N4,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1605_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1604
    );
  rx_output_fifo_N1609_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1609_FFY_SET
    );
  rx_output_fifo_BU362 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N8,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1609_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1608
    );
  mac_control_phystat_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_21_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(4),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_21_FFY_RST,
      O => mac_control_phystat(20)
    );
  mac_control_phystat_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_13_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(12),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_13_FFY_RST,
      O => mac_control_phystat(12)
    );
  rx_input_fifo_fifo_BU76 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1863,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N9_FFX_RST,
      O => rx_input_fifo_fifo_N9
    );
  rx_input_fifo_fifo_N9_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N9_FFX_RST
    );
  q2_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_27_FFY_RST
    );
  memcontroller_Q2_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(26),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_27_FFY_RST,
      O => q2(26)
    );
  rx_input_fifo_fifo_BU113 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2332,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1525_FFY_RST,
      O => rx_input_fifo_fifo_N1526
    );
  rx_input_fifo_fifo_N1525_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1525_FFY_RST
    );
  q2_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_19_FFY_RST
    );
  memcontroller_Q2_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(18),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_19_FFY_RST,
      O => q2(18)
    );
  q3_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_11_FFY_RST
    );
  memcontroller_Q3_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(10),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_11_FFY_RST,
      O => q3(10)
    );
  rx_output_fifo_N1585_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1585_FFY_RST
    );
  rx_output_fifo_BU380 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1552,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1585_FFY_RST,
      O => rx_output_fifo_N1584
    );
  mac_control_phystat_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_23_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(6),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_23_FFY_RST,
      O => mac_control_phystat(22)
    );
  mac_control_phystat_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_31_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(14),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_31_FFY_RST,
      O => mac_control_phystat(30)
    );
  mac_control_phystat_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_15_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(14),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_15_FFY_RST,
      O => mac_control_phystat(14)
    );
  rx_output_fifo_N1571_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1571_FFY_SET
    );
  rx_output_fifo_BU349 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1562,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => rx_output_fifo_N1571_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1570
    );
  q2_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_29_FFY_RST
    );
  memcontroller_Q2_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(28),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_29_FFY_RST,
      O => q2(28)
    );
  q3_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_21_FFY_RST
    );
  memcontroller_Q3_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(20),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_21_FFY_RST,
      O => q3(20)
    );
  q3_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_13_FFY_RST
    );
  memcontroller_Q3_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(12),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_13_FFY_RST,
      O => q3(12)
    );
  rx_output_fifo_N1586_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1586_FFY_SET
    );
  rx_output_fifo_BU468 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3974,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1586_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1587
    );
  rx_output_fifo_BU410 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N1579,
      ADR2 => rx_output_fifo_N1578,
      ADR3 => VCC,
      O => rx_output_fifo_N3974
    );
  rx_output_fifo_N1591_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1591_FFX_SET
    );
  rx_output_fifo_BU460 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3970,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1591_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1591
    );
  rx_output_fifo_BU434 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => rx_output_fifo_N3959,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N1582,
      ADR3 => rx_output_fifo_N1583,
      O => rx_output_fifo_N3970
    );
  rx_output_fifo_BU446 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_output_fifo_N1584,
      ADR1 => rx_output_fifo_N1585,
      ADR2 => rx_output_fifo_N1582,
      ADR3 => rx_output_fifo_N1583,
      O => rx_output_fifo_N1591_GROM
    );
  rx_output_fifo_N1591_YUSED : X_BUF
    port map (
      I => rx_output_fifo_N1591_GROM,
      O => rx_output_fifo_N3958
    );
  rx_output_fifo_N1603_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1603_FFY_SET
    );
  rx_output_fifo_BU374 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N2,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1603_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1602
    );
  rx_output_fifo_N1607_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1607_FFY_SET
    );
  rx_output_fifo_BU366 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N6,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1607_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1606
    );
  mac_control_phystat_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_25_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(8),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_25_FFY_RST,
      O => mac_control_phystat(24)
    );
  mac_control_phystat_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_17_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(0),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_17_FFY_RST,
      O => mac_control_phystat(16)
    );
  rx_input_fifo_fifo_BU151 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1581,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1594_FFY_RST,
      O => rx_input_fifo_fifo_N1595
    );
  rx_input_fifo_fifo_N1594_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1594_FFY_RST
    );
  q3_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_31_FFY_RST
    );
  memcontroller_Q3_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(30),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_31_FFY_RST,
      O => q3(30)
    );
  q3_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_22_FFY_RST
    );
  memcontroller_Q3_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(22),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_22_FFY_RST,
      O => q3(22)
    );
  memcontroller_n00061 : X_LUT4
    generic map(
      INIT => X"0050"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum(1),
      ADR3 => memcontroller_clknum(0),
      O => memcontroller_n0006_FROM
    );
  memcontroller_n00051 : X_LUT4
    generic map(
      INIT => X"0022"
    )
    port map (
      ADR0 => memcontroller_clknum(0),
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum(1),
      O => memcontroller_n0006_GROM
    );
  memcontroller_n0006_XUSED : X_BUF
    port map (
      I => memcontroller_n0006_FROM,
      O => memcontroller_n0006
    );
  memcontroller_n0006_YUSED : X_BUF
    port map (
      I => memcontroller_n0006_GROM,
      O => memcontroller_n0005
    );
  mac_control_phystat_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_19_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(2),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_19_FFY_RST,
      O => mac_control_phystat(18)
    );
  q3_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_25_FFY_RST
    );
  memcontroller_Q3_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(24),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_25_FFY_RST,
      O => q3(24)
    );
  q3_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_17_FFY_RST
    );
  memcontroller_Q3_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(16),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_17_FFY_RST,
      O => q3(16)
    );
  mac_control_phystat_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_29_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(12),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_29_FFY_RST,
      O => mac_control_phystat(28)
    );
  q3_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_27_FFY_RST
    );
  memcontroller_Q3_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(26),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_27_FFY_RST,
      O => q3(26)
    );
  q3_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_19_FFY_RST
    );
  memcontroller_Q3_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(18),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_19_FFY_RST,
      O => q3(18)
    );
  rx_output_fifo_N1581_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1581_FFY_RST
    );
  rx_output_fifo_BU388 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1548,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1581_FFY_RST,
      O => rx_output_fifo_N1580
    );
  q3_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_29_FFY_RST
    );
  memcontroller_Q3_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(28),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_29_FFY_RST,
      O => q3(28)
    );
  tx_output_cs_FFd17_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF_2,
      O => tx_output_cs_FFd17_FFY_SET
    );
  tx_output_cs_FFd17_59 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => tx_output_cs_FFd17_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => tx_output_cs_FFd17_FFY_SET,
      RST => GND,
      O => tx_output_cs_FFd17
    );
  memcontroller_n00091 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_0_1,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_1,
      O => tx_output_cs_FFd17_FROM
    );
  tx_output_cs_FFd17_In1 : X_LUT4
    generic map(
      INIT => X"EAFA"
    )
    port map (
      ADR0 => tx_output_cs_FFd1,
      ADR1 => tx_output_n0006,
      ADR2 => tx_output_cs_FFd17,
      ADR3 => clken2,
      O => tx_output_cs_FFd17_In
    );
  tx_output_cs_FFd17_XUSED : X_BUF
    port map (
      I => tx_output_cs_FFd17_FROM,
      O => clken2
    );
  rx_output_ceinll_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_ceinll_CEMUXNOT
    );
  tx_output_ldata_5_26_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => q2(29),
      ADR1 => q2(13),
      ADR2 => tx_output_cs_FFd4_1,
      ADR3 => tx_output_cs_FFd6_1,
      O => tx_output_data_5_FROM
    );
  tx_output_ldata_5_26 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => q2(21),
      ADR1 => tx_output_CHOICE1694,
      ADR2 => tx_output_cs_FFd5_1,
      ADR3 => tx_output_N81006,
      O => tx_output_ldata(5)
    );
  tx_output_data_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_data_5_CEMUXNOT
    );
  tx_output_data_5_XUSED : X_BUF
    port map (
      I => tx_output_data_5_FROM,
      O => tx_output_N81006
    );
  rx_input_fifo_fifo_BU71 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1862,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N11_FFY_RST,
      O => rx_input_fifo_fifo_N10
    );
  rx_input_fifo_fifo_N11_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N11_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd3_In_SW0 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => MDC_OBUF,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd4,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_cs_FFd3_FROM
    );
  mac_control_PHY_status_MII_Interface_cs_FFd3_In_60 : X_LUT4
    generic map(
      INIT => X"50DC"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_mdccnt_37,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd3,
      ADR2 => mac_control_PHY_status_MII_Interface_N70564,
      ADR3 => mac_control_PHY_status_MII_Interface_n0004,
      O => mac_control_PHY_status_MII_Interface_cs_FFd3_In
    );
  mac_control_PHY_status_MII_Interface_cs_FFd3_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd3_FROM,
      O => mac_control_PHY_status_MII_Interface_N70564
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_170_61 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_37_CYINIT,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_39,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_170
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_391 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_mdccnt_37,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_39
    );
  mac_control_PHY_status_MII_Interface_n00101 : X_LUT4
    generic map(
      INIT => X"3130"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_mdccnt_37,
      ADR1 => RESET_IBUF,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => MDC_OBUF,
      O => mac_control_PHY_status_MII_Interface_mdccnt_37_GROM
    );
  mac_control_PHY_status_MII_Interface_mdccnt_37_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_37_GROM,
      O => mac_control_PHY_status_MII_Interface_n0010
    );
  mac_control_PHY_status_MII_Interface_mdccnt_37_CYINIT_62 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_192,
      O => mac_control_PHY_status_MII_Interface_mdccnt_37_CYINIT
    );
  mac_control_PHY_status_MII_Interface_n00131 : X_LUT4
    generic map(
      INIT => X"3332"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => RESET_IBUF,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd3,
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd4,
      O => mac_control_PHY_status_MII_Interface_n0013_FROM
    );
  mac_control_PHY_status_MII_Interface_n00111 : X_LUT4
    generic map(
      INIT => X"0F0A"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd4,
      ADR1 => VCC,
      ADR2 => RESET_IBUF,
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd3,
      O => mac_control_PHY_status_MII_Interface_n0013_GROM
    );
  mac_control_PHY_status_MII_Interface_n0013_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0013_FROM,
      O => mac_control_PHY_status_MII_Interface_n0013
    );
  mac_control_PHY_status_MII_Interface_n0013_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0013_GROM,
      O => mac_control_PHY_status_MII_Interface_n0011
    );
  tx_output_crc_loigc_Mxor_CO_10_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(2),
      ADR1 => tx_output_crc_loigc_n0118(0),
      ADR2 => tx_output_crc_loigc_Mxor_CO_7_Xo(1),
      ADR3 => tx_output_crc_loigc_n0118(1),
      O => tx_output_crcl_10_FROM
    );
  tx_output_n0034_10_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crc_10_Q,
      O => tx_output_n0034_10_Q
    );
  tx_output_crcl_10_XUSED : X_BUF
    port map (
      I => tx_output_crcl_10_FROM,
      O => tx_output_crc_10_Q
    );
  mac_control_PHY_status_MII_Interface_n00151 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd2,
      O => mac_control_PHY_status_MII_Interface_n0015_GROM
    );
  mac_control_PHY_status_MII_Interface_n0015_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0015_GROM,
      O => mac_control_PHY_status_MII_Interface_n0015
    );
  rx_output_mdl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_11_FFY_RST
    );
  rx_output_mdl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(10),
      CE => rx_output_mdl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_11_FFY_RST,
      O => rx_output_mdl(10)
    );
  rx_output_mdl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_11_CEMUXNOT
    );
  rx_output_mdl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_21_FFY_RST
    );
  rx_output_mdl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(20),
      CE => rx_output_mdl_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_21_FFY_RST,
      O => rx_output_mdl(20)
    );
  rx_output_mdl_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_21_CEMUXNOT
    );
  rx_input_fifo_fifo_BU145 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1583,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1596_FFY_RST,
      O => rx_input_fifo_fifo_N1597
    );
  rx_input_fifo_fifo_N1596_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1596_FFY_RST
    );
  rx_output_mdl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_13_FFY_RST
    );
  rx_output_mdl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(12),
      CE => rx_output_mdl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_13_FFY_RST,
      O => rx_output_mdl(12)
    );
  rx_output_mdl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_13_CEMUXNOT
    );
  rx_input_fifo_fifo_BU154 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N1580,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1594_FFX_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1594
    );
  rx_input_fifo_fifo_N1594_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1594_FFX_SET
    );
  rx_output_mdl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_31_FFY_RST
    );
  rx_output_mdl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(30),
      CE => rx_output_mdl_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_31_FFY_RST,
      O => rx_output_mdl(30)
    );
  rx_output_mdl_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_31_CEMUXNOT
    );
  rx_output_mdl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_23_FFY_RST
    );
  rx_output_mdl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(22),
      CE => rx_output_mdl_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_23_FFY_RST,
      O => rx_output_mdl(22)
    );
  rx_output_mdl_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_23_CEMUXNOT
    );
  rx_input_fifo_fifo_BU120 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2372,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1525_FFX_RST,
      O => rx_input_fifo_fifo_N1525
    );
  rx_input_fifo_fifo_N1525_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1525_FFX_RST
    );
  rx_output_mdl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_15_FFY_RST
    );
  rx_output_mdl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(14),
      CE => rx_output_mdl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_15_FFY_RST,
      O => rx_output_mdl(14)
    );
  rx_output_mdl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_15_CEMUXNOT
    );
  rx_output_mdl_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_25_CEMUXNOT
    );
  rx_output_mdl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_17_FFY_RST
    );
  rx_output_mdl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(16),
      CE => rx_output_mdl_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_17_FFY_RST,
      O => rx_output_mdl(16)
    );
  rx_output_mdl_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_17_CEMUXNOT
    );
  rx_output_mdl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_27_FFY_RST
    );
  rx_output_mdl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(26),
      CE => rx_output_mdl_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_27_FFY_RST,
      O => rx_output_mdl(26)
    );
  rx_output_mdl_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_27_CEMUXNOT
    );
  rx_output_mdl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_19_FFY_RST
    );
  rx_output_mdl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(18),
      CE => rx_output_mdl_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_19_FFY_RST,
      O => rx_output_mdl(18)
    );
  rx_output_mdl_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_19_CEMUXNOT
    );
  rx_output_mdl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_29_FFY_RST
    );
  rx_output_mdl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(28),
      CE => rx_output_mdl_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_29_FFY_RST,
      O => rx_output_mdl(28)
    );
  rx_output_mdl_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_29_CEMUXNOT
    );
  rx_output_lmasell_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lmasell_FFY_RST
    );
  rx_output_lmasell_63 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd7,
      CE => rx_output_lmasell_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lmasell_FFY_RST,
      O => rx_output_lmasell
    );
  rx_output_lmasell_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lmasell_CEMUXNOT
    );
  tx_input_enable_LOGIC_ONE_64 : X_ONE
    port map (
      O => tx_input_enable_LOGIC_ONE
    );
  rx_input_memio_crccomb_Mxor_CO_2_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crc_0_Q,
      ADR1 => rx_input_memio_crccomb_n0124(0),
      ADR2 => rx_input_memio_crccomb_n0122(0),
      ADR3 => rx_input_memio_crccomb_n0118(1),
      O => rx_input_memio_crcl_2_FROM
    );
  rx_input_memio_n0048_2_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_2_Q,
      O => rx_input_memio_n0048_2_Q
    );
  rx_input_memio_crcl_2_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_2_FROM,
      O => rx_input_memio_crc_2_Q
    );
  rx_input_memio_crccomb_Mxor_CO_3_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0118(1),
      ADR1 => rx_input_memio_crccomb_n0122(0),
      ADR2 => rx_input_memio_crccomb_n0124(0),
      ADR3 => rx_input_memio_crccomb_n0124(1),
      O => rx_input_memio_crcl_3_FROM
    );
  rx_input_memio_n0048_3_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_3_Q,
      O => rx_input_memio_n0048_3_Q
    );
  rx_input_memio_crcl_3_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_3_FROM,
      O => rx_input_memio_crc_3_Q
    );
  tx_output_ldata_6_26_SW0 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => q2(30),
      ADR1 => tx_output_cs_FFd4_1,
      ADR2 => tx_output_cs_FFd6_1,
      ADR3 => q2(14),
      O => tx_output_data_6_FROM
    );
  tx_output_ldata_6_26 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => tx_output_CHOICE1670,
      ADR1 => tx_output_cs_FFd5_1,
      ADR2 => q2(22),
      ADR3 => tx_output_N81018,
      O => tx_output_ldata(6)
    );
  tx_output_data_6_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_data_6_CEMUXNOT
    );
  tx_output_data_6_XUSED : X_BUF
    port map (
      I => tx_output_data_6_FROM,
      O => tx_output_N81018
    );
  txfifofull_LOGIC_ONE_65 : X_ONE
    port map (
      O => txfifofull_LOGIC_ONE
    );
  tx_output_ldata_7_26_SW0 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => tx_output_cs_FFd4_1,
      ADR1 => q2(15),
      ADR2 => tx_output_cs_FFd6_1,
      ADR3 => q2(31),
      O => tx_output_data_7_FROM
    );
  tx_output_ldata_7_26 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => q2(23),
      ADR1 => tx_output_cs_FFd5_1,
      ADR2 => tx_output_CHOICE1658,
      ADR3 => tx_output_N81014,
      O => tx_output_ldata(7)
    );
  tx_output_data_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_data_7_CEMUXNOT
    );
  tx_output_data_7_XUSED : X_BUF
    port map (
      I => tx_output_data_7_FROM,
      O => tx_output_N81014
    );
  tx_output_bcntl_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bcntl_2_CEMUXNOT
    );
  tx_output_bcntl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_4_FFY_RST
    );
  tx_output_bcntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_41,
      CE => tx_output_bcntl_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_4_FFY_RST,
      O => tx_output_bcntl(3)
    );
  tx_output_bcntl_4_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bcntl_4_CEMUXNOT
    );
  tx_output_bcntl_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_6_FFY_RST
    );
  tx_output_bcntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_43,
      CE => tx_output_bcntl_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_6_FFY_RST,
      O => tx_output_bcntl(5)
    );
  tx_output_bcntl_6_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bcntl_6_CEMUXNOT
    );
  rxfbbp_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_1_FFY_RST
    );
  rx_output_bpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(0),
      CE => rxfbbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_1_FFY_RST,
      O => rxfbbp(0)
    );
  rxfbbp_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_1_CEMUXNOT
    );
  tx_output_bcntl_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_8_FFY_RST
    );
  tx_output_bcntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_45,
      CE => tx_output_bcntl_8_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_8_FFY_RST,
      O => tx_output_bcntl(7)
    );
  tx_output_bcntl_8_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bcntl_8_CEMUXNOT
    );
  rxfbbp_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_3_FFY_RST
    );
  rx_output_bpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(2),
      CE => rxfbbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_3_FFY_RST,
      O => rxfbbp(2)
    );
  rxfbbp_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_3_CEMUXNOT
    );
  tx_output_datal_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_1_FFY_RST
    );
  tx_output_datal_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(0),
      CE => tx_output_datal_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_1_FFY_RST,
      O => tx_output_datal(0)
    );
  tx_output_datal_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_datal_1_CEMUXNOT
    );
  tx_output_bcntl_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_10_FFY_RST
    );
  tx_output_bcntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_47,
      CE => tx_output_bcntl_10_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_10_FFY_RST,
      O => tx_output_bcntl(9)
    );
  tx_output_bcntl_10_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bcntl_10_CEMUXNOT
    );
  rxfbbp_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_5_FFY_RST
    );
  rx_output_bpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(4),
      CE => rxfbbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_5_FFY_RST,
      O => rxfbbp(4)
    );
  rxfbbp_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_5_CEMUXNOT
    );
  tx_output_datal_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_3_FFY_RST
    );
  tx_output_datal_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(2),
      CE => tx_output_datal_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_3_FFY_RST,
      O => tx_output_datal(2)
    );
  tx_output_datal_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_datal_3_CEMUXNOT
    );
  rxfbbp_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_7_FFY_RST
    );
  rx_output_bpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(6),
      CE => rxfbbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_7_FFY_RST,
      O => rxfbbp(6)
    );
  rxfbbp_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_7_CEMUXNOT
    );
  tx_output_datal_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_5_FFY_RST
    );
  tx_output_datal_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(4),
      CE => tx_output_datal_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_5_FFY_RST,
      O => tx_output_datal(4)
    );
  tx_output_datal_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_datal_5_CEMUXNOT
    );
  tx_output_crcl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_11_FFY_RST
    );
  tx_output_crcl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_11_1_O,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_11_FFY_RST,
      O => tx_output_crcl(11)
    );
  tx_output_crc_loigc_Mxor_CO_11_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0124(1),
      ADR1 => tx_output_crc_loigc_n0115(0),
      ADR2 => tx_output_crc_loigc_Mxor_CO_23_Xo(0),
      ADR3 => tx_output_crcl(3),
      O => tx_output_crcl_11_FROM
    );
  tx_output_n0034_11_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_11_Q,
      O => tx_output_n0034_11_1_O
    );
  tx_output_crcl_11_XUSED : X_BUF
    port map (
      I => tx_output_crcl_11_FROM,
      O => tx_output_crc_11_Q
    );
  rxfbbp_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rxfbbp_9_CEMUXNOT
    );
  rx_input_fifo_fifo_BU99 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2252,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1527_FFY_RST,
      O => rx_input_fifo_fifo_N1528
    );
  rx_input_fifo_fifo_N1527_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1527_FFY_RST
    );
  tx_output_datal_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_7_FFY_RST
    );
  tx_output_datal_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(6),
      CE => tx_output_datal_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_7_FFY_RST,
      O => tx_output_datal(6)
    );
  tx_output_datal_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_datal_7_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_1_FFY_RST
    );
  mac_control_rxfifowerr_cntl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(0),
      CE => mac_control_rxfifowerr_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_1_FFY_RST,
      O => mac_control_rxfifowerr_cntl(0)
    );
  mac_control_rxfifowerr_cntl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_1_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_3_FFY_RST
    );
  mac_control_rxfifowerr_cntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(2),
      CE => mac_control_rxfifowerr_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_3_FFY_RST,
      O => mac_control_rxfifowerr_cntl(2)
    );
  mac_control_rxfifowerr_cntl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_3_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_5_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_7_FFY_RST
    );
  mac_control_rxfifowerr_cntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(6),
      CE => mac_control_rxfifowerr_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_7_FFY_RST,
      O => mac_control_rxfifowerr_cntl(6)
    );
  mac_control_rxfifowerr_cntl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_7_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_9_FFY_RST
    );
  mac_control_rxfifowerr_cntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(8),
      CE => mac_control_rxfifowerr_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_9_FFY_RST,
      O => mac_control_rxfifowerr_cntl(8)
    );
  mac_control_rxfifowerr_cntl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_cntl_9_CEMUXNOT
    );
  rx_output_denll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_denll_FFY_RST
    );
  rx_output_denll_66 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_denl,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => rx_output_denll_FFY_RST,
      O => rx_output_denll
    );
  rx_output_mdl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_1_FFY_RST
    );
  rx_output_mdl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(0),
      CE => rx_output_mdl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_1_FFY_RST,
      O => rx_output_mdl(0)
    );
  rx_output_mdl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_1_CEMUXNOT
    );
  rx_input_fifo_fifo_BU59 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1860,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N13_FFY_RST,
      O => rx_input_fifo_fifo_N12
    );
  rx_input_fifo_fifo_N13_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N13_FFY_RST
    );
  rx_output_len_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_3_FFY_RST
    );
  rx_output_len_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(2),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_3_FFY_RST,
      O => rx_output_len(2)
    );
  rx_input_fifo_fifo_BU65 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1861,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N11_FFX_RST,
      O => rx_input_fifo_fifo_N11
    );
  rx_input_fifo_fifo_N11_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N11_FFX_RST
    );
  rx_output_mdl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_3_FFY_RST
    );
  rx_output_mdl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(2),
      CE => rx_output_mdl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_3_FFY_RST,
      O => rx_output_mdl(2)
    );
  rx_output_mdl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_3_CEMUXNOT
    );
  rx_output_mdl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_5_FFY_RST
    );
  rx_output_mdl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(4),
      CE => rx_output_mdl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_5_FFY_RST,
      O => rx_output_mdl(4)
    );
  rx_output_mdl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_5_CEMUXNOT
    );
  rx_output_len_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_7_FFY_RST
    );
  rx_output_len_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(6),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_7_FFY_RST,
      O => rx_output_len(6)
    );
  rx_output_mdl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_7_FFY_RST
    );
  rx_output_mdl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(6),
      CE => rx_output_mdl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_7_FFY_RST,
      O => rx_output_mdl(6)
    );
  rx_output_mdl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_7_CEMUXNOT
    );
  rx_output_len_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_9_FFY_RST
    );
  rx_output_len_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(8),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_9_FFY_RST,
      O => rx_output_len(8)
    );
  rx_output_mdl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_9_FFY_RST
    );
  rx_output_mdl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(8),
      CE => rx_output_mdl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_9_FFY_RST,
      O => rx_output_mdl(8)
    );
  rx_output_mdl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_mdl_9_CEMUXNOT
    );
  tx_output_ltxd_0_SW0 : X_LUT4
    generic map(
      INIT => X"FCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_datal(0),
      ADR2 => tx_output_outselll(1),
      ADR3 => tx_output_outselll(0),
      O => tx_output_N70308_FROM
    );
  tx_output_ltxd_0_Q : X_LUT4
    generic map(
      INIT => X"FEEE"
    )
    port map (
      ADR0 => tx_output_outselll(2),
      ADR1 => tx_output_N70308,
      ADR2 => tx_output_ncrcbytel(7),
      ADR3 => tx_output_outselll(3),
      O => tx_output_N70308_GROM
    );
  tx_output_N70308_XUSED : X_BUF
    port map (
      I => tx_output_N70308_FROM,
      O => tx_output_N70308
    );
  tx_output_N70308_YUSED : X_BUF
    port map (
      I => tx_output_N70308_GROM,
      O => tx_output_ltxd(0)
    );
  rx_input_GMII_ro_LOGIC_ONE_67 : X_ONE
    port map (
      O => rx_input_GMII_ro_LOGIC_ONE
    );
  rx_input_memio_crccomb_Mxor_CO_4_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0124(1),
      ADR1 => rx_input_memio_crccomb_n0115(0),
      ADR2 => rx_input_memio_crc_0_Q,
      ADR3 => rx_input_memio_crccomb_n0118(1),
      O => rx_input_memio_crcl_4_FROM
    );
  rx_input_memio_n0048_4_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_4_Q,
      O => rx_input_memio_n0048_4_1_O
    );
  rx_input_memio_crcl_4_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_4_FROM,
      O => rx_input_memio_crc_4_Q
    );
  tx_output_outselll_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_outselll_1_CEMUXNOT
    );
  tx_output_outselll_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outselll_3_FFY_RST
    );
  tx_output_outselll_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_outsell(2),
      CE => tx_output_outselll_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outselll_3_FFY_RST,
      O => tx_output_outselll(2)
    );
  tx_output_outselll_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_outselll_3_CEMUXNOT
    );
  tx_output_ltxd_2_SW0 : X_LUT4
    generic map(
      INIT => X"FAF0"
    )
    port map (
      ADR0 => tx_output_datal(2),
      ADR1 => VCC,
      ADR2 => tx_output_outselll(1),
      ADR3 => tx_output_outselll(0),
      O => tx_output_N70281_FROM
    );
  tx_output_ltxd_2_Q : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => tx_output_outselll(3),
      ADR1 => tx_output_outselll(2),
      ADR2 => tx_output_ncrcbytel(5),
      ADR3 => tx_output_N70281,
      O => tx_output_N70281_GROM
    );
  tx_output_N70281_XUSED : X_BUF
    port map (
      I => tx_output_N70281_FROM,
      O => tx_output_N70281
    );
  tx_output_N70281_YUSED : X_BUF
    port map (
      I => tx_output_N70281_GROM,
      O => tx_output_ltxd(2)
    );
  mac_control_txf_cntl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_11_CEMUXNOT
    );
  mac_control_txf_cntl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_21_FFY_RST
    );
  mac_control_txf_cntl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(20),
      CE => mac_control_txf_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_21_FFY_RST,
      O => mac_control_txf_cntl(20)
    );
  mac_control_txf_cntl_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_21_CEMUXNOT
    );
  mac_control_txf_cntl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_13_FFY_RST
    );
  mac_control_txf_cntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(12),
      CE => mac_control_txf_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_13_FFY_RST,
      O => mac_control_txf_cntl(12)
    );
  mac_control_txf_cntl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_13_CEMUXNOT
    );
  tx_output_ltxd_4_SW0 : X_LUT4
    generic map(
      INIT => X"ECEC"
    )
    port map (
      ADR0 => tx_output_outselll(0),
      ADR1 => tx_output_outselll(1),
      ADR2 => tx_output_datal(4),
      ADR3 => VCC,
      O => tx_output_N70254_FROM
    );
  tx_output_ltxd_4_Q : X_LUT4
    generic map(
      INIT => X"FEFC"
    )
    port map (
      ADR0 => tx_output_ncrcbytel(3),
      ADR1 => tx_output_N70254,
      ADR2 => tx_output_outselll(2),
      ADR3 => tx_output_outselll(3),
      O => tx_output_N70254_GROM
    );
  tx_output_N70254_XUSED : X_BUF
    port map (
      I => tx_output_N70254_FROM,
      O => tx_output_N70254
    );
  tx_output_N70254_YUSED : X_BUF
    port map (
      I => tx_output_N70254_GROM,
      O => tx_output_ltxd(4)
    );
  mac_control_txf_cntl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_31_FFY_RST
    );
  mac_control_txf_cntl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(30),
      CE => mac_control_txf_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_31_FFY_RST,
      O => mac_control_txf_cntl(30)
    );
  mac_control_txf_cntl_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_31_CEMUXNOT
    );
  mac_control_txf_cntl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_23_FFY_RST
    );
  mac_control_txf_cntl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(22),
      CE => mac_control_txf_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_23_FFY_RST,
      O => mac_control_txf_cntl(22)
    );
  mac_control_txf_cntl_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_23_CEMUXNOT
    );
  mac_control_txf_cntl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_15_FFY_RST
    );
  mac_control_txf_cntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(14),
      CE => mac_control_txf_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_15_FFY_RST,
      O => mac_control_txf_cntl(14)
    );
  mac_control_txf_cntl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_15_CEMUXNOT
    );
  mac_control_txf_cntl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_25_FFY_RST
    );
  mac_control_txf_cntl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(24),
      CE => mac_control_txf_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_25_FFY_RST,
      O => mac_control_txf_cntl(24)
    );
  mac_control_txf_cntl_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_25_CEMUXNOT
    );
  mac_control_txf_cntl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_17_FFY_RST
    );
  mac_control_txf_cntl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(16),
      CE => mac_control_txf_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_17_FFY_RST,
      O => mac_control_txf_cntl(16)
    );
  mac_control_txf_cntl_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_17_CEMUXNOT
    );
  mac_control_addr_0_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_0_1_FFY_RST
    );
  mac_control_addr_0_1_68 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_Mshreg_sinlll_102,
      CE => mac_control_n0010,
      CLK => clksl,
      SET => GND,
      RST => mac_control_addr_0_1_FFY_RST,
      O => mac_control_addr_0_1
    );
  mac_control_txf_cntl_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_27_CEMUXNOT
    );
  mac_control_txf_cntl_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_19_CEMUXNOT
    );
  mac_control_txf_cntl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_29_FFY_RST
    );
  mac_control_txf_cntl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(28),
      CE => mac_control_txf_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_29_FFY_RST,
      O => mac_control_txf_cntl(28)
    );
  mac_control_txf_cntl_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_29_CEMUXNOT
    );
  tx_output_ldata_2_17 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => q2(2),
      ADR1 => tx_output_cs_FFd4_1,
      ADR2 => tx_output_cs_FFd6_1,
      ADR3 => tx_output_cs_FFd5_1,
      O => tx_output_CHOICE1730_FROM
    );
  tx_output_ldata_0_17 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => q2(0),
      ADR1 => tx_output_cs_FFd4_1,
      ADR2 => tx_output_cs_FFd5_1,
      ADR3 => tx_output_cs_FFd6_1,
      O => tx_output_CHOICE1730_GROM
    );
  tx_output_CHOICE1730_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1730_FROM,
      O => tx_output_CHOICE1730
    );
  tx_output_CHOICE1730_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1730_GROM,
      O => tx_output_CHOICE1742
    );
  tx_output_ldata_5_17 : X_LUT4
    generic map(
      INIT => X"0100"
    )
    port map (
      ADR0 => tx_output_cs_FFd6_1,
      ADR1 => tx_output_cs_FFd4_1,
      ADR2 => tx_output_cs_FFd5_1,
      ADR3 => q2(5),
      O => tx_output_CHOICE1694_FROM
    );
  tx_output_ldata_1_17 : X_LUT4
    generic map(
      INIT => X"0004"
    )
    port map (
      ADR0 => tx_output_cs_FFd4_1,
      ADR1 => q2(1),
      ADR2 => tx_output_cs_FFd5_1,
      ADR3 => tx_output_cs_FFd6_1,
      O => tx_output_CHOICE1694_GROM
    );
  tx_output_CHOICE1694_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1694_FROM,
      O => tx_output_CHOICE1694
    );
  tx_output_CHOICE1694_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1694_GROM,
      O => tx_output_CHOICE1718
    );
  tx_output_ldata_7_17 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => q2(7),
      ADR1 => tx_output_cs_FFd4_1,
      ADR2 => tx_output_cs_FFd5_1,
      ADR3 => tx_output_cs_FFd6_1,
      O => tx_output_CHOICE1658_FROM
    );
  tx_output_ldata_3_17 : X_LUT4
    generic map(
      INIT => X"0010"
    )
    port map (
      ADR0 => tx_output_cs_FFd5_1,
      ADR1 => tx_output_cs_FFd6_1,
      ADR2 => q2(3),
      ADR3 => tx_output_cs_FFd4_1,
      O => tx_output_CHOICE1658_GROM
    );
  tx_output_CHOICE1658_XUSED : X_BUF
    port map (
      I => tx_output_CHOICE1658_FROM,
      O => tx_output_CHOICE1658
    );
  tx_output_CHOICE1658_YUSED : X_BUF
    port map (
      I => tx_output_CHOICE1658_GROM,
      O => tx_output_CHOICE1706
    );
  tx_output_ltxd_6_SW0 : X_LUT4
    generic map(
      INIT => X"EECC"
    )
    port map (
      ADR0 => tx_output_outselll(0),
      ADR1 => tx_output_outselll(1),
      ADR2 => VCC,
      ADR3 => tx_output_datal(6),
      O => tx_output_N70227_FROM
    );
  tx_output_ltxd_6_Q : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => tx_output_outselll(3),
      ADR1 => tx_output_outselll(2),
      ADR2 => tx_output_ncrcbytel(1),
      ADR3 => tx_output_N70227,
      O => tx_output_N70227_GROM
    );
  tx_output_N70227_XUSED : X_BUF
    port map (
      I => tx_output_N70227_FROM,
      O => tx_output_N70227
    );
  tx_output_N70227_YUSED : X_BUF
    port map (
      I => tx_output_N70227_GROM,
      O => tx_output_ltxd(6)
    );
  tx_output_ltxd_7_SW0 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_outselll(0),
      ADR2 => VCC,
      ADR3 => tx_output_datal(7),
      O => tx_output_N70079_FROM
    );
  tx_output_ltxd_7_Q : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => tx_output_outselll(2),
      ADR1 => tx_output_outselll(3),
      ADR2 => tx_output_ncrcbytel(0),
      ADR3 => tx_output_N70079,
      O => tx_output_N70079_GROM
    );
  tx_output_N70079_XUSED : X_BUF
    port map (
      I => tx_output_N70079_FROM,
      O => tx_output_N70079
    );
  tx_output_N70079_YUSED : X_BUF
    port map (
      I => tx_output_N70079_GROM,
      O => tx_output_ltxd(7)
    );
  rx_input_fifo_fifo_BU148 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1582,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1596_FFX_RST,
      O => rx_input_fifo_fifo_N1596
    );
  rx_input_fifo_fifo_N1596_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1596_FFX_RST
    );
  RESET_IBUF_1_69 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => VCC,
      O => RESET_IBUF_1_FROM
    );
  tx_input_n00331 : X_LUT4
    generic map(
      INIT => X"00FE"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => tx_input_cs_FFd5,
      ADR2 => tx_input_cs_FFd9,
      ADR3 => RESET_IBUF_1,
      O => RESET_IBUF_1_GROM
    );
  RESET_IBUF_1_XUSED : X_BUF
    port map (
      I => RESET_IBUF_1_FROM,
      O => RESET_IBUF_1
    );
  RESET_IBUF_1_YUSED : X_BUF
    port map (
      I => RESET_IBUF_1_GROM,
      O => tx_input_n0033
    );
  RESET_IBUF_2_70 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => VCC,
      O => RESET_IBUF_2_FROM
    );
  rx_input_RESET_1_71 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => RESET_IBUF_2,
      O => RESET_IBUF_2_GROM
    );
  RESET_IBUF_2_XUSED : X_BUF
    port map (
      I => RESET_IBUF_2_FROM,
      O => RESET_IBUF_2
    );
  RESET_IBUF_2_YUSED : X_BUF
    port map (
      I => RESET_IBUF_2_GROM,
      O => rx_input_RESET_1
    );
  mac_control_PHY_status_MII_Interface_iobuffer_OBUFT : X_TRI
    port map (
      I => MDIO_OUTMUX,
      CTL => MDIO_ENABLE,
      O => MDIO
    );
  MDIO_ENABLEINV : X_INV
    port map (
      I => MDIO_TORGTS,
      O => MDIO_ENABLE
    );
  MDIO_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => mac_control_PHY_status_MII_Interface_sts,
      O => MDIO_TORGTS
    );
  MDIO_OUTMUX_72 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_sout,
      O => MDIO_OUTMUX
    );
  mac_control_PHY_status_MII_Interface_iobuffer_IBUF : X_BUF
    port map (
      I => MDIO,
      O => mac_control_PHY_status_MII_Interface_sin
    );
  rx_output_DOUT_10_OBUF_73 : X_TRI
    port map (
      I => DOUT_10_OUTMUX,
      CTL => DOUT_10_ENABLE,
      O => DOUT(10)
    );
  DOUT_10_ENABLEINV : X_INV
    port map (
      I => DOUT_10_TORGTS,
      O => DOUT_10_ENABLE
    );
  DOUT_10_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_10_TORGTS
    );
  DOUT_10_OUTMUX_74 : X_BUF
    port map (
      I => rx_output_DOUT_10_OBUF,
      O => DOUT_10_OUTMUX
    );
  DOUT_10_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(10),
      O => DOUT_10_OD
    );
  rx_output_DOUT_11_OBUF_75 : X_TRI
    port map (
      I => DOUT_11_OUTMUX,
      CTL => DOUT_11_ENABLE,
      O => DOUT(11)
    );
  DOUT_11_ENABLEINV : X_INV
    port map (
      I => DOUT_11_TORGTS,
      O => DOUT_11_ENABLE
    );
  DOUT_11_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_11_TORGTS
    );
  DOUT_11_OUTMUX_76 : X_BUF
    port map (
      I => rx_output_DOUT_11_OBUF,
      O => DOUT_11_OUTMUX
    );
  DOUT_11_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(11),
      O => DOUT_11_OD
    );
  rx_output_DOUT_12_OBUF_77 : X_TRI
    port map (
      I => DOUT_12_OUTMUX,
      CTL => DOUT_12_ENABLE,
      O => DOUT(12)
    );
  DOUT_12_ENABLEINV : X_INV
    port map (
      I => DOUT_12_TORGTS,
      O => DOUT_12_ENABLE
    );
  DOUT_12_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_12_TORGTS
    );
  DOUT_12_OUTMUX_78 : X_BUF
    port map (
      I => rx_output_DOUT_12_OBUF,
      O => DOUT_12_OUTMUX
    );
  DOUT_12_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(12),
      O => DOUT_12_OD
    );
  rx_output_DOUT_13_OBUF_79 : X_TRI
    port map (
      I => DOUT_13_OUTMUX,
      CTL => DOUT_13_ENABLE,
      O => DOUT(13)
    );
  DOUT_13_ENABLEINV : X_INV
    port map (
      I => DOUT_13_TORGTS,
      O => DOUT_13_ENABLE
    );
  DOUT_13_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_13_TORGTS
    );
  DOUT_13_OUTMUX_80 : X_BUF
    port map (
      I => rx_output_DOUT_13_OBUF,
      O => DOUT_13_OUTMUX
    );
  DOUT_13_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(13),
      O => DOUT_13_OD
    );
  rx_input_fifo_fifo_BU106 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2292,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1527_FFX_RST,
      O => rx_input_fifo_fifo_N1527
    );
  rx_input_fifo_fifo_N1527_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1527_FFX_RST
    );
  rx_output_DOUT_14_OBUF_81 : X_TRI
    port map (
      I => DOUT_14_OUTMUX,
      CTL => DOUT_14_ENABLE,
      O => DOUT(14)
    );
  DOUT_14_ENABLEINV : X_INV
    port map (
      I => DOUT_14_TORGTS,
      O => DOUT_14_ENABLE
    );
  DOUT_14_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_14_TORGTS
    );
  DOUT_14_OUTMUX_82 : X_BUF
    port map (
      I => rx_output_DOUT_14_OBUF,
      O => DOUT_14_OUTMUX
    );
  DOUT_14_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(14),
      O => DOUT_14_OD
    );
  rx_output_DOUT_15_OBUF_83 : X_TRI
    port map (
      I => DOUT_15_OUTMUX,
      CTL => DOUT_15_ENABLE,
      O => DOUT(15)
    );
  DOUT_15_ENABLEINV : X_INV
    port map (
      I => DOUT_15_TORGTS,
      O => DOUT_15_ENABLE
    );
  DOUT_15_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_15_TORGTS
    );
  DOUT_15_OUTMUX_84 : X_BUF
    port map (
      I => rx_output_DOUT_15_OBUF,
      O => DOUT_15_OUTMUX
    );
  DOUT_15_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(15),
      O => DOUT_15_OD
    );
  MDC_OBUF_85 : X_TRI
    port map (
      I => MDC_OUTMUX,
      CTL => MDC_ENABLE,
      O => MDC
    );
  MDC_ENABLEINV : X_INV
    port map (
      I => MDC_TORGTS,
      O => MDC_ENABLE
    );
  MDC_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MDC_TORGTS
    );
  MDC_OUTMUX_86 : X_BUF
    port map (
      I => MDC_OBUF,
      O => MDC_OUTMUX
    );
  SCS_IMUX : X_BUF
    port map (
      I => SCS_IBUF_1,
      O => SCS_IBUF
    );
  SCS_IBUF_87 : X_BUF
    port map (
      I => SCS,
      O => SCS_IBUF_1
    );
  SIN_IMUX : X_BUF
    port map (
      I => SIN_IBUF_2,
      O => SIN_IBUF
    );
  SIN_IBUF_88 : X_BUF
    port map (
      I => SIN,
      O => SIN_IBUF_2
    );
  mac_control_LED100_OBUF_89 : X_TRI
    port map (
      I => LED100_OUTMUX,
      CTL => LED100_ENABLE,
      O => LED100
    );
  LED100_ENABLEINV : X_INV
    port map (
      I => LED100_TORGTS,
      O => LED100_ENABLE
    );
  LED100_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LED100_TORGTS
    );
  LED100_OUTMUX_90 : X_BUF
    port map (
      I => mac_control_LED100_OBUF,
      O => LED100_OUTMUX
    );
  LED100_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => LED100_OCEMUXNOT
    );
  LED100_OMUX : X_BUF
    port map (
      I => mac_control_n0036,
      O => LED100_OD
    );
  MCLK_OBUF : X_TRI
    port map (
      I => MCLK_OUTMUX,
      CTL => MCLK_ENABLE,
      O => MCLK
    );
  MCLK_ENABLEINV : X_INV
    port map (
      I => MCLK_TORGTS,
      O => MCLK_ENABLE
    );
  MCLK_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MCLK_TORGTS
    );
  MCLK_OUTMUX_91 : X_BUF
    port map (
      I => GTX_CLK_OBUF,
      O => MCLK_OUTMUX
    );
  tx_input_NEWFRAME_IBUF_92 : X_BUF
    port map (
      I => NEWFRAME,
      O => tx_input_NEWFRAME_IBUF
    );
  mac_control_LED1000_OBUF_93 : X_TRI
    port map (
      I => LED1000_OUTMUX,
      CTL => LED1000_ENABLE,
      O => LED1000
    );
  LED1000_ENABLEINV : X_INV
    port map (
      I => LED1000_TORGTS,
      O => LED1000_ENABLE
    );
  LED1000_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LED1000_TORGTS
    );
  LED1000_OUTMUX_94 : X_BUF
    port map (
      I => mac_control_LED1000_OBUF,
      O => LED1000_OUTMUX
    );
  LED1000_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => LED1000_OCEMUXNOT
    );
  LED1000_OMUX : X_BUF
    port map (
      I => mac_control_n0035,
      O => LED1000_OD
    );
  tx_output_TX_EN_OBUF : X_TRI
    port map (
      I => TX_EN_OUTMUX,
      CTL => TX_EN_ENABLE,
      O => TX_EN
    );
  TX_EN_ENABLEINV : X_INV
    port map (
      I => TX_EN_TORGTS,
      O => TX_EN_ENABLE
    );
  TX_EN_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TX_EN_TORGTS
    );
  TX_EN_OUTMUX_95 : X_BUF
    port map (
      I => tx_output_TXEN,
      O => TX_EN_OUTMUX
    );
  TX_EN_OCEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => TX_EN_OCEMUXNOT
    );
  TX_EN_OMUX : X_BUF
    port map (
      I => tx_output_ltxen3,
      O => TX_EN_OD
    );
  rx_output_DOUTEN_OBUF_96 : X_TRI
    port map (
      I => DOUTEN_OUTMUX,
      CTL => DOUTEN_ENABLE,
      O => DOUTEN
    );
  DOUTEN_ENABLEINV : X_INV
    port map (
      I => DOUTEN_TORGTS,
      O => DOUTEN_ENABLE
    );
  DOUTEN_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUTEN_TORGTS
    );
  DOUTEN_OUTMUX_97 : X_BUF
    port map (
      I => rx_output_DOUTEN_OBUF,
      O => DOUTEN_OUTMUX
    );
  DOUTEN_OMUX : X_BUF
    port map (
      I => rx_output_ldouten2,
      O => DOUTEN_OD
    );
  memcontroller_weout : X_TRI
    port map (
      I => MWE_OUTMUX,
      CTL => MWE_ENABLE,
      O => MWE
    );
  MWE_ENABLEINV : X_INV
    port map (
      I => MWE_TORGTS,
      O => MWE_ENABLE
    );
  MWE_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MWE_TORGTS
    );
  MWE_OUTMUX_98 : X_BUF
    port map (
      I => memcontroller_we,
      O => MWE_OUTMUX
    );
  MWE_OMUX : X_BUF
    port map (
      I => memcontroller_n0149,
      O => MWE_OD
    );
  RESET_IMUX : X_BUF
    port map (
      I => RESET_IBUF_3,
      O => RESET_IBUF
    );
  RESET_IBUF_99 : X_BUF
    port map (
      I => RESET,
      O => RESET_IBUF_3
    );
  rx_output_NEXTFRAME_IBUF_100 : X_BUF
    port map (
      I => NEXTFRAME,
      O => rx_output_NEXTFRAME_IBUF
    );
  mac_control_LEDACT_OBUF_101 : X_TRI
    port map (
      I => LEDACT_OUTMUX,
      CTL => LEDACT_ENABLE,
      O => LEDACT
    );
  LEDACT_ENABLEINV : X_INV
    port map (
      I => LEDACT_TORGTS,
      O => LEDACT_ENABLE
    );
  LEDACT_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDACT_TORGTS
    );
  LEDACT_OUTMUX_102 : X_BUF
    port map (
      I => mac_control_LEDACT_OBUF,
      O => LEDACT_OUTMUX
    );
  LEDACT_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => LEDACT_OCEMUXNOT
    );
  LEDACT_OMUX : X_BUF
    port map (
      I => mac_control_phystat(2),
      O => LEDACT_OD
    );
  tx_output_TXD_0_OBUF_103 : X_TRI
    port map (
      I => TXD_0_OUTMUX,
      CTL => TXD_0_ENABLE,
      O => TXD(0)
    );
  TXD_0_ENABLEINV : X_INV
    port map (
      I => TXD_0_TORGTS,
      O => TXD_0_ENABLE
    );
  TXD_0_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_0_TORGTS
    );
  TXD_0_OUTMUX_104 : X_BUF
    port map (
      I => tx_output_TXD_0_OBUF,
      O => TXD_0_OUTMUX
    );
  TXD_0_OCEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => TXD_0_OCEMUXNOT
    );
  TXD_0_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(0),
      O => TXD_0_OD
    );
  tx_output_TXD_1_OBUF_105 : X_TRI
    port map (
      I => TXD_1_OUTMUX,
      CTL => TXD_1_ENABLE,
      O => TXD(1)
    );
  TXD_1_ENABLEINV : X_INV
    port map (
      I => TXD_1_TORGTS,
      O => TXD_1_ENABLE
    );
  TXD_1_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_1_TORGTS
    );
  TXD_1_OUTMUX_106 : X_BUF
    port map (
      I => tx_output_TXD_1_OBUF,
      O => TXD_1_OUTMUX
    );
  TXD_1_OCEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => TXD_1_OCEMUXNOT
    );
  TXD_1_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(1),
      O => TXD_1_OD
    );
  tx_output_TXD_2_OBUF_107 : X_TRI
    port map (
      I => TXD_2_OUTMUX,
      CTL => TXD_2_ENABLE,
      O => TXD(2)
    );
  TXD_2_ENABLEINV : X_INV
    port map (
      I => TXD_2_TORGTS,
      O => TXD_2_ENABLE
    );
  TXD_2_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_2_TORGTS
    );
  TXD_2_OUTMUX_108 : X_BUF
    port map (
      I => tx_output_TXD_2_OBUF,
      O => TXD_2_OUTMUX
    );
  TXD_2_OCEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => TXD_2_OCEMUXNOT
    );
  TXD_2_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(2),
      O => TXD_2_OD
    );
  tx_output_TXD_3_OBUF_109 : X_TRI
    port map (
      I => TXD_3_OUTMUX,
      CTL => TXD_3_ENABLE,
      O => TXD(3)
    );
  TXD_3_ENABLEINV : X_INV
    port map (
      I => TXD_3_TORGTS,
      O => TXD_3_ENABLE
    );
  TXD_3_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_3_TORGTS
    );
  TXD_3_OUTMUX_110 : X_BUF
    port map (
      I => tx_output_TXD_3_OBUF,
      O => TXD_3_OUTMUX
    );
  TXD_3_OCEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => TXD_3_OCEMUXNOT
    );
  TXD_3_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(3),
      O => TXD_3_OD
    );
  tx_output_TXD_4_OBUF_111 : X_TRI
    port map (
      I => TXD_4_OUTMUX,
      CTL => TXD_4_ENABLE,
      O => TXD(4)
    );
  TXD_4_ENABLEINV : X_INV
    port map (
      I => TXD_4_TORGTS,
      O => TXD_4_ENABLE
    );
  TXD_4_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_4_TORGTS
    );
  TXD_4_OUTMUX_112 : X_BUF
    port map (
      I => tx_output_TXD_4_OBUF,
      O => TXD_4_OUTMUX
    );
  TXD_4_OCEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => TXD_4_OCEMUXNOT
    );
  TXD_4_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(4),
      O => TXD_4_OD
    );
  tx_output_TXD_5_OBUF_113 : X_TRI
    port map (
      I => TXD_5_OUTMUX,
      CTL => TXD_5_ENABLE,
      O => TXD(5)
    );
  TXD_5_ENABLEINV : X_INV
    port map (
      I => TXD_5_TORGTS,
      O => TXD_5_ENABLE
    );
  TXD_5_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_5_TORGTS
    );
  TXD_5_OUTMUX_114 : X_BUF
    port map (
      I => tx_output_TXD_5_OBUF,
      O => TXD_5_OUTMUX
    );
  TXD_5_OCEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => TXD_5_OCEMUXNOT
    );
  TXD_5_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(5),
      O => TXD_5_OD
    );
  tx_output_TXD_6_OBUF_115 : X_TRI
    port map (
      I => TXD_6_OUTMUX,
      CTL => TXD_6_ENABLE,
      O => TXD(6)
    );
  TXD_6_ENABLEINV : X_INV
    port map (
      I => TXD_6_TORGTS,
      O => TXD_6_ENABLE
    );
  TXD_6_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_6_TORGTS
    );
  TXD_6_OUTMUX_116 : X_BUF
    port map (
      I => tx_output_TXD_6_OBUF,
      O => TXD_6_OUTMUX
    );
  TXD_6_OCEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => TXD_6_OCEMUXNOT
    );
  TXD_6_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(6),
      O => TXD_6_OD
    );
  tx_output_TXD_7_OBUF_117 : X_TRI
    port map (
      I => TXD_7_OUTMUX,
      CTL => TXD_7_ENABLE,
      O => TXD(7)
    );
  TXD_7_ENABLEINV : X_INV
    port map (
      I => TXD_7_TORGTS,
      O => TXD_7_ENABLE
    );
  TXD_7_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => TXD_7_TORGTS
    );
  TXD_7_OUTMUX_118 : X_BUF
    port map (
      I => tx_output_TXD_7_OBUF,
      O => TXD_7_OUTMUX
    );
  TXD_7_OCEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => TXD_7_OCEMUXNOT
    );
  TXD_7_OMUX : X_BUF
    port map (
      I => tx_output_ltxd(7),
      O => TXD_7_OD
    );
  mac_control_LEDDPX_OBUF_119 : X_TRI
    port map (
      I => LEDDPX_OUTMUX,
      CTL => LEDDPX_ENABLE,
      O => LEDDPX
    );
  LEDDPX_ENABLEINV : X_INV
    port map (
      I => LEDDPX_TORGTS,
      O => LEDDPX_ENABLE
    );
  LEDDPX_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDDPX_TORGTS
    );
  LEDDPX_OUTMUX_120 : X_BUF
    port map (
      I => mac_control_LEDDPX_OBUF,
      O => LEDDPX_OUTMUX
    );
  LEDDPX_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => LEDDPX_OCEMUXNOT
    );
  LEDDPX_OMUX : X_BUF
    port map (
      I => mac_control_phystat(1),
      O => LEDDPX_OD
    );
  rx_input_GMII_RXD_0_IBUF_121 : X_BUF
    port map (
      I => RXD(0),
      O => rx_input_GMII_RXD_0_IBUF
    );
  rx_input_GMII_RXD_1_IBUF_122 : X_BUF
    port map (
      I => RXD(1),
      O => rx_input_GMII_RXD_1_IBUF
    );
  rx_input_GMII_RXD_2_IBUF_123 : X_BUF
    port map (
      I => RXD(2),
      O => rx_input_GMII_RXD_2_IBUF
    );
  rx_input_GMII_RXD_3_IBUF_124 : X_BUF
    port map (
      I => RXD(3),
      O => rx_input_GMII_RXD_3_IBUF
    );
  rx_input_GMII_RXD_4_IBUF_125 : X_BUF
    port map (
      I => RXD(4),
      O => rx_input_GMII_RXD_4_IBUF
    );
  rx_input_GMII_RXD_5_IBUF_126 : X_BUF
    port map (
      I => RXD(5),
      O => rx_input_GMII_RXD_5_IBUF
    );
  rx_input_GMII_RXD_6_IBUF_127 : X_BUF
    port map (
      I => RXD(6),
      O => rx_input_GMII_RXD_6_IBUF
    );
  rx_input_GMII_RXD_7_IBUF_128 : X_BUF
    port map (
      I => RXD(7),
      O => rx_input_GMII_RXD_7_IBUF
    );
  tx_input_DIN_10_IBUF_129 : X_BUF
    port map (
      I => DIN(10),
      O => tx_input_DIN_10_IBUF
    );
  tx_input_DIN_11_IBUF_130 : X_BUF
    port map (
      I => DIN(11),
      O => tx_input_DIN_11_IBUF
    );
  tx_input_DIN_12_IBUF_131 : X_BUF
    port map (
      I => DIN(12),
      O => tx_input_DIN_12_IBUF
    );
  rx_input_fifo_fifo_BU92 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2212,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1530_FFY_RST,
      O => rx_input_fifo_fifo_N1529
    );
  rx_input_fifo_fifo_N1530_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1530_FFY_RST
    );
  tx_input_DIN_13_IBUF_132 : X_BUF
    port map (
      I => DIN(13),
      O => tx_input_DIN_13_IBUF
    );
  rx_input_fifo_fifo_BU53 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1859,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N13_FFX_RST,
      O => rx_input_fifo_fifo_N13
    );
  rx_input_fifo_fifo_N13_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N13_FFX_RST
    );
  tx_input_DIN_14_IBUF_133 : X_BUF
    port map (
      I => DIN(14),
      O => tx_input_DIN_14_IBUF
    );
  tx_input_DIN_15_IBUF_134 : X_BUF
    port map (
      I => DIN(15),
      O => tx_input_DIN_15_IBUF
    );
  rx_output_DOUT_0_OBUF_135 : X_TRI
    port map (
      I => DOUT_0_OUTMUX,
      CTL => DOUT_0_ENABLE,
      O => DOUT(0)
    );
  DOUT_0_ENABLEINV : X_INV
    port map (
      I => DOUT_0_TORGTS,
      O => DOUT_0_ENABLE
    );
  DOUT_0_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_0_TORGTS
    );
  DOUT_0_OUTMUX_136 : X_BUF
    port map (
      I => rx_output_DOUT_0_OBUF,
      O => DOUT_0_OUTMUX
    );
  DOUT_0_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(0),
      O => DOUT_0_OD
    );
  rx_input_fifo_fifo_BU142 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1584,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1598_FFY_RST,
      O => rx_input_fifo_fifo_N1598
    );
  rx_input_fifo_fifo_N1598_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1598_FFY_RST
    );
  rx_output_DOUT_1_OBUF_137 : X_TRI
    port map (
      I => DOUT_1_OUTMUX,
      CTL => DOUT_1_ENABLE,
      O => DOUT(1)
    );
  DOUT_1_ENABLEINV : X_INV
    port map (
      I => DOUT_1_TORGTS,
      O => DOUT_1_ENABLE
    );
  DOUT_1_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_1_TORGTS
    );
  DOUT_1_OUTMUX_138 : X_BUF
    port map (
      I => rx_output_DOUT_1_OBUF,
      O => DOUT_1_OUTMUX
    );
  DOUT_1_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(1),
      O => DOUT_1_OD
    );
  rx_output_DOUT_2_OBUF_139 : X_TRI
    port map (
      I => DOUT_2_OUTMUX,
      CTL => DOUT_2_ENABLE,
      O => DOUT(2)
    );
  DOUT_2_ENABLEINV : X_INV
    port map (
      I => DOUT_2_TORGTS,
      O => DOUT_2_ENABLE
    );
  DOUT_2_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_2_TORGTS
    );
  DOUT_2_OUTMUX_140 : X_BUF
    port map (
      I => rx_output_DOUT_2_OBUF,
      O => DOUT_2_OUTMUX
    );
  DOUT_2_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(2),
      O => DOUT_2_OD
    );
  rx_output_DOUT_3_OBUF_141 : X_TRI
    port map (
      I => DOUT_3_OUTMUX,
      CTL => DOUT_3_ENABLE,
      O => DOUT(3)
    );
  DOUT_3_ENABLEINV : X_INV
    port map (
      I => DOUT_3_TORGTS,
      O => DOUT_3_ENABLE
    );
  DOUT_3_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_3_TORGTS
    );
  DOUT_3_OUTMUX_142 : X_BUF
    port map (
      I => rx_output_DOUT_3_OBUF,
      O => DOUT_3_OUTMUX
    );
  DOUT_3_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(3),
      O => DOUT_3_OD
    );
  rx_output_DOUT_4_OBUF_143 : X_TRI
    port map (
      I => DOUT_4_OUTMUX,
      CTL => DOUT_4_ENABLE,
      O => DOUT(4)
    );
  DOUT_4_ENABLEINV : X_INV
    port map (
      I => DOUT_4_TORGTS,
      O => DOUT_4_ENABLE
    );
  DOUT_4_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_4_TORGTS
    );
  DOUT_4_OUTMUX_144 : X_BUF
    port map (
      I => rx_output_DOUT_4_OBUF,
      O => DOUT_4_OUTMUX
    );
  DOUT_4_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(4),
      O => DOUT_4_OD
    );
  rx_output_DOUT_5_OBUF_145 : X_TRI
    port map (
      I => DOUT_5_OUTMUX,
      CTL => DOUT_5_ENABLE,
      O => DOUT(5)
    );
  DOUT_5_ENABLEINV : X_INV
    port map (
      I => DOUT_5_TORGTS,
      O => DOUT_5_ENABLE
    );
  DOUT_5_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_5_TORGTS
    );
  DOUT_5_OUTMUX_146 : X_BUF
    port map (
      I => rx_output_DOUT_5_OBUF,
      O => DOUT_5_OUTMUX
    );
  DOUT_5_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(5),
      O => DOUT_5_OD
    );
  rx_output_DOUT_6_OBUF_147 : X_TRI
    port map (
      I => DOUT_6_OUTMUX,
      CTL => DOUT_6_ENABLE,
      O => DOUT(6)
    );
  DOUT_6_ENABLEINV : X_INV
    port map (
      I => DOUT_6_TORGTS,
      O => DOUT_6_ENABLE
    );
  DOUT_6_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_6_TORGTS
    );
  DOUT_6_OUTMUX_148 : X_BUF
    port map (
      I => rx_output_DOUT_6_OBUF,
      O => DOUT_6_OUTMUX
    );
  DOUT_6_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(6),
      O => DOUT_6_OD
    );
  rx_output_DOUT_7_OBUF_149 : X_TRI
    port map (
      I => DOUT_7_OUTMUX,
      CTL => DOUT_7_ENABLE,
      O => DOUT(7)
    );
  DOUT_7_ENABLEINV : X_INV
    port map (
      I => DOUT_7_TORGTS,
      O => DOUT_7_ENABLE
    );
  DOUT_7_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_7_TORGTS
    );
  DOUT_7_OUTMUX_150 : X_BUF
    port map (
      I => rx_output_DOUT_7_OBUF,
      O => DOUT_7_OUTMUX
    );
  DOUT_7_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(7),
      O => DOUT_7_OD
    );
  rx_output_DOUT_8_OBUF_151 : X_TRI
    port map (
      I => DOUT_8_OUTMUX,
      CTL => DOUT_8_ENABLE,
      O => DOUT(8)
    );
  DOUT_8_ENABLEINV : X_INV
    port map (
      I => DOUT_8_TORGTS,
      O => DOUT_8_ENABLE
    );
  DOUT_8_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_8_TORGTS
    );
  DOUT_8_OUTMUX_152 : X_BUF
    port map (
      I => rx_output_DOUT_8_OBUF,
      O => DOUT_8_OUTMUX
    );
  DOUT_8_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(8),
      O => DOUT_8_OD
    );
  rx_output_DOUT_9_OBUF_153 : X_TRI
    port map (
      I => DOUT_9_OUTMUX,
      CTL => DOUT_9_ENABLE,
      O => DOUT(9)
    );
  DOUT_9_ENABLEINV : X_INV
    port map (
      I => DOUT_9_TORGTS,
      O => DOUT_9_ENABLE
    );
  DOUT_9_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => DOUT_9_TORGTS
    );
  DOUT_9_OUTMUX_154 : X_BUF
    port map (
      I => rx_output_DOUT_9_OBUF,
      O => DOUT_9_OUTMUX
    );
  DOUT_9_OMUX : X_BUF
    port map (
      I => rx_output_fifodout(9),
      O => DOUT_9_OD
    );
  mac_control_SOUT_OBUF_155 : X_TRI
    port map (
      I => SOUT_OUTMUX,
      CTL => SOUT_ENABLE,
      O => SOUT
    );
  SOUT_ENABLEINV : X_INV
    port map (
      I => SOUT_TORGTS,
      O => SOUT_ENABLE
    );
  SOUT_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => SOUT_TORGTS
    );
  SOUT_OUTMUX_156 : X_BUF
    port map (
      I => mac_control_SOUT_OBUF,
      O => SOUT_OUTMUX
    );
  SOUT_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => SOUT_OCEMUXNOT
    );
  SOUT_OMUX : X_BUF
    port map (
      I => mac_control_dout(31),
      O => SOUT_OD
    );
  SCLK_ICEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => SCLK_ICEMUXNOT
    );
  mac_control_SCLK_IBUF_157 : X_BUF
    port map (
      I => SCLK,
      O => mac_control_SCLK_IBUF
    );
  SCLK_DELAY : X_BUF
    port map (
      I => mac_control_SCLK_IBUF,
      O => SCLK_IDELAY
    );
  mac_control_LEDRX_OBUF_158 : X_TRI
    port map (
      I => LEDRX_OUTMUX,
      CTL => LEDRX_ENABLE,
      O => LEDRX
    );
  LEDRX_ENABLEINV : X_INV
    port map (
      I => LEDRX_TORGTS,
      O => LEDRX_ENABLE
    );
  LEDRX_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDRX_TORGTS
    );
  LEDRX_OUTMUX_159 : X_BUF
    port map (
      I => mac_control_LEDRX_OBUF,
      O => LEDRX_OUTMUX
    );
  LEDRX_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => LEDRX_OCEMUXNOT
    );
  LEDRX_OMUX : X_BUF
    port map (
      I => mac_control_n0040,
      O => LEDRX_OD
    );
  mac_control_LEDTX_OBUF_160 : X_TRI
    port map (
      I => LEDTX_OUTMUX,
      CTL => LEDTX_ENABLE,
      O => LEDTX
    );
  LEDTX_ENABLEINV : X_INV
    port map (
      I => LEDTX_TORGTS,
      O => LEDTX_ENABLE
    );
  LEDTX_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => LEDTX_TORGTS
    );
  LEDTX_OUTMUX_161 : X_BUF
    port map (
      I => mac_control_LEDTX_OBUF,
      O => LEDTX_OUTMUX
    );
  LEDTX_OCEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => LEDTX_OCEMUXNOT
    );
  LEDTX_OMUX : X_BUF
    port map (
      I => mac_control_n0038,
      O => LEDTX_OD
    );
  tx_input_DIN_0_IBUF_162 : X_BUF
    port map (
      I => DIN(0),
      O => tx_input_DIN_0_IBUF
    );
  tx_input_DIN_1_IBUF_163 : X_BUF
    port map (
      I => DIN(1),
      O => tx_input_DIN_1_IBUF
    );
  tx_input_DIN_2_IBUF_164 : X_BUF
    port map (
      I => DIN(2),
      O => tx_input_DIN_2_IBUF
    );
  tx_input_DIN_3_IBUF_165 : X_BUF
    port map (
      I => DIN(3),
      O => tx_input_DIN_3_IBUF
    );
  tx_input_DIN_4_IBUF_166 : X_BUF
    port map (
      I => DIN(4),
      O => tx_input_DIN_4_IBUF
    );
  tx_input_DIN_5_IBUF_167 : X_BUF
    port map (
      I => DIN(5),
      O => tx_input_DIN_5_IBUF
    );
  tx_input_DIN_6_IBUF_168 : X_BUF
    port map (
      I => DIN(6),
      O => tx_input_DIN_6_IBUF
    );
  tx_input_DIN_7_IBUF_169 : X_BUF
    port map (
      I => DIN(7),
      O => tx_input_DIN_7_IBUF
    );
  tx_input_DIN_8_IBUF_170 : X_BUF
    port map (
      I => DIN(8),
      O => tx_input_DIN_8_IBUF
    );
  tx_input_DIN_9_IBUF_171 : X_BUF
    port map (
      I => DIN(9),
      O => tx_input_DIN_9_IBUF
    );
  rx_input_GMII_RX_ER_IBUF_172 : X_BUF
    port map (
      I => RX_ER,
      O => rx_input_GMII_RX_ER_IBUF
    );
  rx_input_GMII_RX_DV_IBUF_173 : X_BUF
    port map (
      I => RX_DV,
      O => rx_input_GMII_RX_DV_IBUF
    );
  memcontroller_addrout10 : X_TRI
    port map (
      I => MA_10_OUTMUX,
      CTL => MA_10_ENABLE,
      O => MA(10)
    );
  MA_10_ENABLEINV : X_INV
    port map (
      I => MA_10_TORGTS,
      O => MA_10_ENABLE
    );
  MA_10_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_10_TORGTS
    );
  MA_10_OUTMUX_174 : X_BUF
    port map (
      I => memcontroller_addr(10),
      O => MA_10_OUTMUX
    );
  MA_10_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(10),
      O => MA_10_OD
    );
  rx_input_fifo_fifo_BU85 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N2172,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N1530_FFX_RST,
      O => rx_input_fifo_fifo_N1530
    );
  rx_input_fifo_fifo_N1530_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1530_FFX_RST
    );
  memcontroller_addrout11 : X_TRI
    port map (
      I => MA_11_OUTMUX,
      CTL => MA_11_ENABLE,
      O => MA(11)
    );
  MA_11_ENABLEINV : X_INV
    port map (
      I => MA_11_TORGTS,
      O => MA_11_ENABLE
    );
  MA_11_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_11_TORGTS
    );
  MA_11_OUTMUX_175 : X_BUF
    port map (
      I => memcontroller_addr(11),
      O => MA_11_OUTMUX
    );
  MA_11_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(11),
      O => MA_11_OD
    );
  memcontroller_addrout12 : X_TRI
    port map (
      I => MA_12_OUTMUX,
      CTL => MA_12_ENABLE,
      O => MA(12)
    );
  MA_12_ENABLEINV : X_INV
    port map (
      I => MA_12_TORGTS,
      O => MA_12_ENABLE
    );
  MA_12_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_12_TORGTS
    );
  MA_12_OUTMUX_176 : X_BUF
    port map (
      I => memcontroller_addr(12),
      O => MA_12_OUTMUX
    );
  MA_12_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(12),
      O => MA_12_OD
    );
  memcontroller_addrout13 : X_TRI
    port map (
      I => MA_13_OUTMUX,
      CTL => MA_13_ENABLE,
      O => MA(13)
    );
  MA_13_ENABLEINV : X_INV
    port map (
      I => MA_13_TORGTS,
      O => MA_13_ENABLE
    );
  MA_13_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_13_TORGTS
    );
  MA_13_OUTMUX_177 : X_BUF
    port map (
      I => memcontroller_addr(13),
      O => MA_13_OUTMUX
    );
  MA_13_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(13),
      O => MA_13_OD
    );
  memcontroller_addrout14 : X_TRI
    port map (
      I => MA_14_OUTMUX,
      CTL => MA_14_ENABLE,
      O => MA(14)
    );
  MA_14_ENABLEINV : X_INV
    port map (
      I => MA_14_TORGTS,
      O => MA_14_ENABLE
    );
  MA_14_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_14_TORGTS
    );
  MA_14_OUTMUX_178 : X_BUF
    port map (
      I => memcontroller_addr(14),
      O => MA_14_OUTMUX
    );
  MA_14_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(14),
      O => MA_14_OD
    );
  memcontroller_addrout15 : X_TRI
    port map (
      I => MA_15_OUTMUX,
      CTL => MA_15_ENABLE,
      O => MA(15)
    );
  MA_15_ENABLEINV : X_INV
    port map (
      I => MA_15_TORGTS,
      O => MA_15_ENABLE
    );
  MA_15_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_15_TORGTS
    );
  MA_15_OUTMUX_179 : X_BUF
    port map (
      I => memcontroller_addr(15),
      O => MA_15_OUTMUX
    );
  MA_15_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(15),
      O => MA_15_OD
    );
  memcontroller_addrout16 : X_TRI
    port map (
      I => MA_16_OUTMUX,
      CTL => MA_16_ENABLE,
      O => MA(16)
    );
  MA_16_ENABLEINV : X_INV
    port map (
      I => MA_16_TORGTS,
      O => MA_16_ENABLE
    );
  MA_16_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_16_TORGTS
    );
  MA_16_OUTMUX_180 : X_BUF
    port map (
      I => memcontroller_addr(16),
      O => MA_16_OUTMUX
    );
  MA_16_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(16),
      O => MA_16_OD
    );
  memcontroller_qdout10_OBUFT : X_TRI
    port map (
      I => MD_10_OUTMUX,
      CTL => MD_10_ENABLE,
      O => MD(10)
    );
  MD_10_ENABLEINV : X_INV
    port map (
      I => MD_10_TORGTS,
      O => MD_10_ENABLE
    );
  MD_10_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_10_TORGTS
    );
  MD_10_OUTMUX_181 : X_BUF
    port map (
      I => memcontroller_dnout(10),
      O => MD_10_OUTMUX
    );
  MD_10_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(10),
      O => MD_10_OD
    );
  memcontroller_qdout10_IBUF : X_BUF
    port map (
      I => MD(10),
      O => memcontroller_q(10)
    );
  memcontroller_qdout11_OBUFT : X_TRI
    port map (
      I => MD_11_OUTMUX,
      CTL => MD_11_ENABLE,
      O => MD(11)
    );
  MD_11_ENABLEINV : X_INV
    port map (
      I => MD_11_TORGTS,
      O => MD_11_ENABLE
    );
  MD_11_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_11_TORGTS
    );
  MD_11_OUTMUX_182 : X_BUF
    port map (
      I => memcontroller_dnout(11),
      O => MD_11_OUTMUX
    );
  MD_11_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(11),
      O => MD_11_OD
    );
  memcontroller_qdout11_IBUF : X_BUF
    port map (
      I => MD(11),
      O => memcontroller_q(11)
    );
  rx_input_fifo_fifo_BU133 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_fifo_N1586,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => rx_input_fifo_fifo_N1599_FFY_SET,
      RST => GND,
      O => rx_input_fifo_fifo_N1600
    );
  rx_input_fifo_fifo_N1599_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_fifo_RESET_1,
      O => rx_input_fifo_fifo_N1599_FFY_SET
    );
  memcontroller_qdout20_OBUFT : X_TRI
    port map (
      I => MD_20_OUTMUX,
      CTL => MD_20_ENABLE,
      O => MD(20)
    );
  MD_20_ENABLEINV : X_INV
    port map (
      I => MD_20_TORGTS,
      O => MD_20_ENABLE
    );
  MD_20_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_20_TORGTS
    );
  MD_20_OUTMUX_183 : X_BUF
    port map (
      I => memcontroller_dnout(20),
      O => MD_20_OUTMUX
    );
  MD_20_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(20),
      O => MD_20_OD
    );
  memcontroller_qdout20_IBUF : X_BUF
    port map (
      I => MD(20),
      O => memcontroller_q(20)
    );
  memcontroller_qdout12_OBUFT : X_TRI
    port map (
      I => MD_12_OUTMUX,
      CTL => MD_12_ENABLE,
      O => MD(12)
    );
  MD_12_ENABLEINV : X_INV
    port map (
      I => MD_12_TORGTS,
      O => MD_12_ENABLE
    );
  MD_12_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_12_TORGTS
    );
  MD_12_OUTMUX_184 : X_BUF
    port map (
      I => memcontroller_dnout(12),
      O => MD_12_OUTMUX
    );
  MD_12_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(12),
      O => MD_12_OD
    );
  memcontroller_qdout12_IBUF : X_BUF
    port map (
      I => MD(12),
      O => memcontroller_q(12)
    );
  memcontroller_qdout21_OBUFT : X_TRI
    port map (
      I => MD_21_OUTMUX,
      CTL => MD_21_ENABLE,
      O => MD(21)
    );
  MD_21_ENABLEINV : X_INV
    port map (
      I => MD_21_TORGTS,
      O => MD_21_ENABLE
    );
  MD_21_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_21_TORGTS
    );
  MD_21_OUTMUX_185 : X_BUF
    port map (
      I => memcontroller_dnout(21),
      O => MD_21_OUTMUX
    );
  MD_21_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(21),
      O => MD_21_OD
    );
  memcontroller_qdout21_IBUF : X_BUF
    port map (
      I => MD(21),
      O => memcontroller_q(21)
    );
  memcontroller_qdout13_OBUFT : X_TRI
    port map (
      I => MD_13_OUTMUX,
      CTL => MD_13_ENABLE,
      O => MD(13)
    );
  MD_13_ENABLEINV : X_INV
    port map (
      I => MD_13_TORGTS,
      O => MD_13_ENABLE
    );
  MD_13_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_13_TORGTS
    );
  MD_13_OUTMUX_186 : X_BUF
    port map (
      I => memcontroller_dnout(13),
      O => MD_13_OUTMUX
    );
  MD_13_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(13),
      O => MD_13_OD
    );
  memcontroller_qdout13_IBUF : X_BUF
    port map (
      I => MD(13),
      O => memcontroller_q(13)
    );
  memcontroller_qdout22_OBUFT : X_TRI
    port map (
      I => MD_22_OUTMUX,
      CTL => MD_22_ENABLE,
      O => MD(22)
    );
  MD_22_ENABLEINV : X_INV
    port map (
      I => MD_22_TORGTS,
      O => MD_22_ENABLE
    );
  MD_22_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_22_TORGTS
    );
  MD_22_OUTMUX_187 : X_BUF
    port map (
      I => memcontroller_dnout(22),
      O => MD_22_OUTMUX
    );
  MD_22_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(22),
      O => MD_22_OD
    );
  memcontroller_qdout22_IBUF : X_BUF
    port map (
      I => MD(22),
      O => memcontroller_q(22)
    );
  memcontroller_qdout14_OBUFT : X_TRI
    port map (
      I => MD_14_OUTMUX,
      CTL => MD_14_ENABLE,
      O => MD(14)
    );
  MD_14_ENABLEINV : X_INV
    port map (
      I => MD_14_TORGTS,
      O => MD_14_ENABLE
    );
  MD_14_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_14_TORGTS
    );
  MD_14_OUTMUX_188 : X_BUF
    port map (
      I => memcontroller_dnout(14),
      O => MD_14_OUTMUX
    );
  MD_14_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(14),
      O => MD_14_OD
    );
  memcontroller_qdout14_IBUF : X_BUF
    port map (
      I => MD(14),
      O => memcontroller_q(14)
    );
  memcontroller_qdout30_OBUFT : X_TRI
    port map (
      I => MD_30_OUTMUX,
      CTL => MD_30_ENABLE,
      O => MD(30)
    );
  MD_30_ENABLEINV : X_INV
    port map (
      I => MD_30_TORGTS,
      O => MD_30_ENABLE
    );
  MD_30_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_30_TORGTS
    );
  MD_30_OUTMUX_189 : X_BUF
    port map (
      I => memcontroller_dnout(30),
      O => MD_30_OUTMUX
    );
  MD_30_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(30),
      O => MD_30_OD
    );
  memcontroller_qdout30_IBUF : X_BUF
    port map (
      I => MD(30),
      O => memcontroller_q(30)
    );
  rx_input_fifo_fifo_BU47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1858,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N15_FFY_RST,
      O => rx_input_fifo_fifo_N14
    );
  rx_input_fifo_fifo_N15_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N15_FFY_RST
    );
  memcontroller_qdout23_OBUFT : X_TRI
    port map (
      I => MD_23_OUTMUX,
      CTL => MD_23_ENABLE,
      O => MD(23)
    );
  MD_23_ENABLEINV : X_INV
    port map (
      I => MD_23_TORGTS,
      O => MD_23_ENABLE
    );
  MD_23_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_23_TORGTS
    );
  MD_23_OUTMUX_190 : X_BUF
    port map (
      I => memcontroller_dnout(23),
      O => MD_23_OUTMUX
    );
  MD_23_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(23),
      O => MD_23_OD
    );
  memcontroller_qdout23_IBUF : X_BUF
    port map (
      I => MD(23),
      O => memcontroller_q(23)
    );
  memcontroller_qdout15_OBUFT : X_TRI
    port map (
      I => MD_15_OUTMUX,
      CTL => MD_15_ENABLE,
      O => MD(15)
    );
  MD_15_ENABLEINV : X_INV
    port map (
      I => MD_15_TORGTS,
      O => MD_15_ENABLE
    );
  MD_15_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_15_TORGTS
    );
  MD_15_OUTMUX_191 : X_BUF
    port map (
      I => memcontroller_dnout(15),
      O => MD_15_OUTMUX
    );
  MD_15_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(15),
      O => MD_15_OD
    );
  memcontroller_qdout15_IBUF : X_BUF
    port map (
      I => MD(15),
      O => memcontroller_q(15)
    );
  memcontroller_qdout31_OBUFT : X_TRI
    port map (
      I => MD_31_OUTMUX,
      CTL => MD_31_ENABLE,
      O => MD(31)
    );
  MD_31_ENABLEINV : X_INV
    port map (
      I => MD_31_TORGTS,
      O => MD_31_ENABLE
    );
  MD_31_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_31_TORGTS
    );
  MD_31_OUTMUX_192 : X_BUF
    port map (
      I => memcontroller_dnout(31),
      O => MD_31_OUTMUX
    );
  MD_31_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(31),
      O => MD_31_OD
    );
  memcontroller_qdout31_IBUF : X_BUF
    port map (
      I => MD(31),
      O => memcontroller_q(31)
    );
  memcontroller_qdout24_OBUFT : X_TRI
    port map (
      I => MD_24_OUTMUX,
      CTL => MD_24_ENABLE,
      O => MD(24)
    );
  MD_24_ENABLEINV : X_INV
    port map (
      I => MD_24_TORGTS,
      O => MD_24_ENABLE
    );
  MD_24_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_24_TORGTS
    );
  MD_24_OUTMUX_193 : X_BUF
    port map (
      I => memcontroller_dnout(24),
      O => MD_24_OUTMUX
    );
  MD_24_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(24),
      O => MD_24_OD
    );
  memcontroller_qdout24_IBUF : X_BUF
    port map (
      I => MD(24),
      O => memcontroller_q(24)
    );
  memcontroller_qdout16_OBUFT : X_TRI
    port map (
      I => MD_16_OUTMUX,
      CTL => MD_16_ENABLE,
      O => MD(16)
    );
  MD_16_ENABLEINV : X_INV
    port map (
      I => MD_16_TORGTS,
      O => MD_16_ENABLE
    );
  MD_16_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_16_TORGTS
    );
  MD_16_OUTMUX_194 : X_BUF
    port map (
      I => memcontroller_dnout(16),
      O => MD_16_OUTMUX
    );
  MD_16_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(16),
      O => MD_16_OD
    );
  memcontroller_qdout16_IBUF : X_BUF
    port map (
      I => MD(16),
      O => memcontroller_q(16)
    );
  memcontroller_qdout17_OBUFT : X_TRI
    port map (
      I => MD_17_OUTMUX,
      CTL => MD_17_ENABLE,
      O => MD(17)
    );
  MD_17_ENABLEINV : X_INV
    port map (
      I => MD_17_TORGTS,
      O => MD_17_ENABLE
    );
  MD_17_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_17_TORGTS
    );
  MD_17_OUTMUX_195 : X_BUF
    port map (
      I => memcontroller_dnout(17),
      O => MD_17_OUTMUX
    );
  MD_17_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(17),
      O => MD_17_OD
    );
  memcontroller_qdout17_IBUF : X_BUF
    port map (
      I => MD(17),
      O => memcontroller_q(17)
    );
  memcontroller_qdout25_OBUFT : X_TRI
    port map (
      I => MD_25_OUTMUX,
      CTL => MD_25_ENABLE,
      O => MD(25)
    );
  MD_25_ENABLEINV : X_INV
    port map (
      I => MD_25_TORGTS,
      O => MD_25_ENABLE
    );
  MD_25_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_25_TORGTS
    );
  MD_25_OUTMUX_196 : X_BUF
    port map (
      I => memcontroller_dnout(25),
      O => MD_25_OUTMUX
    );
  MD_25_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(25),
      O => MD_25_OD
    );
  memcontroller_qdout25_IBUF : X_BUF
    port map (
      I => MD(25),
      O => memcontroller_q(25)
    );
  memcontroller_qdout18_OBUFT : X_TRI
    port map (
      I => MD_18_OUTMUX,
      CTL => MD_18_ENABLE,
      O => MD(18)
    );
  MD_18_ENABLEINV : X_INV
    port map (
      I => MD_18_TORGTS,
      O => MD_18_ENABLE
    );
  MD_18_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_18_TORGTS
    );
  MD_18_OUTMUX_197 : X_BUF
    port map (
      I => memcontroller_dnout(18),
      O => MD_18_OUTMUX
    );
  MD_18_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(18),
      O => MD_18_OD
    );
  memcontroller_qdout18_IBUF : X_BUF
    port map (
      I => MD(18),
      O => memcontroller_q(18)
    );
  memcontroller_qdout26_OBUFT : X_TRI
    port map (
      I => MD_26_OUTMUX,
      CTL => MD_26_ENABLE,
      O => MD(26)
    );
  MD_26_ENABLEINV : X_INV
    port map (
      I => MD_26_TORGTS,
      O => MD_26_ENABLE
    );
  MD_26_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_26_TORGTS
    );
  MD_26_OUTMUX_198 : X_BUF
    port map (
      I => memcontroller_dnout(26),
      O => MD_26_OUTMUX
    );
  MD_26_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(26),
      O => MD_26_OD
    );
  memcontroller_qdout26_IBUF : X_BUF
    port map (
      I => MD(26),
      O => memcontroller_q(26)
    );
  memcontroller_qdout19_OBUFT : X_TRI
    port map (
      I => MD_19_OUTMUX,
      CTL => MD_19_ENABLE,
      O => MD(19)
    );
  MD_19_ENABLEINV : X_INV
    port map (
      I => MD_19_TORGTS,
      O => MD_19_ENABLE
    );
  MD_19_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_19_TORGTS
    );
  MD_19_OUTMUX_199 : X_BUF
    port map (
      I => memcontroller_dnout(19),
      O => MD_19_OUTMUX
    );
  MD_19_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(19),
      O => MD_19_OD
    );
  memcontroller_qdout19_IBUF : X_BUF
    port map (
      I => MD(19),
      O => memcontroller_q(19)
    );
  memcontroller_qdout27_OBUFT : X_TRI
    port map (
      I => MD_27_OUTMUX,
      CTL => MD_27_ENABLE,
      O => MD(27)
    );
  MD_27_ENABLEINV : X_INV
    port map (
      I => MD_27_TORGTS,
      O => MD_27_ENABLE
    );
  MD_27_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_27_TORGTS
    );
  MD_27_OUTMUX_200 : X_BUF
    port map (
      I => memcontroller_dnout(27),
      O => MD_27_OUTMUX
    );
  MD_27_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(27),
      O => MD_27_OD
    );
  memcontroller_qdout27_IBUF : X_BUF
    port map (
      I => MD(27),
      O => memcontroller_q(27)
    );
  memcontroller_qdout28_OBUFT : X_TRI
    port map (
      I => MD_28_OUTMUX,
      CTL => MD_28_ENABLE,
      O => MD(28)
    );
  MD_28_ENABLEINV : X_INV
    port map (
      I => MD_28_TORGTS,
      O => MD_28_ENABLE
    );
  MD_28_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_28_TORGTS
    );
  MD_28_OUTMUX_201 : X_BUF
    port map (
      I => memcontroller_dnout(28),
      O => MD_28_OUTMUX
    );
  MD_28_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(28),
      O => MD_28_OD
    );
  memcontroller_qdout28_IBUF : X_BUF
    port map (
      I => MD(28),
      O => memcontroller_q(28)
    );
  memcontroller_qdout29_OBUFT : X_TRI
    port map (
      I => MD_29_OUTMUX,
      CTL => MD_29_ENABLE,
      O => MD(29)
    );
  MD_29_ENABLEINV : X_INV
    port map (
      I => MD_29_TORGTS,
      O => MD_29_ENABLE
    );
  MD_29_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_29_TORGTS
    );
  MD_29_OUTMUX_202 : X_BUF
    port map (
      I => memcontroller_dnout(29),
      O => MD_29_OUTMUX
    );
  MD_29_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(29),
      O => MD_29_OD
    );
  memcontroller_qdout29_IBUF : X_BUF
    port map (
      I => MD(29),
      O => memcontroller_q(29)
    );
  memcontroller_addrout0 : X_TRI
    port map (
      I => MA_0_OUTMUX,
      CTL => MA_0_ENABLE,
      O => MA(0)
    );
  MA_0_ENABLEINV : X_INV
    port map (
      I => MA_0_TORGTS,
      O => MA_0_ENABLE
    );
  MA_0_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_0_TORGTS
    );
  MA_0_OUTMUX_203 : X_BUF
    port map (
      I => memcontroller_addr(0),
      O => MA_0_OUTMUX
    );
  MA_0_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(0),
      O => MA_0_OD
    );
  memcontroller_addrout1 : X_TRI
    port map (
      I => MA_1_OUTMUX,
      CTL => MA_1_ENABLE,
      O => MA(1)
    );
  MA_1_ENABLEINV : X_INV
    port map (
      I => MA_1_TORGTS,
      O => MA_1_ENABLE
    );
  MA_1_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_1_TORGTS
    );
  MA_1_OUTMUX_204 : X_BUF
    port map (
      I => memcontroller_addr(1),
      O => MA_1_OUTMUX
    );
  MA_1_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(1),
      O => MA_1_OD
    );
  memcontroller_addrout2 : X_TRI
    port map (
      I => MA_2_OUTMUX,
      CTL => MA_2_ENABLE,
      O => MA(2)
    );
  MA_2_ENABLEINV : X_INV
    port map (
      I => MA_2_TORGTS,
      O => MA_2_ENABLE
    );
  MA_2_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_2_TORGTS
    );
  MA_2_OUTMUX_205 : X_BUF
    port map (
      I => memcontroller_addr(2),
      O => MA_2_OUTMUX
    );
  MA_2_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(2),
      O => MA_2_OD
    );
  memcontroller_addrout3 : X_TRI
    port map (
      I => MA_3_OUTMUX,
      CTL => MA_3_ENABLE,
      O => MA(3)
    );
  MA_3_ENABLEINV : X_INV
    port map (
      I => MA_3_TORGTS,
      O => MA_3_ENABLE
    );
  MA_3_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_3_TORGTS
    );
  MA_3_OUTMUX_206 : X_BUF
    port map (
      I => memcontroller_addr(3),
      O => MA_3_OUTMUX
    );
  MA_3_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(3),
      O => MA_3_OD
    );
  memcontroller_addrout4 : X_TRI
    port map (
      I => MA_4_OUTMUX,
      CTL => MA_4_ENABLE,
      O => MA(4)
    );
  MA_4_ENABLEINV : X_INV
    port map (
      I => MA_4_TORGTS,
      O => MA_4_ENABLE
    );
  MA_4_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_4_TORGTS
    );
  MA_4_OUTMUX_207 : X_BUF
    port map (
      I => memcontroller_addr(4),
      O => MA_4_OUTMUX
    );
  MA_4_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(4),
      O => MA_4_OD
    );
  memcontroller_addrout5 : X_TRI
    port map (
      I => MA_5_OUTMUX,
      CTL => MA_5_ENABLE,
      O => MA(5)
    );
  MA_5_ENABLEINV : X_INV
    port map (
      I => MA_5_TORGTS,
      O => MA_5_ENABLE
    );
  MA_5_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_5_TORGTS
    );
  MA_5_OUTMUX_208 : X_BUF
    port map (
      I => memcontroller_addr(5),
      O => MA_5_OUTMUX
    );
  MA_5_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(5),
      O => MA_5_OD
    );
  memcontroller_addrout6 : X_TRI
    port map (
      I => MA_6_OUTMUX,
      CTL => MA_6_ENABLE,
      O => MA(6)
    );
  MA_6_ENABLEINV : X_INV
    port map (
      I => MA_6_TORGTS,
      O => MA_6_ENABLE
    );
  MA_6_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_6_TORGTS
    );
  MA_6_OUTMUX_209 : X_BUF
    port map (
      I => memcontroller_addr(6),
      O => MA_6_OUTMUX
    );
  MA_6_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(6),
      O => MA_6_OD
    );
  memcontroller_addrout7 : X_TRI
    port map (
      I => MA_7_OUTMUX,
      CTL => MA_7_ENABLE,
      O => MA(7)
    );
  MA_7_ENABLEINV : X_INV
    port map (
      I => MA_7_TORGTS,
      O => MA_7_ENABLE
    );
  MA_7_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_7_TORGTS
    );
  MA_7_OUTMUX_210 : X_BUF
    port map (
      I => memcontroller_addr(7),
      O => MA_7_OUTMUX
    );
  MA_7_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(7),
      O => MA_7_OD
    );
  memcontroller_addrout8 : X_TRI
    port map (
      I => MA_8_OUTMUX,
      CTL => MA_8_ENABLE,
      O => MA(8)
    );
  MA_8_ENABLEINV : X_INV
    port map (
      I => MA_8_TORGTS,
      O => MA_8_ENABLE
    );
  MA_8_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_8_TORGTS
    );
  MA_8_OUTMUX_211 : X_BUF
    port map (
      I => memcontroller_addr(8),
      O => MA_8_OUTMUX
    );
  MA_8_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(8),
      O => MA_8_OD
    );
  mac_control_phyaddr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_9_FFY_RST,
      O => mac_control_phyaddr(8)
    );
  mac_control_phyaddr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_9_FFY_RST
    );
  memcontroller_addrout9 : X_TRI
    port map (
      I => MA_9_OUTMUX,
      CTL => MA_9_ENABLE,
      O => MA(9)
    );
  MA_9_ENABLEINV : X_INV
    port map (
      I => MA_9_TORGTS,
      O => MA_9_ENABLE
    );
  MA_9_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => MA_9_TORGTS
    );
  MA_9_OUTMUX_212 : X_BUF
    port map (
      I => memcontroller_addr(9),
      O => MA_9_OUTMUX
    );
  MA_9_OMUX : X_BUF
    port map (
      I => memcontroller_addrn(9),
      O => MA_9_OD
    );
  mac_control_PHYRESET_OBUF_213 : X_TRI
    port map (
      I => PHYRESET_OUTMUX,
      CTL => PHYRESET_ENABLE,
      O => PHYRESET
    );
  PHYRESET_ENABLEINV : X_INV
    port map (
      I => PHYRESET_TORGTS,
      O => PHYRESET_ENABLE
    );
  PHYRESET_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => PHYRESET_TORGTS
    );
  PHYRESET_OUTMUX_214 : X_BUF
    port map (
      I => mac_control_PHYRESET_OBUF,
      O => PHYRESET_OUTMUX
    );
  PHYRESET_OMUX : X_BUF
    port map (
      I => mac_control_n0034,
      O => PHYRESET_OD
    );
  memcontroller_qdout0_OBUFT : X_TRI
    port map (
      I => MD_0_OUTMUX,
      CTL => MD_0_ENABLE,
      O => MD(0)
    );
  MD_0_ENABLEINV : X_INV
    port map (
      I => MD_0_TORGTS,
      O => MD_0_ENABLE
    );
  MD_0_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_0_TORGTS
    );
  MD_0_OUTMUX_215 : X_BUF
    port map (
      I => memcontroller_dnout(0),
      O => MD_0_OUTMUX
    );
  MD_0_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(0),
      O => MD_0_OD
    );
  memcontroller_qdout0_IBUF : X_BUF
    port map (
      I => MD(0),
      O => memcontroller_q(0)
    );
  memcontroller_qdout1_OBUFT : X_TRI
    port map (
      I => MD_1_OUTMUX,
      CTL => MD_1_ENABLE,
      O => MD(1)
    );
  MD_1_ENABLEINV : X_INV
    port map (
      I => MD_1_TORGTS,
      O => MD_1_ENABLE
    );
  MD_1_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_1_TORGTS
    );
  MD_1_OUTMUX_216 : X_BUF
    port map (
      I => memcontroller_dnout(1),
      O => MD_1_OUTMUX
    );
  MD_1_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(1),
      O => MD_1_OD
    );
  memcontroller_qdout1_IBUF : X_BUF
    port map (
      I => MD(1),
      O => memcontroller_q(1)
    );
  rx_input_fifo_fifo_BU41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1857,
      CE => rx_input_fifo_fifo_N1495,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_fifo_N15_FFX_RST,
      O => rx_input_fifo_fifo_N15
    );
  rx_input_fifo_fifo_N15_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N15_FFX_RST
    );
  memcontroller_qdout2_OBUFT : X_TRI
    port map (
      I => MD_2_OUTMUX,
      CTL => MD_2_ENABLE,
      O => MD(2)
    );
  MD_2_ENABLEINV : X_INV
    port map (
      I => MD_2_TORGTS,
      O => MD_2_ENABLE
    );
  MD_2_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_2_TORGTS
    );
  MD_2_OUTMUX_217 : X_BUF
    port map (
      I => memcontroller_dnout(2),
      O => MD_2_OUTMUX
    );
  MD_2_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(2),
      O => MD_2_OD
    );
  memcontroller_qdout2_IBUF : X_BUF
    port map (
      I => MD(2),
      O => memcontroller_q(2)
    );
  memcontroller_qdout3_OBUFT : X_TRI
    port map (
      I => MD_3_OUTMUX,
      CTL => MD_3_ENABLE,
      O => MD(3)
    );
  MD_3_ENABLEINV : X_INV
    port map (
      I => MD_3_TORGTS,
      O => MD_3_ENABLE
    );
  MD_3_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_3_TORGTS
    );
  MD_3_OUTMUX_218 : X_BUF
    port map (
      I => memcontroller_dnout(3),
      O => MD_3_OUTMUX
    );
  MD_3_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(3),
      O => MD_3_OD
    );
  memcontroller_qdout3_IBUF : X_BUF
    port map (
      I => MD(3),
      O => memcontroller_q(3)
    );
  memcontroller_qdout4_OBUFT : X_TRI
    port map (
      I => MD_4_OUTMUX,
      CTL => MD_4_ENABLE,
      O => MD(4)
    );
  MD_4_ENABLEINV : X_INV
    port map (
      I => MD_4_TORGTS,
      O => MD_4_ENABLE
    );
  MD_4_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_4_TORGTS
    );
  MD_4_OUTMUX_219 : X_BUF
    port map (
      I => memcontroller_dnout(4),
      O => MD_4_OUTMUX
    );
  MD_4_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(4),
      O => MD_4_OD
    );
  memcontroller_qdout4_IBUF : X_BUF
    port map (
      I => MD(4),
      O => memcontroller_q(4)
    );
  memcontroller_qdout5_OBUFT : X_TRI
    port map (
      I => MD_5_OUTMUX,
      CTL => MD_5_ENABLE,
      O => MD(5)
    );
  MD_5_ENABLEINV : X_INV
    port map (
      I => MD_5_TORGTS,
      O => MD_5_ENABLE
    );
  MD_5_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_5_TORGTS
    );
  MD_5_OUTMUX_220 : X_BUF
    port map (
      I => memcontroller_dnout(5),
      O => MD_5_OUTMUX
    );
  MD_5_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(5),
      O => MD_5_OD
    );
  memcontroller_qdout5_IBUF : X_BUF
    port map (
      I => MD(5),
      O => memcontroller_q(5)
    );
  memcontroller_qdout6_OBUFT : X_TRI
    port map (
      I => MD_6_OUTMUX,
      CTL => MD_6_ENABLE,
      O => MD(6)
    );
  MD_6_ENABLEINV : X_INV
    port map (
      I => MD_6_TORGTS,
      O => MD_6_ENABLE
    );
  MD_6_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_6_TORGTS
    );
  MD_6_OUTMUX_221 : X_BUF
    port map (
      I => memcontroller_dnout(6),
      O => MD_6_OUTMUX
    );
  MD_6_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(6),
      O => MD_6_OD
    );
  memcontroller_qdout6_IBUF : X_BUF
    port map (
      I => MD(6),
      O => memcontroller_q(6)
    );
  memcontroller_qdout7_OBUFT : X_TRI
    port map (
      I => MD_7_OUTMUX,
      CTL => MD_7_ENABLE,
      O => MD(7)
    );
  MD_7_ENABLEINV : X_INV
    port map (
      I => MD_7_TORGTS,
      O => MD_7_ENABLE
    );
  MD_7_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_7_TORGTS
    );
  MD_7_OUTMUX_222 : X_BUF
    port map (
      I => memcontroller_dnout(7),
      O => MD_7_OUTMUX
    );
  MD_7_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(7),
      O => MD_7_OD
    );
  memcontroller_qdout7_IBUF : X_BUF
    port map (
      I => MD(7),
      O => memcontroller_q(7)
    );
  memcontroller_qdout8_OBUFT : X_TRI
    port map (
      I => MD_8_OUTMUX,
      CTL => MD_8_ENABLE,
      O => MD(8)
    );
  MD_8_ENABLEINV : X_INV
    port map (
      I => MD_8_TORGTS,
      O => MD_8_ENABLE
    );
  MD_8_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_8_TORGTS
    );
  MD_8_OUTMUX_223 : X_BUF
    port map (
      I => memcontroller_dnout(8),
      O => MD_8_OUTMUX
    );
  MD_8_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(8),
      O => MD_8_OD
    );
  memcontroller_qdout8_IBUF : X_BUF
    port map (
      I => MD(8),
      O => memcontroller_q(8)
    );
  memcontroller_qdout9_OBUFT : X_TRI
    port map (
      I => MD_9_OUTMUX,
      CTL => MD_9_ENABLE,
      O => MD(9)
    );
  MD_9_ENABLEINV : X_INV
    port map (
      I => MD_9_TORGTS,
      O => MD_9_ENABLE
    );
  MD_9_GTS_OR : X_OR2
    port map (
      I0 => GTS,
      I1 => memcontroller_ts(0),
      O => MD_9_TORGTS
    );
  MD_9_OUTMUX_224 : X_BUF
    port map (
      I => memcontroller_dnout(9),
      O => MD_9_OUTMUX
    );
  MD_9_OMUX : X_BUF
    port map (
      I => memcontroller_dnl2(9),
      O => MD_9_OD
    );
  memcontroller_qdout9_IBUF : X_BUF
    port map (
      I => MD(9),
      O => memcontroller_q(9)
    );
  GTX_CLK_OBUF_225 : X_TRI
    port map (
      I => GTX_CLK_OUTMUX,
      CTL => GTX_CLK_ENABLE,
      O => GTX_CLK
    );
  GTX_CLK_ENABLEINV : X_INV
    port map (
      I => GTX_CLK_TORGTS,
      O => GTX_CLK_ENABLE
    );
  GTX_CLK_GTS_OR : X_BUF
    port map (
      I => GTS,
      O => GTX_CLK_TORGTS
    );
  GTX_CLK_OUTMUX_226 : X_BUF
    port map (
      I => GTX_CLK_OBUF,
      O => GTX_CLK_OUTMUX
    );
  clkio_dll : X_CLKDLLE
    generic map(
      CLKDV_DIVIDE => 4.0,
      DUTY_CYCLE_CORRECTION => TRUE,
      MAXPERCLKIN => 40000 ps
    )
    port map (
      CLKIN => CLKIOIN_IBUFG,
      CLKFB => clkio,
      RST => RESET_IBUF,
      CLK0 => clkio_to_bufg,
      CLK90 => clkio_dll_CLK90,
      CLK180 => clkio_dll_CLK180,
      CLK270 => clkio_dll_CLK270,
      CLK2X => clkio_dll_CLK2X,
      CLK2X180 => clkio_dll_CLK2X180,
      CLKDV => clkio_dll_CLKDV,
      LOCKED => clkio_dll_LOCKED
    );
  clk_dll : X_CLKDLLE
    generic map(
      CLKDV_DIVIDE => 4.0,
      DUTY_CYCLE_CORRECTION => TRUE,
      MAXPERCLKIN => 40000 ps
    )
    port map (
      CLKIN => CLKIN_IBUFG,
      CLKFB => GTX_CLK_OBUF,
      RST => RESET_IBUF,
      CLK0 => clk_to_bufg,
      CLK90 => clk_dll_CLK90,
      CLK180 => clk_dll_CLK180,
      CLK270 => clk_dll_CLK270,
      CLK2X => clk_dll_CLK2X,
      CLK2X180 => clk_dll_CLK2X180,
      CLKDV => clksl,
      LOCKED => clk_dll_LOCKED
    );
  clkrx_dll : X_CLKDLLE
    generic map(
      CLKDV_DIVIDE => 4.0,
      DUTY_CYCLE_CORRECTION => TRUE,
      MAXPERCLKIN => 40000 ps
    )
    port map (
      CLKIN => RX_CLK_IBUFG,
      CLKFB => clkrx,
      RST => RESET_IBUF,
      CLK0 => clkrx_to_bufg,
      CLK90 => clkrx_dll_CLK90,
      CLK180 => clkrx_dll_CLK180,
      CLK270 => clkrx_dll_CLK270,
      CLK2X => clkrx_dll_CLK2X,
      CLK2X180 => clkrx_dll_CLK2X180,
      CLKDV => clkrx_dll_CLKDV,
      LOCKED => clkrx_dll_LOCKED
    );
  rx_input_fifo_fifo_B7_LOGIC_ONE_227 : X_ONE
    port map (
      O => rx_input_fifo_fifo_B7_LOGIC_ONE
    );
  rx_input_fifo_fifo_B7_LOGIC_ZERO_228 : X_ZERO
    port map (
      O => rx_input_fifo_fifo_B7_LOGIC_ZERO
    );
  rx_input_fifo_fifo_B7 : X_RAMB4_S16_S16
    generic map(
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      SETUP_ALL => 3025 ps,
      XON => FALSE
    )
    port map (
      CLKA => clkrx,
      CLKB => GTX_CLK_OBUF,
      ENA => rx_input_fifo_fifo_B7_LOGIC_ONE,
      ENB => rx_input_fifo_fifo_N16,
      RSTA => rx_input_fifo_fifo_B7_LOGIC_ZERO,
      RSTB => rx_input_fifo_fifo_B7_LOGIC_ZERO,
      WEA => rx_input_fifo_fifo_N17,
      WEB => rx_input_fifo_fifo_B7_LOGIC_ZERO,
      GSR => GSR,
      ADDRA(7) => GLOBAL_LOGIC0_1,
      ADDRA(6) => rx_input_fifo_fifo_N2,
      ADDRA(5) => rx_input_fifo_fifo_N3,
      ADDRA(4) => rx_input_fifo_fifo_N4,
      ADDRA(3) => rx_input_fifo_fifo_N5,
      ADDRA(2) => rx_input_fifo_fifo_N6,
      ADDRA(1) => rx_input_fifo_fifo_N7,
      ADDRA(0) => rx_input_fifo_fifo_N8,
      ADDRB(7) => GLOBAL_LOGIC0_1,
      ADDRB(6) => rx_input_fifo_fifo_N9,
      ADDRB(5) => rx_input_fifo_fifo_N10,
      ADDRB(4) => rx_input_fifo_fifo_N11,
      ADDRB(3) => rx_input_fifo_fifo_N12,
      ADDRB(2) => rx_input_fifo_fifo_N13,
      ADDRB(1) => rx_input_fifo_fifo_N14,
      ADDRB(0) => rx_input_fifo_fifo_N15,
      DIA(15) => GLOBAL_LOGIC0_1,
      DIA(14) => GLOBAL_LOGIC0_1,
      DIA(13) => GLOBAL_LOGIC0_1,
      DIA(12) => GLOBAL_LOGIC0_1,
      DIA(11) => GLOBAL_LOGIC0_1,
      DIA(10) => GLOBAL_LOGIC0_1,
      DIA(9) => GLOBAL_LOGIC0_1,
      DIA(8) => rx_input_endfin,
      DIA(7) => rx_input_fifoin(7),
      DIA(6) => rx_input_fifoin(6),
      DIA(5) => rx_input_fifoin(5),
      DIA(4) => rx_input_fifoin(4),
      DIA(3) => rx_input_fifoin(3),
      DIA(2) => rx_input_fifoin(2),
      DIA(1) => rx_input_fifoin(1),
      DIA(0) => rx_input_fifoin(0),
      DIB(15) => GLOBAL_LOGIC0_1,
      DIB(14) => GLOBAL_LOGIC0_1,
      DIB(13) => GLOBAL_LOGIC0_1,
      DIB(12) => GLOBAL_LOGIC0_1,
      DIB(11) => GLOBAL_LOGIC0_1,
      DIB(10) => GLOBAL_LOGIC0_1,
      DIB(9) => GLOBAL_LOGIC0_1,
      DIB(8) => GLOBAL_LOGIC0_1,
      DIB(7) => GLOBAL_LOGIC0_1,
      DIB(6) => GLOBAL_LOGIC0_1,
      DIB(5) => GLOBAL_LOGIC0_1,
      DIB(4) => GLOBAL_LOGIC0_1,
      DIB(3) => GLOBAL_LOGIC0_1,
      DIB(2) => GLOBAL_LOGIC0_1,
      DIB(1) => GLOBAL_LOGIC0_1,
      DIB(0) => GLOBAL_LOGIC0_1,
      DOA(15) => rx_input_fifo_fifo_B7_DOA15,
      DOA(14) => rx_input_fifo_fifo_B7_DOA14,
      DOA(13) => rx_input_fifo_fifo_B7_DOA13,
      DOA(12) => rx_input_fifo_fifo_B7_DOA12,
      DOA(11) => rx_input_fifo_fifo_B7_DOA11,
      DOA(10) => rx_input_fifo_fifo_B7_DOA10,
      DOA(9) => rx_input_fifo_fifo_B7_DOA9,
      DOA(8) => rx_input_fifo_fifo_B7_DOA8,
      DOA(7) => rx_input_fifo_fifo_B7_DOA7,
      DOA(6) => rx_input_fifo_fifo_B7_DOA6,
      DOA(5) => rx_input_fifo_fifo_B7_DOA5,
      DOA(4) => rx_input_fifo_fifo_B7_DOA4,
      DOA(3) => rx_input_fifo_fifo_B7_DOA3,
      DOA(2) => rx_input_fifo_fifo_B7_DOA2,
      DOA(1) => rx_input_fifo_fifo_B7_DOA1,
      DOA(0) => rx_input_fifo_fifo_B7_DOA0,
      DOB(15) => rx_input_fifo_fifo_B7_DOB15,
      DOB(14) => rx_input_fifo_fifo_B7_DOB14,
      DOB(13) => rx_input_fifo_fifo_B7_DOB13,
      DOB(12) => rx_input_fifo_fifo_B7_DOB12,
      DOB(11) => rx_input_fifo_fifo_B7_DOB11,
      DOB(10) => rx_input_fifo_fifo_B7_DOB10,
      DOB(9) => rx_input_fifo_fifo_B7_DOB9,
      DOB(8) => rx_input_fifo_fifodout(8),
      DOB(7) => rx_input_fifo_fifodout(7),
      DOB(6) => rx_input_fifo_fifodout(6),
      DOB(5) => rx_input_fifo_fifodout(5),
      DOB(4) => rx_input_fifo_fifodout(4),
      DOB(3) => rx_input_fifo_fifodout(3),
      DOB(2) => rx_input_fifo_fifodout(2),
      DOB(1) => rx_input_fifo_fifodout(1),
      DOB(0) => rx_input_fifo_fifodout(0)
    );
  rx_output_fifo_B7_LOGIC_ONE_229 : X_ONE
    port map (
      O => rx_output_fifo_B7_LOGIC_ONE
    );
  rx_output_fifo_B7_LOGIC_ZERO_230 : X_ZERO
    port map (
      O => rx_output_fifo_B7_LOGIC_ZERO
    );
  rx_output_fifo_B7 : X_RAMB4_S16_S16
    generic map(
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      SETUP_ALL => 3025 ps,
      XON => FALSE
    )
    port map (
      CLKA => GTX_CLK_OBUF,
      CLKB => clkio,
      ENA => rx_output_fifo_B7_LOGIC_ONE,
      ENB => rx_output_fifo_N18,
      RSTA => rx_output_fifo_B7_LOGIC_ZERO,
      RSTB => rx_output_fifo_B7_LOGIC_ZERO,
      WEA => rx_output_fifo_N19,
      WEB => rx_output_fifo_B7_LOGIC_ZERO,
      GSR => GSR,
      ADDRA(7) => rx_output_fifo_N2,
      ADDRA(6) => rx_output_fifo_N3,
      ADDRA(5) => rx_output_fifo_N4,
      ADDRA(4) => rx_output_fifo_N5,
      ADDRA(3) => rx_output_fifo_N6,
      ADDRA(2) => rx_output_fifo_N7,
      ADDRA(1) => rx_output_fifo_N8,
      ADDRA(0) => rx_output_fifo_N9,
      ADDRB(7) => rx_output_fifo_N10,
      ADDRB(6) => rx_output_fifo_N11,
      ADDRB(5) => rx_output_fifo_N12,
      ADDRB(4) => rx_output_fifo_N13,
      ADDRB(3) => rx_output_fifo_N14,
      ADDRB(2) => rx_output_fifo_N15,
      ADDRB(1) => rx_output_fifo_N16,
      ADDRB(0) => rx_output_fifo_N17,
      DIA(15) => rx_output_fifodin(15),
      DIA(14) => rx_output_fifodin(14),
      DIA(13) => rx_output_fifodin(13),
      DIA(12) => rx_output_fifodin(12),
      DIA(11) => rx_output_fifodin(11),
      DIA(10) => rx_output_fifodin(10),
      DIA(9) => rx_output_fifodin(9),
      DIA(8) => rx_output_fifodin(8),
      DIA(7) => rx_output_fifodin(7),
      DIA(6) => rx_output_fifodin(6),
      DIA(5) => rx_output_fifodin(5),
      DIA(4) => rx_output_fifodin(4),
      DIA(3) => rx_output_fifodin(3),
      DIA(2) => rx_output_fifodin(2),
      DIA(1) => rx_output_fifodin(1),
      DIA(0) => rx_output_fifodin(0),
      DIB(15) => GLOBAL_LOGIC0_46,
      DIB(14) => GLOBAL_LOGIC0_46,
      DIB(13) => GLOBAL_LOGIC0_46,
      DIB(12) => GLOBAL_LOGIC0_46,
      DIB(11) => GLOBAL_LOGIC0_47,
      DIB(10) => GLOBAL_LOGIC0_46,
      DIB(9) => GLOBAL_LOGIC0_47,
      DIB(8) => GLOBAL_LOGIC0_46,
      DIB(7) => GLOBAL_LOGIC0_46,
      DIB(6) => GLOBAL_LOGIC0_46,
      DIB(5) => GLOBAL_LOGIC0_46,
      DIB(4) => GLOBAL_LOGIC0_46,
      DIB(3) => GLOBAL_LOGIC0_48,
      DIB(2) => GLOBAL_LOGIC0_46,
      DIB(1) => GLOBAL_LOGIC0_47,
      DIB(0) => GLOBAL_LOGIC0_46,
      DOA(15) => rx_output_fifo_B7_DOA15,
      DOA(14) => rx_output_fifo_B7_DOA14,
      DOA(13) => rx_output_fifo_B7_DOA13,
      DOA(12) => rx_output_fifo_B7_DOA12,
      DOA(11) => rx_output_fifo_B7_DOA11,
      DOA(10) => rx_output_fifo_B7_DOA10,
      DOA(9) => rx_output_fifo_B7_DOA9,
      DOA(8) => rx_output_fifo_B7_DOA8,
      DOA(7) => rx_output_fifo_B7_DOA7,
      DOA(6) => rx_output_fifo_B7_DOA6,
      DOA(5) => rx_output_fifo_B7_DOA5,
      DOA(4) => rx_output_fifo_B7_DOA4,
      DOA(3) => rx_output_fifo_B7_DOA3,
      DOA(2) => rx_output_fifo_B7_DOA2,
      DOA(1) => rx_output_fifo_B7_DOA1,
      DOA(0) => rx_output_fifo_B7_DOA0,
      DOB(15) => rx_output_fifodout(15),
      DOB(14) => rx_output_fifodout(14),
      DOB(13) => rx_output_fifodout(13),
      DOB(12) => rx_output_fifodout(12),
      DOB(11) => rx_output_fifodout(11),
      DOB(10) => rx_output_fifodout(10),
      DOB(9) => rx_output_fifodout(9),
      DOB(8) => rx_output_fifodout(8),
      DOB(7) => rx_output_fifodout(7),
      DOB(6) => rx_output_fifodout(6),
      DOB(5) => rx_output_fifodout(5),
      DOB(4) => rx_output_fifodout(4),
      DOB(3) => rx_output_fifodout(3),
      DOB(2) => rx_output_fifodout(2),
      DOB(1) => rx_output_fifodout(1),
      DOB(0) => rx_output_fifodout(0)
    );
  mac_control_Mmux_n0016_Result_20_80 : X_MUX2
    port map (
      IA => mac_control_dout_19_rt,
      IB => mac_control_N81880,
      SEL => mac_control_n0044,
      O => mac_control_n0016(20)
    );
  mac_control_Mmux_n0016_Result_20_80_G : X_LUT4
    generic map(
      INIT => X"00EA"
    )
    port map (
      ADR0 => mac_control_CHOICE2142,
      ADR1 => mac_control_phystat(20),
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_addr(5),
      O => mac_control_N81880
    );
  mac_control_dout_19_rt_231 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_dout(19),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_dout_19_rt
    );
  mac_control_Mmux_n0016_Result_21_84 : X_MUX2
    port map (
      IA => mac_control_dout_20_rt,
      IB => mac_control_N81872,
      SEL => mac_control_n0044,
      O => mac_control_n0016(21)
    );
  mac_control_Mmux_n0016_Result_21_84_G : X_LUT4
    generic map(
      INIT => X"3222"
    )
    port map (
      ADR0 => mac_control_CHOICE2375,
      ADR1 => mac_control_addr(5),
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_phystat(21),
      O => mac_control_N81872
    );
  mac_control_dout_20_rt_232 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_dout(20),
      ADR3 => VCC,
      O => mac_control_dout_20_rt
    );
  mac_control_Mmux_n0016_Result_22_80 : X_MUX2
    port map (
      IA => mac_control_dout_21_rt,
      IB => mac_control_N81896,
      SEL => mac_control_n0044,
      O => mac_control_n0016(22)
    );
  mac_control_Mmux_n0016_Result_22_80_G : X_LUT4
    generic map(
      INIT => X"5450"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_phystat(22),
      ADR2 => mac_control_CHOICE2119,
      ADR3 => mac_control_n0057,
      O => mac_control_N81896
    );
  mac_control_dout_21_rt_233 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_dout(21),
      O => mac_control_dout_21_rt
    );
  mac_control_Mmux_n0016_Result_30_80 : X_MUX2
    port map (
      IA => mac_control_dout_29_rt,
      IB => mac_control_N81884,
      SEL => mac_control_n0044,
      O => mac_control_n0016(30)
    );
  mac_control_Mmux_n0016_Result_30_80_G : X_LUT4
    generic map(
      INIT => X"5450"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_n0057,
      ADR2 => mac_control_CHOICE2303,
      ADR3 => mac_control_phystat(30),
      O => mac_control_N81884
    );
  mac_control_dout_29_rt_234 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_dout(29),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_dout_29_rt
    );
  mac_control_Mmux_n0016_Result_23_80 : X_MUX2
    port map (
      IA => mac_control_dout_22_rt,
      IB => mac_control_N81856,
      SEL => mac_control_n0044,
      O => mac_control_n0016(23)
    );
  mac_control_Mmux_n0016_Result_23_80_G : X_LUT4
    generic map(
      INIT => X"5540"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_phystat(23),
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_CHOICE2165,
      O => mac_control_N81856
    );
  mac_control_dout_22_rt_235 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_dout(22),
      O => mac_control_dout_22_rt
    );
  mac_control_Mmux_n0016_Result_16_84 : X_MUX2
    port map (
      IA => mac_control_dout_15_rt,
      IB => mac_control_N81900,
      SEL => mac_control_n0044,
      O => mac_control_n0016(16)
    );
  mac_control_Mmux_n0016_Result_16_84_G : X_LUT4
    generic map(
      INIT => X"00F8"
    )
    port map (
      ADR0 => mac_control_phystat(16),
      ADR1 => mac_control_n0057,
      ADR2 => mac_control_CHOICE2327,
      ADR3 => mac_control_addr(5),
      O => mac_control_N81900
    );
  mac_control_dout_15_rt_236 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_dout(15),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_dout_15_rt
    );
  rx_input_fifo_fifo_BU136 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifo_N1585,
      CE => rx_input_fifo_fifo_N1497,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_fifo_fifo_N1599_FFX_RST,
      O => rx_input_fifo_fifo_N1599
    );
  rx_input_fifo_fifo_N1599_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_RESET_1,
      I1 => GSR,
      O => rx_input_fifo_fifo_N1599_FFX_RST
    );
  mac_control_Mmux_n0016_Result_24_84 : X_MUX2
    port map (
      IA => mac_control_dout_23_rt,
      IB => mac_control_N81852,
      SEL => mac_control_n0044,
      O => mac_control_n0016(24)
    );
  mac_control_Mmux_n0016_Result_24_84_G : X_LUT4
    generic map(
      INIT => X"0E0A"
    )
    port map (
      ADR0 => mac_control_CHOICE2399,
      ADR1 => mac_control_phystat(24),
      ADR2 => mac_control_addr(5),
      ADR3 => mac_control_n0057,
      O => mac_control_N81852
    );
  mac_control_dout_23_rt_237 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_dout(23),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_dout_23_rt
    );
  mac_control_Mmux_n0016_Result_25_80 : X_MUX2
    port map (
      IA => mac_control_dout_24_rt,
      IB => mac_control_N81876,
      SEL => mac_control_n0044,
      O => mac_control_n0016(25)
    );
  mac_control_Mmux_n0016_Result_25_80_G : X_LUT4
    generic map(
      INIT => X"0E0C"
    )
    port map (
      ADR0 => mac_control_phystat(25),
      ADR1 => mac_control_CHOICE2211,
      ADR2 => mac_control_addr(5),
      ADR3 => mac_control_n0057,
      O => mac_control_N81876
    );
  mac_control_dout_24_rt_238 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_dout(24),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_dout_24_rt
    );
  mac_control_Mmux_n0016_Result_17_84 : X_MUX2
    port map (
      IA => mac_control_dout_16_rt,
      IB => mac_control_N81904,
      SEL => mac_control_n0044,
      O => mac_control_n0016(17)
    );
  mac_control_Mmux_n0016_Result_17_84_G : X_LUT4
    generic map(
      INIT => X"00F8"
    )
    port map (
      ADR0 => mac_control_n0057,
      ADR1 => mac_control_phystat(17),
      ADR2 => mac_control_CHOICE2351,
      ADR3 => mac_control_addr(5),
      O => mac_control_N81904
    );
  mac_control_dout_16_rt_239 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_dout(16),
      ADR3 => VCC,
      O => mac_control_dout_16_rt
    );
  mac_control_Mmux_n0016_Result_26_80 : X_MUX2
    port map (
      IA => mac_control_dout_25_rt,
      IB => mac_control_N81908,
      SEL => mac_control_n0044,
      O => mac_control_n0016(26)
    );
  mac_control_Mmux_n0016_Result_26_80_G : X_LUT4
    generic map(
      INIT => X"5450"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_n0057,
      ADR2 => mac_control_CHOICE2188,
      ADR3 => mac_control_phystat(26),
      O => mac_control_N81908
    );
  mac_control_dout_25_rt_240 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_dout(25),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_dout_25_rt
    );
  mac_control_Mmux_n0016_Result_18_80 : X_MUX2
    port map (
      IA => mac_control_dout_17_rt,
      IB => mac_control_N81868,
      SEL => mac_control_n0044,
      O => mac_control_n0016(18)
    );
  mac_control_Mmux_n0016_Result_18_80_G : X_LUT4
    generic map(
      INIT => X"3222"
    )
    port map (
      ADR0 => mac_control_CHOICE2073,
      ADR1 => mac_control_addr(5),
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_phystat(18),
      O => mac_control_N81868
    );
  mac_control_dout_17_rt_241 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_dout(17),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_dout_17_rt
    );
  mac_control_Mmux_n0016_Result_19_80 : X_MUX2
    port map (
      IA => mac_control_dout_18_rt,
      IB => mac_control_N81892,
      SEL => mac_control_n0044,
      O => mac_control_n0016(19)
    );
  mac_control_Mmux_n0016_Result_19_80_G : X_LUT4
    generic map(
      INIT => X"0E0C"
    )
    port map (
      ADR0 => mac_control_n0057,
      ADR1 => mac_control_CHOICE2096,
      ADR2 => mac_control_addr(5),
      ADR3 => mac_control_phystat(19),
      O => mac_control_N81892
    );
  mac_control_dout_18_rt_242 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_dout(18),
      ADR3 => VCC,
      O => mac_control_dout_18_rt
    );
  mac_control_Mmux_n0016_Result_27_80 : X_MUX2
    port map (
      IA => mac_control_dout_26_rt,
      IB => mac_control_N81860,
      SEL => mac_control_n0044,
      O => mac_control_n0016(27)
    );
  mac_control_Mmux_n0016_Result_27_80_G : X_LUT4
    generic map(
      INIT => X"00EC"
    )
    port map (
      ADR0 => mac_control_n0057,
      ADR1 => mac_control_CHOICE2234,
      ADR2 => mac_control_phystat(27),
      ADR3 => mac_control_addr(5),
      O => mac_control_N81860
    );
  mac_control_dout_26_rt_243 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_dout(26),
      O => mac_control_dout_26_rt
    );
  mac_control_Mmux_n0016_Result_28_80 : X_MUX2
    port map (
      IA => mac_control_dout_27_rt,
      IB => mac_control_N81888,
      SEL => mac_control_n0044,
      O => mac_control_n0016(28)
    );
  mac_control_Mmux_n0016_Result_28_80_G : X_LUT4
    generic map(
      INIT => X"0E0A"
    )
    port map (
      ADR0 => mac_control_CHOICE2257,
      ADR1 => mac_control_phystat(28),
      ADR2 => mac_control_addr(5),
      ADR3 => mac_control_n0057,
      O => mac_control_N81888
    );
  mac_control_dout_27_rt_244 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_dout(27),
      ADR3 => VCC,
      O => mac_control_dout_27_rt
    );
  mac_control_Mmux_n0016_Result_29_80 : X_MUX2
    port map (
      IA => mac_control_dout_28_rt,
      IB => mac_control_N81864,
      SEL => mac_control_n0044,
      O => mac_control_n0016(29)
    );
  mac_control_Mmux_n0016_Result_29_80_G : X_LUT4
    generic map(
      INIT => X"00EC"
    )
    port map (
      ADR0 => mac_control_n0057,
      ADR1 => mac_control_CHOICE2280,
      ADR2 => mac_control_phystat(29),
      ADR3 => mac_control_addr(5),
      O => mac_control_N81864
    );
  mac_control_dout_28_rt_245 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_dout(28),
      O => mac_control_dout_28_rt
    );
  mac_control_phyaddr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_9_FFX_RST,
      O => mac_control_phyaddr(9)
    );
  mac_control_phyaddr_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_9_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_sout414 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_N81846,
      IB => mac_control_PHY_status_MII_Interface_N81848,
      SEL => mac_control_PHY_status_MII_Interface_statecnt(4),
      O => mac_control_PHY_status_MII_Interface_CHOICE977_F5MUX
    );
  mac_control_PHY_status_MII_Interface_sout414_G : X_LUT4
    generic map(
      INIT => X"4540"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_din(9),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR3 => mac_control_PHY_status_din(13),
      O => mac_control_PHY_status_MII_Interface_N81848
    );
  mac_control_PHY_status_MII_Interface_sout414_F : X_LUT4
    generic map(
      INIT => X"0011"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_miirw,
      O => mac_control_PHY_status_MII_Interface_N81846
    );
  mac_control_PHY_status_MII_Interface_CHOICE977_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE977_F5MUX,
      O => mac_control_PHY_status_MII_Interface_CHOICE977
    );
  memcontroller_Mmux_addrn_inst_mux_f5_32111 : X_MUX2
    port map (
      IA => memcontroller_N81726,
      IB => memcontroller_N81728,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_0_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_32111_G : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => addr4ext(0),
      ADR1 => addr2ext(0),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81728
    );
  memcontroller_Mmux_addrn_inst_mux_f5_32111_F : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(0),
      ADR2 => addr1ext(0),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81726
    );
  memcontroller_addrn_0_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_0_F5MUX,
      O => memcontroller_addrn(0)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_40111 : X_MUX2
    port map (
      IA => memcontroller_N81686,
      IB => memcontroller_N81688,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_8_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_40111_G : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr4ext(8),
      ADR2 => addr2ext(8),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81688
    );
  memcontroller_Mmux_addrn_inst_mux_f5_40111_F : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(8),
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => addr1ext(8),
      O => memcontroller_N81686
    );
  memcontroller_addrn_8_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_8_F5MUX,
      O => memcontroller_addrn(8)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_33111 : X_MUX2
    port map (
      IA => memcontroller_N81721,
      IB => memcontroller_N81723,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_1_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_33111_G : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => addr2ext(1),
      ADR1 => VCC,
      ADR2 => addr4ext(1),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81723
    );
  memcontroller_Mmux_addrn_inst_mux_f5_33111_F : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => addr3ext(1),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => addr1ext(1),
      O => memcontroller_N81721
    );
  memcontroller_addrn_1_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_1_F5MUX,
      O => memcontroller_addrn(1)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_41111 : X_MUX2
    port map (
      IA => memcontroller_N81681,
      IB => memcontroller_N81683,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_9_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_41111_G : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(9),
      ADR2 => addr4ext(9),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81683
    );
  memcontroller_Mmux_addrn_inst_mux_f5_41111_F : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr1ext(9),
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => addr3ext(9),
      O => memcontroller_N81681
    );
  memcontroller_addrn_9_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_9_F5MUX,
      O => memcontroller_addrn(9)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_34111 : X_MUX2
    port map (
      IA => memcontroller_N81716,
      IB => memcontroller_N81718,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_2_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_34111_G : X_LUT4
    generic map(
      INIT => X"F3C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_1,
      ADR2 => addr4ext(2),
      ADR3 => addr2ext(2),
      O => memcontroller_N81718
    );
  memcontroller_Mmux_addrn_inst_mux_f5_34111_F : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(2),
      ADR2 => addr1ext(2),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81716
    );
  memcontroller_addrn_2_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_2_F5MUX,
      O => memcontroller_addrn(2)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_42111 : X_MUX2
    port map (
      IA => memcontroller_N81676,
      IB => memcontroller_N81678,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_10_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_42111_G : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => addr4ext(10),
      ADR1 => addr2ext(10),
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => VCC,
      O => memcontroller_N81678
    );
  memcontroller_Mmux_addrn_inst_mux_f5_42111_F : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => addr1ext(10),
      ADR1 => addr3ext(10),
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => VCC,
      O => memcontroller_N81676
    );
  memcontroller_addrn_10_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_10_F5MUX,
      O => memcontroller_addrn(10)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_35111 : X_MUX2
    port map (
      IA => memcontroller_N81711,
      IB => memcontroller_N81713,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_3_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_35111_G : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => addr4ext(3),
      ADR1 => addr2ext(3),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81713
    );
  memcontroller_Mmux_addrn_inst_mux_f5_35111_F : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => addr3ext(3),
      ADR1 => addr1ext(3),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81711
    );
  memcontroller_addrn_3_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_3_F5MUX,
      O => memcontroller_addrn(3)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_43111 : X_MUX2
    port map (
      IA => memcontroller_N81671,
      IB => memcontroller_N81673,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_11_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_43111_G : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => addr2ext(11),
      ADR1 => addr4ext(11),
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => VCC,
      O => memcontroller_N81673
    );
  memcontroller_Mmux_addrn_inst_mux_f5_43111_F : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => addr3ext(11),
      ADR1 => VCC,
      ADR2 => addr1ext(11),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81671
    );
  memcontroller_addrn_11_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_11_F5MUX,
      O => memcontroller_addrn(11)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_36111 : X_MUX2
    port map (
      IA => memcontroller_N81706,
      IB => memcontroller_N81708,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_4_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_36111_G : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(4),
      ADR2 => addr4ext(4),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81708
    );
  memcontroller_Mmux_addrn_inst_mux_f5_36111_F : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => addr1ext(4),
      ADR1 => addr3ext(4),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81706
    );
  memcontroller_addrn_4_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_4_F5MUX,
      O => memcontroller_addrn(4)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_44111 : X_MUX2
    port map (
      IA => memcontroller_N81666,
      IB => memcontroller_N81668,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_12_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_44111_G : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => addr4ext(12),
      ADR1 => memcontroller_clknum_1_1,
      ADR2 => VCC,
      ADR3 => addr2ext(12),
      O => memcontroller_N81668
    );
  memcontroller_Mmux_addrn_inst_mux_f5_44111_F : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(12),
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => addr1ext(12),
      O => memcontroller_N81666
    );
  memcontroller_addrn_12_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_12_F5MUX,
      O => memcontroller_addrn(12)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_37111 : X_MUX2
    port map (
      IA => memcontroller_N81701,
      IB => memcontroller_N81703,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_5_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_37111_G : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => addr2ext(5),
      ADR1 => addr4ext(5),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81703
    );
  memcontroller_Mmux_addrn_inst_mux_f5_37111_F : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => addr3ext(5),
      ADR1 => VCC,
      ADR2 => addr1ext(5),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81701
    );
  memcontroller_addrn_5_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_5_F5MUX,
      O => memcontroller_addrn(5)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_45111 : X_MUX2
    port map (
      IA => memcontroller_N81606,
      IB => memcontroller_N81608,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_13_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_45111_G : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => addr4ext(13),
      ADR1 => addr2ext(13),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81608
    );
  memcontroller_Mmux_addrn_inst_mux_f5_45111_F : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => memcontroller_clknum_1_1,
      ADR1 => addr1ext(13),
      ADR2 => VCC,
      ADR3 => addr3ext(13),
      O => memcontroller_N81606
    );
  memcontroller_addrn_13_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_13_F5MUX,
      O => memcontroller_addrn(13)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_38111 : X_MUX2
    port map (
      IA => memcontroller_N81696,
      IB => memcontroller_N81698,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_6_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_38111_G : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => addr2ext(6),
      ADR1 => addr4ext(6),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81698
    );
  memcontroller_Mmux_addrn_inst_mux_f5_38111_F : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => addr1ext(6),
      ADR1 => addr3ext(6),
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => VCC,
      O => memcontroller_N81696
    );
  memcontroller_addrn_6_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_6_F5MUX,
      O => memcontroller_addrn(6)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_46111 : X_MUX2
    port map (
      IA => memcontroller_N81601,
      IB => memcontroller_N81603,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_14_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_46111_G : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(14),
      ADR2 => memcontroller_clknum_1_1,
      ADR3 => addr4ext(14),
      O => memcontroller_N81603
    );
  memcontroller_Mmux_addrn_inst_mux_f5_46111_F : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => addr1ext(14),
      ADR1 => VCC,
      ADR2 => addr3ext(14),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81601
    );
  memcontroller_addrn_14_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_14_F5MUX,
      O => memcontroller_addrn(14)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_39111 : X_MUX2
    port map (
      IA => memcontroller_N81691,
      IB => memcontroller_N81693,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_7_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_39111_G : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr4ext(7),
      ADR2 => addr2ext(7),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81693
    );
  memcontroller_Mmux_addrn_inst_mux_f5_39111_F : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => addr3ext(7),
      ADR1 => VCC,
      ADR2 => addr1ext(7),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81691
    );
  memcontroller_addrn_7_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_7_F5MUX,
      O => memcontroller_addrn(7)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_47111 : X_MUX2
    port map (
      IA => memcontroller_N81611,
      IB => memcontroller_N81613,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_15_F5MUX
    );
  memcontroller_Mmux_addrn_inst_mux_f5_47111_G : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(15),
      ADR2 => addr4ext(15),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81613
    );
  memcontroller_Mmux_addrn_inst_mux_f5_47111_F : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(15),
      ADR2 => addr1ext(15),
      ADR3 => memcontroller_clknum_1_1,
      O => memcontroller_N81611
    );
  memcontroller_addrn_15_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_15_F5MUX,
      O => memcontroller_addrn(15)
    );
  memcontroller_Mmux_addrn_inst_mux_f5_48111 : X_MUX2
    port map (
      IA => memcontroller_addrn_16_GROM,
      IB => memcontroller_addrn_16_FROM,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_addrn_16_F5MUX
    );
  memcontroller_addrn_16_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_addrn_16_FROM
    );
  memcontroller_addrn_16_G : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_addrn_16_GROM
    );
  memcontroller_addrn_16_XUSED : X_BUF
    port map (
      I => memcontroller_addrn_16_F5MUX,
      O => memcontroller_addrn(16)
    );
  memcontroller_Mmux_dn_inst_mux_f5_10111 : X_MUX2
    port map (
      IA => memcontroller_N81826,
      IB => memcontroller_N81828,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(10)
    );
  memcontroller_Mmux_dn_inst_mux_f5_10111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => d4(10),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_3,
      ADR3 => VCC,
      O => memcontroller_N81828
    );
  memcontroller_Mmux_dn_inst_mux_f5_10111_F : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => memcontroller_clknum_1_3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(10),
      O => memcontroller_N81826
    );
  memcontroller_dnl1_10_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_10_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_11011 : X_MUX2
    port map (
      IA => memcontroller_N81781,
      IB => memcontroller_N81783,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(1)
    );
  memcontroller_Mmux_dn_inst_mux_f5_11011_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_3,
      O => memcontroller_N81783
    );
  memcontroller_Mmux_dn_inst_mux_f5_11011_F : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(1),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_3,
      O => memcontroller_N81781
    );
  memcontroller_dnl1_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_1_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_11111 : X_MUX2
    port map (
      IA => memcontroller_N81831,
      IB => memcontroller_N81833,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(11)
    );
  memcontroller_Mmux_dn_inst_mux_f5_11111_G : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(11),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_3,
      O => memcontroller_N81833
    );
  memcontroller_Mmux_dn_inst_mux_f5_11111_F : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_3,
      ADR2 => d1(11),
      ADR3 => VCC,
      O => memcontroller_N81831
    );
  memcontroller_dnl1_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_11_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_0111 : X_MUX2
    port map (
      IA => memcontroller_N81776,
      IB => memcontroller_N81778,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(0)
    );
  memcontroller_Mmux_dn_inst_mux_f5_0111_G : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => d4(0),
      ADR1 => memcontroller_clknum_1_3,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N81778
    );
  memcontroller_Mmux_dn_inst_mux_f5_0111_F : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_3,
      ADR2 => VCC,
      ADR3 => d1(0),
      O => memcontroller_N81776
    );
  memcontroller_dnl1_0_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_0_CEMUXNOT
    );
  rx_input_memio_addrchk_n0052_SW0 : X_LUT4
    generic map(
      INIT => X"8800"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_maceq(5),
      ADR1 => rx_input_memio_addrchk_maceq(4),
      ADR2 => VCC,
      ADR3 => rx_input_memio_addrchk_maceq(3),
      O => rx_input_memio_addrchk_validucast_FROM
    );
  rx_input_memio_addrchk_n0052_246 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_maceq(0),
      ADR1 => rx_input_memio_addrchk_maceq(1),
      ADR2 => rx_input_memio_addrchk_maceq(2),
      ADR3 => rx_input_memio_addrchk_N70335,
      O => rx_input_memio_addrchk_n0052
    );
  rx_input_memio_addrchk_validucast_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_validucast_CEMUXNOT
    );
  rx_input_memio_addrchk_validucast_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_validucast_FROM,
      O => rx_input_memio_addrchk_N70335
    );
  mac_control_rxfifowerr_cntl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(19),
      CE => mac_control_rxfifowerr_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_19_FFX_RST,
      O => mac_control_rxfifowerr_cntl(19)
    );
  mac_control_rxfifowerr_cntl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_19_FFX_RST
    );
  rx_input_memio_bpen_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_bpen_CEMUXNOT
    );
  rx_input_memio_addrchk_n0053_SW0 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_rxbcastl,
      ADR1 => rx_input_memio_addrchk_validmcast,
      ADR2 => rx_input_memio_addrchk_validbcast,
      ADR3 => rx_input_memio_addrchk_rxmcastl,
      O => rx_input_memio_destok_FROM
    );
  rx_input_memio_addrchk_n0053_247 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_rxallfl,
      ADR1 => rx_input_memio_addrchk_rxucastl,
      ADR2 => rx_input_memio_addrchk_validucast,
      ADR3 => rx_input_memio_addrchk_N72932,
      O => rx_input_memio_addrchk_n0053
    );
  rx_input_memio_destok_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_destok_CEMUXNOT
    );
  rx_input_memio_destok_XUSED : X_BUF
    port map (
      I => rx_input_memio_destok_FROM,
      O => rx_input_memio_addrchk_N72932
    );
  rx_output_cs_FFd10_In4 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_output_cs_FFd3,
      ADR1 => rx_output_cs_FFd4,
      ADR2 => rx_output_cs_FFd2,
      ADR3 => rx_output_cs_FFd5,
      O => rx_output_cs_FFd10_FROM
    );
  rx_output_cs_FFd10_In26 : X_LUT4
    generic map(
      INIT => X"3332"
    )
    port map (
      ADR0 => rx_output_CHOICE1800,
      ADR1 => rx_output_nf,
      ADR2 => rx_output_N34486,
      ADR3 => rx_output_CHOICE1797,
      O => rx_output_cs_FFd10_In
    );
  rx_output_cs_FFd10_XUSED : X_BUF
    port map (
      I => rx_output_cs_FFd10_FROM,
      O => rx_output_CHOICE1797
    );
  tx_output_crc_loigc_Mxor_CO_26_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(3),
      ADR1 => tx_output_crcl(24),
      ADR2 => tx_output_crcl(28),
      ADR3 => tx_output_data(7),
      O => tx_output_crc_loigc_Mxor_CO_26_Xo_1_GROM
    );
  tx_output_crc_loigc_Mxor_CO_26_Xo_1_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_26_Xo_1_GROM,
      O => tx_output_crc_loigc_Mxor_CO_26_Xo(1)
    );
  tx_output_crc_loigc_Mxor_CO_18_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(0),
      ADR1 => tx_output_crc_loigc_Mxor_CO_18_Xo(0),
      ADR2 => tx_output_crcl(10),
      ADR3 => tx_output_crcl(31),
      O => tx_output_crcl_18_FROM
    );
  tx_output_n0034_18_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16_1,
      ADR2 => VCC,
      ADR3 => tx_output_crc_18_Q,
      O => tx_output_n0034_18_Q
    );
  tx_output_crcl_18_XUSED : X_BUF
    port map (
      I => tx_output_crcl_18_FROM,
      O => tx_output_crc_18_Q
    );
  tx_output_crc_loigc_Mxor_CO_26_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0124(1),
      ADR1 => tx_output_crcl(18),
      ADR2 => tx_output_crc_loigc_n0104(0),
      ADR3 => tx_output_crc_loigc_Mxor_CO_26_Xo(1),
      O => tx_output_crcl_26_FROM
    );
  tx_output_n0034_26_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_26_Q,
      O => tx_output_n0034_26_Q
    );
  tx_output_crcl_26_XUSED : X_BUF
    port map (
      I => tx_output_crcl_26_FROM,
      O => tx_output_crc_26_Q
    );
  mac_control_rxfifowerr_cntl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(29),
      CE => mac_control_rxfifowerr_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_29_FFX_RST,
      O => mac_control_rxfifowerr_cntl(29)
    );
  mac_control_rxfifowerr_cntl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_29_FFX_RST
    );
  rx_input_memio_crccomb_Mxor_CO_13_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_datal(0),
      ADR1 => rx_input_memio_datal(4),
      ADR2 => rx_input_memio_crcl(27),
      ADR3 => rx_input_memio_crcl(31),
      O => rx_input_memio_crcl_19_FROM
    );
  rx_input_memio_n0048_19_1 : X_LUT4
    generic map(
      INIT => X"F5FA"
    )
    port map (
      ADR0 => rx_input_memio_crcl(11),
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crccomb_Mxor_CO_13_Xo(2),
      O => rx_input_memio_n0048_19_Q
    );
  rx_input_memio_crcl_19_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_19_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_13_Xo(2)
    );
  rx_input_memio_crccomb_Mxor_CO_13_Xo_5_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(5),
      ADR1 => rx_input_memio_crccomb_Mxor_CO_18_Xo(0),
      ADR2 => rx_input_memio_crccomb_Mxor_n0007_Xo(0),
      ADR3 => rx_input_memio_crccomb_Mxor_CO_13_Xo(2),
      O => rx_input_memio_crcl_13_FROM
    );
  rx_input_memio_n0048_13_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_13_Q,
      O => rx_input_memio_n0048_13_Q
    );
  rx_input_memio_crcl_13_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_13_FROM,
      O => rx_input_memio_crc_13_Q
    );
  tx_output_crc_loigc_Mxor_CO_27_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0118(0),
      ADR1 => tx_output_crc_loigc_Mxor_CO_9_Xo(0),
      ADR2 => tx_output_crc_loigc_n0124(0),
      ADR3 => tx_output_crcl(19),
      O => tx_output_crcl_27_FROM
    );
  tx_output_n0034_27_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16_1,
      ADR3 => tx_output_crc_27_Q,
      O => tx_output_n0034_27_Q
    );
  tx_output_crcl_27_XUSED : X_BUF
    port map (
      I => tx_output_crcl_27_FROM,
      O => tx_output_crc_27_Q
    );
  rx_output_cs_FFd6_In10 : X_LUT4
    generic map(
      INIT => X"FF8C"
    )
    port map (
      ADR0 => rx_output_fifo_nearfull,
      ADR1 => rx_output_cs_FFd6,
      ADR2 => clken3,
      ADR3 => rx_output_CHOICE1106,
      O => rx_output_cs_FFd6_FROM
    );
  rx_output_cs_FFd6_In12 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rx_output_nf,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_CHOICE1110,
      O => rx_output_cs_FFd6_In
    );
  rx_output_cs_FFd6_XUSED : X_BUF
    port map (
      I => rx_output_cs_FFd6_FROM,
      O => rx_output_CHOICE1110
    );
  rx_input_memio_crccomb_Mxor_CO_30_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(22),
      ADR1 => rx_input_memio_datal(0),
      ADR2 => rx_input_memio_crccomb_n0115(0),
      ADR3 => rx_input_memio_crcl(31),
      O => rx_input_memio_crcl_30_FROM
    );
  rx_input_memio_n0048_30_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_30_Q,
      O => rx_input_memio_n0048_30_1_O
    );
  rx_input_memio_crcl_30_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_30_FROM,
      O => rx_input_memio_crc_30_Q
    );
  rx_input_memio_crccomb_Mxor_CO_14_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(26),
      ADR1 => rx_input_memio_crccomb_N81261,
      ADR2 => rx_input_memio_crccomb_n0104(0),
      ADR3 => rx_input_memio_crccomb_Mxor_CO_13_Xo(2),
      O => rx_input_memio_crcl_14_FROM
    );
  rx_input_memio_n0048_14_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_14_Q,
      O => rx_input_memio_n0048_14_Q
    );
  rx_input_memio_crcl_14_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_14_FROM,
      O => rx_input_memio_crc_14_Q
    );
  tx_input_cs_FFd12_In_SW0 : X_LUT4
    generic map(
      INIT => X"FAFA"
    )
    port map (
      ADR0 => txfifowerr,
      ADR1 => VCC,
      ADR2 => tx_input_DONE,
      ADR3 => VCC,
      O => tx_input_cs_FFd12_FROM
    );
  tx_input_cs_FFd12_In_248 : X_LUT4
    generic map(
      INIT => X"FF4C"
    )
    port map (
      ADR0 => tx_input_den,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => tx_input_newfint,
      ADR3 => tx_input_N70123,
      O => tx_input_cs_FFd12_In
    );
  tx_input_cs_FFd12_XUSED : X_BUF
    port map (
      I => tx_input_cs_FFd12_FROM,
      O => tx_input_N70123
    );
  mac_control_rxcrcerr_cntl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_1_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_3_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_5_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_7_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_9_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_11_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_11_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_21_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(20),
      CE => rx_input_memio_addrchk_macaddrl_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_21_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(20)
    );
  rx_input_memio_addrchk_macaddrl_21_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_21_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_13_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(12),
      CE => rx_input_memio_addrchk_macaddrl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_13_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(12)
    );
  rx_input_memio_addrchk_macaddrl_13_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_13_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_31_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(30),
      CE => rx_input_memio_addrchk_macaddrl_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_31_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(30)
    );
  rx_input_memio_addrchk_macaddrl_31_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_31_CEMUXNOT
    );
  tx_input_fifofulll_249 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfifofull,
      CE => tx_input_fifofulll_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_fifofulll_FFY_RST,
      O => tx_input_fifofulll
    );
  tx_input_fifofulll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_fifofulll_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_23_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(22),
      CE => rx_input_memio_addrchk_macaddrl_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_23_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(22)
    );
  rx_input_memio_addrchk_macaddrl_23_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_23_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_15_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(14),
      CE => rx_input_memio_addrchk_macaddrl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_15_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(14)
    );
  rx_input_memio_addrchk_macaddrl_15_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_15_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_41_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_41_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_33_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_32 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(32),
      CE => rx_input_memio_addrchk_macaddrl_33_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_33_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(32)
    );
  rx_input_memio_addrchk_macaddrl_33_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_33_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_25_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(24),
      CE => rx_input_memio_addrchk_macaddrl_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_25_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(24)
    );
  rx_input_memio_addrchk_macaddrl_25_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_25_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_17_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(16),
      CE => rx_input_memio_addrchk_macaddrl_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_17_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(16)
    );
  rx_input_memio_addrchk_macaddrl_17_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_17_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_43_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_42 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(42),
      CE => rx_input_memio_addrchk_macaddrl_43_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_43_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(42)
    );
  rx_input_memio_addrchk_macaddrl_43_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_43_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_12111 : X_MUX2
    port map (
      IA => memcontroller_N81836,
      IB => memcontroller_N81838,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(12)
    );
  memcontroller_Mmux_dn_inst_mux_f5_12111_G : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_3,
      ADR2 => d4(12),
      ADR3 => VCC,
      O => memcontroller_N81838
    );
  memcontroller_Mmux_dn_inst_mux_f5_12111_F : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_3,
      ADR3 => d1(12),
      O => memcontroller_N81836
    );
  memcontroller_dnl1_12_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_12_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_20111 : X_MUX2
    port map (
      IA => memcontroller_N81651,
      IB => memcontroller_N81653,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(20)
    );
  memcontroller_Mmux_dn_inst_mux_f5_20111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(20),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_3,
      O => memcontroller_N81653
    );
  memcontroller_Mmux_dn_inst_mux_f5_20111_F : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => memcontroller_clknum_1_3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(20),
      O => memcontroller_N81651
    );
  memcontroller_dnl1_20_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_20_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_21011 : X_MUX2
    port map (
      IA => memcontroller_N81786,
      IB => memcontroller_N81788,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(2)
    );
  memcontroller_Mmux_dn_inst_mux_f5_21011_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => memcontroller_clknum_1_3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d4(2),
      O => memcontroller_N81788
    );
  memcontroller_Mmux_dn_inst_mux_f5_21011_F : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => memcontroller_clknum_1_3,
      ADR1 => d1(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N81786
    );
  memcontroller_dnl1_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_2_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_21111 : X_MUX2
    port map (
      IA => memcontroller_N81656,
      IB => memcontroller_N81658,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(21)
    );
  memcontroller_Mmux_dn_inst_mux_f5_21111_G : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_3,
      ADR2 => VCC,
      ADR3 => d4(21),
      O => memcontroller_N81658
    );
  memcontroller_Mmux_dn_inst_mux_f5_21111_F : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_3,
      ADR3 => d1(21),
      O => memcontroller_N81656
    );
  memcontroller_dnl1_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_21_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_13111 : X_MUX2
    port map (
      IA => memcontroller_N81841,
      IB => memcontroller_N81843,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(13)
    );
  memcontroller_Mmux_dn_inst_mux_f5_13111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d4(13),
      ADR3 => memcontroller_clknum_1_3,
      O => memcontroller_N81843
    );
  memcontroller_Mmux_dn_inst_mux_f5_13111_F : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_3,
      ADR2 => VCC,
      ADR3 => d1(13),
      O => memcontroller_N81841
    );
  memcontroller_dnl1_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_13_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_30111 : X_MUX2
    port map (
      IA => memcontroller_N81736,
      IB => memcontroller_N81738,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(30)
    );
  memcontroller_Mmux_dn_inst_mux_f5_30111_G : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => d4(30),
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N81738
    );
  memcontroller_Mmux_dn_inst_mux_f5_30111_F : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => d1(30),
      ADR3 => VCC,
      O => memcontroller_N81736
    );
  memcontroller_dnl1_30_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_30_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_22111 : X_MUX2
    port map (
      IA => memcontroller_N81661,
      IB => memcontroller_N81663,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(22)
    );
  memcontroller_Mmux_dn_inst_mux_f5_22111_G : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(22),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_3,
      O => memcontroller_N81663
    );
  memcontroller_Mmux_dn_inst_mux_f5_22111_F : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_3,
      ADR2 => d1(22),
      ADR3 => VCC,
      O => memcontroller_N81661
    );
  memcontroller_dnl1_22_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_22_CEMUXNOT
    );
  rx_input_memio_dout_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_1_FFY_RST,
      O => rx_input_memio_dout(0)
    );
  rx_input_memio_dout_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_1_FFY_RST
    );
  memcontroller_Mmux_dn_inst_mux_f5_14111 : X_MUX2
    port map (
      IA => memcontroller_N81621,
      IB => memcontroller_N81623,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(14)
    );
  memcontroller_Mmux_dn_inst_mux_f5_14111_G : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => memcontroller_clknum_1_3,
      ADR1 => d4(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N81623
    );
  memcontroller_Mmux_dn_inst_mux_f5_14111_F : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => memcontroller_clknum_1_3,
      ADR1 => VCC,
      ADR2 => d1(14),
      ADR3 => VCC,
      O => memcontroller_N81621
    );
  memcontroller_dnl1_14_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_14_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_31111 : X_MUX2
    port map (
      IA => memcontroller_N81771,
      IB => memcontroller_N81773,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(31)
    );
  memcontroller_Mmux_dn_inst_mux_f5_31111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => d4(31),
      ADR3 => VCC,
      O => memcontroller_N81773
    );
  memcontroller_Mmux_dn_inst_mux_f5_31111_F : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => d1(31),
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N81771
    );
  memcontroller_dnl1_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_31_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_15111 : X_MUX2
    port map (
      IA => memcontroller_N81626,
      IB => memcontroller_N81628,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(15)
    );
  memcontroller_Mmux_dn_inst_mux_f5_15111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d4(15),
      ADR3 => memcontroller_clknum_1_3,
      O => memcontroller_N81628
    );
  memcontroller_Mmux_dn_inst_mux_f5_15111_F : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => memcontroller_clknum_1_3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(15),
      O => memcontroller_N81626
    );
  memcontroller_dnl1_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_15_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_23111 : X_MUX2
    port map (
      IA => memcontroller_N81616,
      IB => memcontroller_N81618,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(23)
    );
  memcontroller_Mmux_dn_inst_mux_f5_23111_G : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(23),
      ADR2 => memcontroller_clknum_1_3,
      ADR3 => VCC,
      O => memcontroller_N81618
    );
  memcontroller_Mmux_dn_inst_mux_f5_23111_F : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(23),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N81616
    );
  memcontroller_dnl1_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_23_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_3211 : X_MUX2
    port map (
      IA => memcontroller_N81791,
      IB => memcontroller_N81793,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(3)
    );
  memcontroller_Mmux_dn_inst_mux_f5_3211_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d4(3),
      O => memcontroller_N81793
    );
  memcontroller_Mmux_dn_inst_mux_f5_3211_F : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d1(3),
      O => memcontroller_N81791
    );
  memcontroller_dnl1_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_3_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_4111 : X_MUX2
    port map (
      IA => memcontroller_N81796,
      IB => memcontroller_N81798,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(4)
    );
  memcontroller_Mmux_dn_inst_mux_f5_4111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => d4(4),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N81798
    );
  memcontroller_Mmux_dn_inst_mux_f5_4111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(4),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N81796
    );
  memcontroller_dnl1_4_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_4_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_24111 : X_MUX2
    port map (
      IA => memcontroller_N81766,
      IB => memcontroller_N81768,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(24)
    );
  memcontroller_Mmux_dn_inst_mux_f5_24111_G : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(24),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N81768
    );
  memcontroller_Mmux_dn_inst_mux_f5_24111_F : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d1(24),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N81766
    );
  memcontroller_dnl1_24_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_24_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_16111 : X_MUX2
    port map (
      IA => memcontroller_N81631,
      IB => memcontroller_N81633,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(16)
    );
  memcontroller_Mmux_dn_inst_mux_f5_16111_G : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d4(16),
      ADR2 => memcontroller_clknum_1_3,
      ADR3 => VCC,
      O => memcontroller_N81633
    );
  memcontroller_Mmux_dn_inst_mux_f5_16111_F : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => memcontroller_clknum_1_3,
      ADR1 => VCC,
      ADR2 => d1(16),
      ADR3 => VCC,
      O => memcontroller_N81631
    );
  memcontroller_dnl1_16_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_16_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_5111 : X_MUX2
    port map (
      IA => memcontroller_N81801,
      IB => memcontroller_N81803,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(5)
    );
  memcontroller_Mmux_dn_inst_mux_f5_5111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d4(5),
      O => memcontroller_N81803
    );
  memcontroller_Mmux_dn_inst_mux_f5_5111_F : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(5),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N81801
    );
  memcontroller_dnl1_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_5_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_25111 : X_MUX2
    port map (
      IA => memcontroller_N81761,
      IB => memcontroller_N81763,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(25)
    );
  memcontroller_Mmux_dn_inst_mux_f5_25111_G : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => d4(25),
      ADR3 => VCC,
      O => memcontroller_N81763
    );
  memcontroller_Mmux_dn_inst_mux_f5_25111_F : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d1(25),
      O => memcontroller_N81761
    );
  memcontroller_dnl1_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_25_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_17111 : X_MUX2
    port map (
      IA => memcontroller_N81636,
      IB => memcontroller_N81638,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(17)
    );
  memcontroller_Mmux_dn_inst_mux_f5_17111_G : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => memcontroller_clknum_1_3,
      ADR1 => d4(17),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N81638
    );
  memcontroller_Mmux_dn_inst_mux_f5_17111_F : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => d1(17),
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_3,
      ADR3 => VCC,
      O => memcontroller_N81636
    );
  memcontroller_dnl1_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_17_CEMUXNOT
    );
  tx_output_FBBP_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(10),
      CE => txfbbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_11_FFY_RST,
      O => txfbbp(10)
    );
  txfbbp_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_11_FFY_RST
    );
  memcontroller_Mmux_dn_inst_mux_f5_6111 : X_MUX2
    port map (
      IA => memcontroller_N81806,
      IB => memcontroller_N81808,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(6)
    );
  memcontroller_Mmux_dn_inst_mux_f5_6111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d4(6),
      O => memcontroller_N81808
    );
  memcontroller_Mmux_dn_inst_mux_f5_6111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(6),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N81806
    );
  memcontroller_dnl1_6_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_6_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_26111 : X_MUX2
    port map (
      IA => memcontroller_N81756,
      IB => memcontroller_N81758,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(26)
    );
  memcontroller_Mmux_dn_inst_mux_f5_26111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d4(26),
      O => memcontroller_N81758
    );
  memcontroller_Mmux_dn_inst_mux_f5_26111_F : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => d1(26),
      ADR3 => VCC,
      O => memcontroller_N81756
    );
  memcontroller_dnl1_26_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_26_CEMUXNOT
    );
  rx_input_memio_dout_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_1_FFX_RST,
      O => rx_input_memio_dout(1)
    );
  rx_input_memio_dout_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_1_FFX_RST
    );
  memcontroller_Mmux_dn_inst_mux_f5_18111 : X_MUX2
    port map (
      IA => memcontroller_N81641,
      IB => memcontroller_N81643,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(18)
    );
  memcontroller_Mmux_dn_inst_mux_f5_18111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(18),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_3,
      O => memcontroller_N81643
    );
  memcontroller_Mmux_dn_inst_mux_f5_18111_F : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => memcontroller_clknum_1_3,
      ADR1 => d1(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N81641
    );
  memcontroller_dnl1_18_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_18_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_7111 : X_MUX2
    port map (
      IA => memcontroller_N81811,
      IB => memcontroller_N81813,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(7)
    );
  memcontroller_Mmux_dn_inst_mux_f5_7111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d4(7),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N81813
    );
  memcontroller_Mmux_dn_inst_mux_f5_7111_F : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => d1(7),
      O => memcontroller_N81811
    );
  memcontroller_dnl1_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_7_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_27111 : X_MUX2
    port map (
      IA => memcontroller_N81751,
      IB => memcontroller_N81753,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(27)
    );
  memcontroller_Mmux_dn_inst_mux_f5_27111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => d4(27),
      O => memcontroller_N81753
    );
  memcontroller_Mmux_dn_inst_mux_f5_27111_F : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => memcontroller_clknum_1_2,
      ADR1 => VCC,
      ADR2 => d1(27),
      ADR3 => VCC,
      O => memcontroller_N81751
    );
  memcontroller_dnl1_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_27_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_19111 : X_MUX2
    port map (
      IA => memcontroller_N81646,
      IB => memcontroller_N81648,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(19)
    );
  memcontroller_Mmux_dn_inst_mux_f5_19111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d4(19),
      ADR3 => memcontroller_clknum_1_3,
      O => memcontroller_N81648
    );
  memcontroller_Mmux_dn_inst_mux_f5_19111_F : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_3,
      ADR2 => VCC,
      ADR3 => d1(19),
      O => memcontroller_N81646
    );
  memcontroller_dnl1_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_19_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_8111 : X_MUX2
    port map (
      IA => memcontroller_N81816,
      IB => memcontroller_N81818,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(8)
    );
  memcontroller_Mmux_dn_inst_mux_f5_8111_G : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => d4(8),
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N81818
    );
  memcontroller_Mmux_dn_inst_mux_f5_8111_F : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(8),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N81816
    );
  memcontroller_dnl1_8_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_8_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_28111 : X_MUX2
    port map (
      IA => memcontroller_N81746,
      IB => memcontroller_N81748,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(28)
    );
  memcontroller_Mmux_dn_inst_mux_f5_28111_G : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => d4(28),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N81748
    );
  memcontroller_Mmux_dn_inst_mux_f5_28111_F : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(28),
      ADR2 => VCC,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_N81746
    );
  memcontroller_dnl1_28_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_28_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_9111 : X_MUX2
    port map (
      IA => memcontroller_N81821,
      IB => memcontroller_N81823,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(9)
    );
  memcontroller_Mmux_dn_inst_mux_f5_9111_G : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => VCC,
      ADR3 => d4(9),
      O => memcontroller_N81823
    );
  memcontroller_Mmux_dn_inst_mux_f5_9111_F : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => VCC,
      ADR3 => d1(9),
      O => memcontroller_N81821
    );
  memcontroller_dnl1_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_9_CEMUXNOT
    );
  memcontroller_Mmux_dn_inst_mux_f5_29111 : X_MUX2
    port map (
      IA => memcontroller_N81741,
      IB => memcontroller_N81743,
      SEL => memcontroller_clknum_0_1,
      O => memcontroller_dn(29)
    );
  memcontroller_Mmux_dn_inst_mux_f5_29111_G : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => d4(29),
      ADR1 => memcontroller_clknum_1_2,
      ADR2 => VCC,
      ADR3 => VCC,
      O => memcontroller_N81743
    );
  memcontroller_Mmux_dn_inst_mux_f5_29111_F : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => d1(29),
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_N81741
    );
  memcontroller_dnl1_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl1_29_CEMUXNOT
    );
  mac_control_PHY_status_MII_Interface_n0076_1_LOGIC_ZERO_250 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_n0076_1_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_181_251 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_31,
      IB => mac_control_PHY_status_MII_Interface_n0076_1_LOGIC_ZERO,
      SEL => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_lut2_127,
      O => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_181
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_lut2_1271 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_31,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_lut2_127
    );
  mac_control_PHY_status_MII_Interface_n0076_1_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_45,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(1),
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_n0076_1_GROM
    );
  mac_control_PHY_status_MII_Interface_n0076_1_COUTUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0076_1_CYMUXG,
      O => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_182
    );
  mac_control_PHY_status_MII_Interface_n0076_1_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0076_1_XORG,
      O => mac_control_PHY_status_MII_Interface_n0076(1)
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_182_252 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_45,
      IB => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_181,
      SEL => mac_control_PHY_status_MII_Interface_n0076_1_GROM,
      O => mac_control_PHY_status_MII_Interface_n0076_1_CYMUXG
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_sum_160 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_181,
      I1 => mac_control_PHY_status_MII_Interface_n0076_1_GROM,
      O => mac_control_PHY_status_MII_Interface_n0076_1_XORG
    );
  mac_control_PHY_status_MII_Interface_n0076_2_LOGIC_ZERO_253 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_n0076_2_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_183_254 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_n0076_2_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_n0076_2_CYINIT,
      SEL => mac_control_PHY_status_MII_Interface_n0076_2_FROM,
      O => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_183
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_sum_161 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_n0076_2_CYINIT,
      I1 => mac_control_PHY_status_MII_Interface_n0076_2_FROM,
      O => mac_control_PHY_status_MII_Interface_n0076_2_XORF
    );
  mac_control_PHY_status_MII_Interface_n0076_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(2),
      O => mac_control_PHY_status_MII_Interface_n0076_2_FROM
    );
  mac_control_PHY_status_MII_Interface_n0076_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_n0076_2_GROM
    );
  mac_control_PHY_status_MII_Interface_n0076_2_COUTUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0076_2_CYMUXG,
      O => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_184
    );
  mac_control_PHY_status_MII_Interface_n0076_2_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0076_2_XORF,
      O => mac_control_PHY_status_MII_Interface_n0076(2)
    );
  mac_control_PHY_status_MII_Interface_n0076_2_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0076_2_XORG,
      O => mac_control_PHY_status_MII_Interface_n0076(3)
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_184_255 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_n0076_2_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_183,
      SEL => mac_control_PHY_status_MII_Interface_n0076_2_GROM,
      O => mac_control_PHY_status_MII_Interface_n0076_2_CYMUXG
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_sum_162 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_183,
      I1 => mac_control_PHY_status_MII_Interface_n0076_2_GROM,
      O => mac_control_PHY_status_MII_Interface_n0076_2_XORG
    );
  mac_control_PHY_status_MII_Interface_n0076_2_CYINIT_256 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_182,
      O => mac_control_PHY_status_MII_Interface_n0076_2_CYINIT
    );
  mac_control_PHY_status_MII_Interface_n0076_4_LOGIC_ZERO_257 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_n0076_4_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_185_258 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_n0076_4_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_n0076_4_CYINIT,
      SEL => mac_control_PHY_status_MII_Interface_n0076_4_FROM,
      O => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_185
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_sum_163 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_n0076_4_CYINIT,
      I1 => mac_control_PHY_status_MII_Interface_n0076_4_FROM,
      O => mac_control_PHY_status_MII_Interface_n0076_4_XORF
    );
  mac_control_PHY_status_MII_Interface_n0076_4_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(4),
      O => mac_control_PHY_status_MII_Interface_n0076_4_FROM
    );
  mac_control_PHY_status_MII_Interface_statecnt_5_rt_259 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_statecnt_5_rt
    );
  mac_control_PHY_status_MII_Interface_n0076_4_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0076_4_XORF,
      O => mac_control_PHY_status_MII_Interface_n0076(4)
    );
  mac_control_PHY_status_MII_Interface_n0076_4_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_n0076_4_XORG,
      O => mac_control_PHY_status_MII_Interface_n0076(5)
    );
  mac_control_PHY_status_MII_Interface_Madd_n0076_inst_sum_164 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_185,
      I1 => mac_control_PHY_status_MII_Interface_statecnt_5_rt,
      O => mac_control_PHY_status_MII_Interface_n0076_4_XORG
    );
  mac_control_PHY_status_MII_Interface_n0076_4_CYINIT_260 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_Madd_n0076_inst_cy_184,
      O => mac_control_PHY_status_MII_Interface_n0076_4_CYINIT
    );
  tx_output_FBBP_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(11),
      CE => txfbbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_11_FFX_RST,
      O => txfbbp(11)
    );
  txfbbp_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_11_FFX_RST
    );
  addr2ext_0_LOGIC_ZERO_261 : X_ZERO
    port map (
      O => addr2ext_0_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_0_262 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_8,
      IB => addr2ext_0_LOGIC_ZERO,
      SEL => tx_output_addr_Madd_n0000_inst_lut2_0,
      O => tx_output_addr_Madd_n0000_inst_cy_0
    );
  tx_output_addr_Madd_n0000_inst_lut2_01 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_8,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(0),
      O => tx_output_addr_Madd_n0000_inst_lut2_0
    );
  addr2ext_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_15,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(1),
      O => addr2ext_0_GROM
    );
  addr2ext_0_COUTUSED : X_BUF
    port map (
      I => addr2ext_0_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_1
    );
  tx_output_addr_Madd_n0000_inst_cy_1_263 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_15,
      IB => tx_output_addr_Madd_n0000_inst_cy_0,
      SEL => addr2ext_0_GROM,
      O => addr2ext_0_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_1 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_0,
      I1 => addr2ext_0_GROM,
      O => tx_output_addr_n0000(1)
    );
  addr2ext_2_LOGIC_ZERO_264 : X_ZERO
    port map (
      O => addr2ext_2_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_2_265 : X_MUX2
    port map (
      IA => addr2ext_2_LOGIC_ZERO,
      IB => addr2ext_2_CYINIT,
      SEL => addr2ext_2_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_2
    );
  tx_output_addr_Madd_n0000_inst_sum_2 : X_XOR2
    port map (
      I0 => addr2ext_2_CYINIT,
      I1 => addr2ext_2_FROM,
      O => tx_output_addr_n0000(2)
    );
  addr2ext_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(2),
      O => addr2ext_2_FROM
    );
  addr2ext_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(3),
      O => addr2ext_2_GROM
    );
  addr2ext_2_COUTUSED : X_BUF
    port map (
      I => addr2ext_2_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_3
    );
  tx_output_addr_Madd_n0000_inst_cy_3_266 : X_MUX2
    port map (
      IA => addr2ext_2_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_2,
      SEL => addr2ext_2_GROM,
      O => addr2ext_2_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_3 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_2,
      I1 => addr2ext_2_GROM,
      O => tx_output_addr_n0000(3)
    );
  addr2ext_2_CYINIT_267 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_1,
      O => addr2ext_2_CYINIT
    );
  addr2ext_4_LOGIC_ZERO_268 : X_ZERO
    port map (
      O => addr2ext_4_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_4_269 : X_MUX2
    port map (
      IA => addr2ext_4_LOGIC_ZERO,
      IB => addr2ext_4_CYINIT,
      SEL => addr2ext_4_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_4
    );
  tx_output_addr_Madd_n0000_inst_sum_4 : X_XOR2
    port map (
      I0 => addr2ext_4_CYINIT,
      I1 => addr2ext_4_FROM,
      O => tx_output_addr_n0000(4)
    );
  addr2ext_4_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr2ext(4),
      ADR3 => VCC,
      O => addr2ext_4_FROM
    );
  addr2ext_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr2ext(5),
      ADR3 => VCC,
      O => addr2ext_4_GROM
    );
  addr2ext_4_COUTUSED : X_BUF
    port map (
      I => addr2ext_4_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_5
    );
  tx_output_addr_Madd_n0000_inst_cy_5_270 : X_MUX2
    port map (
      IA => addr2ext_4_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_4,
      SEL => addr2ext_4_GROM,
      O => addr2ext_4_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_5 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_4,
      I1 => addr2ext_4_GROM,
      O => tx_output_addr_n0000(5)
    );
  addr2ext_4_CYINIT_271 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_3,
      O => addr2ext_4_CYINIT
    );
  addr2ext_6_LOGIC_ZERO_272 : X_ZERO
    port map (
      O => addr2ext_6_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_6_273 : X_MUX2
    port map (
      IA => addr2ext_6_LOGIC_ZERO,
      IB => addr2ext_6_CYINIT,
      SEL => addr2ext_6_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_6
    );
  tx_output_addr_Madd_n0000_inst_sum_6 : X_XOR2
    port map (
      I0 => addr2ext_6_CYINIT,
      I1 => addr2ext_6_FROM,
      O => tx_output_addr_n0000(6)
    );
  addr2ext_6_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(6),
      O => addr2ext_6_FROM
    );
  addr2ext_6_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(7),
      O => addr2ext_6_GROM
    );
  addr2ext_6_COUTUSED : X_BUF
    port map (
      I => addr2ext_6_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_7
    );
  tx_output_addr_Madd_n0000_inst_cy_7_274 : X_MUX2
    port map (
      IA => addr2ext_6_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_6,
      SEL => addr2ext_6_GROM,
      O => addr2ext_6_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_7 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_6,
      I1 => addr2ext_6_GROM,
      O => tx_output_addr_n0000(7)
    );
  addr2ext_6_CYINIT_275 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_5,
      O => addr2ext_6_CYINIT
    );
  addr2ext_8_LOGIC_ZERO_276 : X_ZERO
    port map (
      O => addr2ext_8_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_8_277 : X_MUX2
    port map (
      IA => addr2ext_8_LOGIC_ZERO,
      IB => addr2ext_8_CYINIT,
      SEL => addr2ext_8_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_8
    );
  tx_output_addr_Madd_n0000_inst_sum_8 : X_XOR2
    port map (
      I0 => addr2ext_8_CYINIT,
      I1 => addr2ext_8_FROM,
      O => tx_output_addr_n0000(8)
    );
  addr2ext_8_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr2ext(8),
      ADR3 => VCC,
      O => addr2ext_8_FROM
    );
  addr2ext_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr2ext(9),
      ADR3 => VCC,
      O => addr2ext_8_GROM
    );
  addr2ext_8_COUTUSED : X_BUF
    port map (
      I => addr2ext_8_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_9
    );
  tx_output_addr_Madd_n0000_inst_cy_9_278 : X_MUX2
    port map (
      IA => addr2ext_8_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_8,
      SEL => addr2ext_8_GROM,
      O => addr2ext_8_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_9 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_8,
      I1 => addr2ext_8_GROM,
      O => tx_output_addr_n0000(9)
    );
  addr2ext_8_CYINIT_279 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_7,
      O => addr2ext_8_CYINIT
    );
  addr2ext_10_LOGIC_ZERO_280 : X_ZERO
    port map (
      O => addr2ext_10_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_10_281 : X_MUX2
    port map (
      IA => addr2ext_10_LOGIC_ZERO,
      IB => addr2ext_10_CYINIT,
      SEL => addr2ext_10_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_10
    );
  tx_output_addr_Madd_n0000_inst_sum_10 : X_XOR2
    port map (
      I0 => addr2ext_10_CYINIT,
      I1 => addr2ext_10_FROM,
      O => tx_output_addr_n0000(10)
    );
  addr2ext_10_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(10),
      O => addr2ext_10_FROM
    );
  addr2ext_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(11),
      O => addr2ext_10_GROM
    );
  addr2ext_10_COUTUSED : X_BUF
    port map (
      I => addr2ext_10_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_11
    );
  tx_output_addr_Madd_n0000_inst_cy_11_282 : X_MUX2
    port map (
      IA => addr2ext_10_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_10,
      SEL => addr2ext_10_GROM,
      O => addr2ext_10_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_11 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_10,
      I1 => addr2ext_10_GROM,
      O => tx_output_addr_n0000(11)
    );
  addr2ext_10_CYINIT_283 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_9,
      O => addr2ext_10_CYINIT
    );
  addr2ext_12_LOGIC_ZERO_284 : X_ZERO
    port map (
      O => addr2ext_12_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_12_285 : X_MUX2
    port map (
      IA => addr2ext_12_LOGIC_ZERO,
      IB => addr2ext_12_CYINIT,
      SEL => addr2ext_12_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_12
    );
  tx_output_addr_Madd_n0000_inst_sum_12 : X_XOR2
    port map (
      I0 => addr2ext_12_CYINIT,
      I1 => addr2ext_12_FROM,
      O => tx_output_addr_n0000(12)
    );
  addr2ext_12_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => addr2ext(12),
      ADR3 => VCC,
      O => addr2ext_12_FROM
    );
  addr2ext_12_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(13),
      O => addr2ext_12_GROM
    );
  addr2ext_12_COUTUSED : X_BUF
    port map (
      I => addr2ext_12_CYMUXG,
      O => tx_output_addr_Madd_n0000_inst_cy_13
    );
  tx_output_addr_Madd_n0000_inst_cy_13_286 : X_MUX2
    port map (
      IA => addr2ext_12_LOGIC_ZERO,
      IB => tx_output_addr_Madd_n0000_inst_cy_12,
      SEL => addr2ext_12_GROM,
      O => addr2ext_12_CYMUXG
    );
  tx_output_addr_Madd_n0000_inst_sum_13 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_12,
      I1 => addr2ext_12_GROM,
      O => tx_output_addr_n0000(13)
    );
  addr2ext_12_CYINIT_287 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_11,
      O => addr2ext_12_CYINIT
    );
  addr2ext_14_LOGIC_ZERO_288 : X_ZERO
    port map (
      O => addr2ext_14_LOGIC_ZERO
    );
  tx_output_addr_Madd_n0000_inst_cy_14_289 : X_MUX2
    port map (
      IA => addr2ext_14_LOGIC_ZERO,
      IB => addr2ext_14_CYINIT,
      SEL => addr2ext_14_FROM,
      O => tx_output_addr_Madd_n0000_inst_cy_14
    );
  tx_output_addr_Madd_n0000_inst_sum_14 : X_XOR2
    port map (
      I0 => addr2ext_14_CYINIT,
      I1 => addr2ext_14_FROM,
      O => tx_output_addr_n0000(14)
    );
  addr2ext_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr2ext(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => addr2ext_14_FROM
    );
  addr2ext_15_rt_290 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => addr2ext(15),
      O => addr2ext_15_rt
    );
  tx_output_addr_Madd_n0000_inst_sum_15 : X_XOR2
    port map (
      I0 => tx_output_addr_Madd_n0000_inst_cy_14,
      I1 => addr2ext_15_rt,
      O => tx_output_addr_n0000(15)
    );
  addr2ext_14_CYINIT_291 : X_BUF
    port map (
      I => tx_output_addr_Madd_n0000_inst_cy_13,
      O => addr2ext_14_CYINIT
    );
  rx_input_memio_bcnt_86_LOGIC_ZERO_292 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_86_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_270_293 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_6,
      IB => rx_input_memio_bcnt_86_LOGIC_ZERO,
      SEL => rx_input_memio_cs_FFd16_2_rt,
      O => rx_input_memio_bcnt_inst_cy_270
    );
  rx_input_memio_cs_FFd16_2_rt_294 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_6,
      ADR1 => rx_input_memio_cs_FFd16_2,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_cs_FFd16_2_rt
    );
  rx_input_memio_bcnt_inst_lut3_721 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_3,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => rx_input_memio_bcnt_86,
      O => rx_input_memio_bcnt_inst_lut3_72
    );
  rx_input_memio_bcnt_86_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_86_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_271
    );
  rx_input_memio_bcnt_inst_cy_271_295 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_3,
      IB => rx_input_memio_bcnt_inst_cy_270,
      SEL => rx_input_memio_bcnt_inst_lut3_72,
      O => rx_input_memio_bcnt_86_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_235_296 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_270,
      I1 => rx_input_memio_bcnt_inst_lut3_72,
      O => rx_input_memio_bcnt_inst_sum_235
    );
  rx_input_memio_bcnt_87_LOGIC_ZERO_297 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_87_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_272_298 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_87_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_87_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_73,
      O => rx_input_memio_bcnt_inst_cy_272
    );
  rx_input_memio_bcnt_inst_sum_236_299 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_87_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_73,
      O => rx_input_memio_bcnt_inst_sum_236
    );
  rx_input_memio_bcnt_inst_lut3_731 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd16_1,
      ADR3 => rx_input_memio_bcnt_87,
      O => rx_input_memio_bcnt_inst_lut3_73
    );
  rx_input_memio_bcnt_inst_lut3_741 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcnt_88,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_74
    );
  rx_input_memio_bcnt_87_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_87_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_273
    );
  rx_input_memio_bcnt_87_YUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_87_XORG,
      O => rx_input_memio_bcnt_inst_sum_237
    );
  rx_input_memio_bcnt_inst_cy_273_300 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_87_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_272,
      SEL => rx_input_memio_bcnt_inst_lut3_74,
      O => rx_input_memio_bcnt_87_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_237_301 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_272,
      I1 => rx_input_memio_bcnt_inst_lut3_74,
      O => rx_input_memio_bcnt_87_XORG
    );
  rx_input_memio_bcnt_87_CYINIT_302 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_271,
      O => rx_input_memio_bcnt_87_CYINIT
    );
  rx_input_memio_bcnt_89_LOGIC_ZERO_303 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_89_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_274_304 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_89_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_89_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_75,
      O => rx_input_memio_bcnt_inst_cy_274
    );
  rx_input_memio_bcnt_inst_sum_238_305 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_89_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_75,
      O => rx_input_memio_bcnt_inst_sum_238
    );
  rx_input_memio_bcnt_inst_lut3_751 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => rx_input_memio_bcnt_89,
      O => rx_input_memio_bcnt_inst_lut3_75
    );
  rx_input_memio_bcnt_inst_lut3_761 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcnt_90,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_76
    );
  rx_input_memio_bcnt_89_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_89_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_275
    );
  rx_input_memio_bcnt_inst_cy_275_306 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_89_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_274,
      SEL => rx_input_memio_bcnt_inst_lut3_76,
      O => rx_input_memio_bcnt_89_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_239_307 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_274,
      I1 => rx_input_memio_bcnt_inst_lut3_76,
      O => rx_input_memio_bcnt_inst_sum_239
    );
  rx_input_memio_bcnt_89_CYINIT_308 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_273,
      O => rx_input_memio_bcnt_89_CYINIT
    );
  rx_input_memio_bcnt_91_LOGIC_ZERO_309 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_91_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_276_310 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_91_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_91_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_77,
      O => rx_input_memio_bcnt_inst_cy_276
    );
  rx_input_memio_bcnt_inst_sum_240_311 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_91_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_77,
      O => rx_input_memio_bcnt_inst_sum_240
    );
  rx_input_memio_bcnt_inst_lut3_771 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcnt_91,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_77
    );
  rx_input_memio_bcnt_inst_lut3_781 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcnt_92,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_78
    );
  rx_input_memio_bcnt_91_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_91_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_277
    );
  rx_input_memio_bcnt_inst_cy_277_312 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_91_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_276,
      SEL => rx_input_memio_bcnt_inst_lut3_78,
      O => rx_input_memio_bcnt_91_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_241_313 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_276,
      I1 => rx_input_memio_bcnt_inst_lut3_78,
      O => rx_input_memio_bcnt_inst_sum_241
    );
  rx_input_memio_bcnt_91_CYINIT_314 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_275,
      O => rx_input_memio_bcnt_91_CYINIT
    );
  rx_input_memio_bcnt_93_LOGIC_ZERO_315 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_93_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_278_316 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_93_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_93_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_79,
      O => rx_input_memio_bcnt_inst_cy_278
    );
  rx_input_memio_bcnt_inst_sum_242_317 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_93_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_79,
      O => rx_input_memio_bcnt_inst_sum_242
    );
  rx_input_memio_bcnt_inst_lut3_791 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcnt_93,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_79
    );
  rx_input_memio_bcnt_inst_lut3_801 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bcnt_94,
      O => rx_input_memio_bcnt_inst_lut3_80
    );
  rx_input_memio_bcnt_93_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_93_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_279
    );
  rx_input_memio_bcnt_inst_cy_279_318 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_93_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_278,
      SEL => rx_input_memio_bcnt_inst_lut3_80,
      O => rx_input_memio_bcnt_93_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_243_319 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_278,
      I1 => rx_input_memio_bcnt_inst_lut3_80,
      O => rx_input_memio_bcnt_inst_sum_243
    );
  rx_input_memio_bcnt_93_CYINIT_320 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_277,
      O => rx_input_memio_bcnt_93_CYINIT
    );
  rx_input_memio_dout_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_3_FFX_RST,
      O => rx_input_memio_dout(3)
    );
  rx_input_memio_dout_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_3_FFX_RST
    );
  rx_input_memio_bcnt_95_LOGIC_ZERO_321 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_95_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_280_322 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_95_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_95_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_81,
      O => rx_input_memio_bcnt_inst_cy_280
    );
  rx_input_memio_bcnt_inst_sum_244_323 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_95_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_81,
      O => rx_input_memio_bcnt_inst_sum_244
    );
  rx_input_memio_bcnt_inst_lut3_811 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bcnt_95,
      O => rx_input_memio_bcnt_inst_lut3_81
    );
  rx_input_memio_bcnt_inst_lut3_821 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcnt_96,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_82
    );
  rx_input_memio_bcnt_95_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_95_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_281
    );
  rx_input_memio_bcnt_inst_cy_281_324 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_95_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_280,
      SEL => rx_input_memio_bcnt_inst_lut3_82,
      O => rx_input_memio_bcnt_95_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_245_325 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_280,
      I1 => rx_input_memio_bcnt_inst_lut3_82,
      O => rx_input_memio_bcnt_inst_sum_245
    );
  rx_input_memio_bcnt_95_CYINIT_326 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_279,
      O => rx_input_memio_bcnt_95_CYINIT
    );
  rx_input_memio_bcnt_97_LOGIC_ZERO_327 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_97_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_282_328 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_97_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_97_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_83,
      O => rx_input_memio_bcnt_inst_cy_282
    );
  rx_input_memio_bcnt_inst_sum_246_329 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_97_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_83,
      O => rx_input_memio_bcnt_inst_sum_246
    );
  rx_input_memio_bcnt_inst_lut3_831 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcnt_97,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_83
    );
  rx_input_memio_bcnt_inst_lut3_841 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => rx_input_memio_bcnt_98,
      ADR3 => VCC,
      O => rx_input_memio_bcnt_inst_lut3_84
    );
  rx_input_memio_bcnt_97_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_97_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_283
    );
  rx_input_memio_bcnt_inst_cy_283_330 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_97_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_282,
      SEL => rx_input_memio_bcnt_inst_lut3_84,
      O => rx_input_memio_bcnt_97_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_247_331 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_282,
      I1 => rx_input_memio_bcnt_inst_lut3_84,
      O => rx_input_memio_bcnt_inst_sum_247
    );
  rx_input_memio_bcnt_97_CYINIT_332 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_281,
      O => rx_input_memio_bcnt_97_CYINIT
    );
  rx_input_memio_bcnt_99_LOGIC_ZERO_333 : X_ZERO
    port map (
      O => rx_input_memio_bcnt_99_LOGIC_ZERO
    );
  rx_input_memio_bcnt_inst_cy_284_334 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_99_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_99_CYINIT,
      SEL => rx_input_memio_bcnt_inst_lut3_85,
      O => rx_input_memio_bcnt_inst_cy_284
    );
  rx_input_memio_bcnt_inst_sum_248_335 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_99_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_85,
      O => rx_input_memio_bcnt_inst_sum_248
    );
  rx_input_memio_bcnt_inst_lut3_851 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_99,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_85
    );
  rx_input_memio_bcnt_inst_lut3_861 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd16,
      ADR3 => rx_input_memio_bcnt_100,
      O => rx_input_memio_bcnt_inst_lut3_86
    );
  rx_input_memio_bcnt_99_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcnt_99_CYMUXG,
      O => rx_input_memio_bcnt_inst_cy_285
    );
  rx_input_memio_bcnt_inst_cy_285_336 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_99_LOGIC_ZERO,
      IB => rx_input_memio_bcnt_inst_cy_284,
      SEL => rx_input_memio_bcnt_inst_lut3_86,
      O => rx_input_memio_bcnt_99_CYMUXG
    );
  rx_input_memio_bcnt_inst_sum_249_337 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_inst_cy_284,
      I1 => rx_input_memio_bcnt_inst_lut3_86,
      O => rx_input_memio_bcnt_inst_sum_249
    );
  rx_input_memio_bcnt_99_CYINIT_338 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_283,
      O => rx_input_memio_bcnt_99_CYINIT
    );
  rx_input_memio_bcnt_inst_sum_250_339 : X_XOR2
    port map (
      I0 => rx_input_memio_bcnt_101_CYINIT,
      I1 => rx_input_memio_bcnt_inst_lut3_87,
      O => rx_input_memio_bcnt_inst_sum_250
    );
  rx_input_memio_bcnt_inst_lut3_871 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcnt_101,
      ADR3 => rx_input_memio_cs_FFd16,
      O => rx_input_memio_bcnt_inst_lut3_87
    );
  rx_input_memio_bcnt_101_CYINIT_340 : X_BUF
    port map (
      I => rx_input_memio_bcnt_inst_cy_285,
      O => rx_input_memio_bcnt_101_CYINIT
    );
  rx_output_Madd_n0060_inst_cy_49_LOGIC_ZERO_341 : X_ZERO
    port map (
      O => rx_output_Madd_n0060_inst_cy_49_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_48_342 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_17,
      IB => rx_output_Madd_n0060_inst_cy_49_LOGIC_ZERO,
      SEL => rx_output_Madd_n0060_inst_lut2_4811_O,
      O => rx_output_Madd_n0060_inst_cy_48
    );
  rx_output_Madd_n0060_inst_lut2_4811 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_17,
      ADR1 => VCC,
      ADR2 => rx_output_len(0),
      ADR3 => VCC,
      O => rx_output_Madd_n0060_inst_lut2_4811_O
    );
  rx_output_Madd_n0060_inst_lut2_491 : X_LUT4
    generic map(
      INIT => X"EEEE"
    )
    port map (
      ADR0 => rx_output_len(1),
      ADR1 => rx_output_len(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_Madd_n0060_inst_lut2_491_O
    );
  rx_output_Madd_n0060_inst_cy_49_COUTUSED : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_49_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_49
    );
  rx_output_Madd_n0060_inst_cy_49_343 : X_MUX2
    port map (
      IA => rx_output_len(1),
      IB => rx_output_Madd_n0060_inst_cy_48,
      SEL => rx_output_Madd_n0060_inst_lut2_491_O,
      O => rx_output_Madd_n0060_inst_cy_49_CYMUXG
    );
  rx_output_n0060_2_LOGIC_ZERO_344 : X_ZERO
    port map (
      O => rx_output_n0060_2_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_50_345 : X_MUX2
    port map (
      IA => rx_output_n0060_2_LOGIC_ZERO,
      IB => rx_output_n0060_2_CYINIT,
      SEL => rx_output_n0060_2_FROM,
      O => rx_output_Madd_n0060_inst_cy_50
    );
  rx_output_Madd_n0060_inst_sum_50 : X_XOR2
    port map (
      I0 => rx_output_n0060_2_CYINIT,
      I1 => rx_output_n0060_2_FROM,
      O => rx_output_n0060_2_XORF
    );
  rx_output_n0060_2_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(2),
      ADR3 => VCC,
      O => rx_output_n0060_2_FROM
    );
  rx_output_n0060_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(3),
      O => rx_output_n0060_2_GROM
    );
  rx_output_n0060_2_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_2_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_51
    );
  rx_output_n0060_2_XUSED : X_BUF
    port map (
      I => rx_output_n0060_2_XORF,
      O => rx_output_n0060(2)
    );
  rx_output_n0060_2_YUSED : X_BUF
    port map (
      I => rx_output_n0060_2_XORG,
      O => rx_output_n0060(3)
    );
  rx_output_Madd_n0060_inst_cy_51_346 : X_MUX2
    port map (
      IA => rx_output_n0060_2_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_50,
      SEL => rx_output_n0060_2_GROM,
      O => rx_output_n0060_2_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_51 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_50,
      I1 => rx_output_n0060_2_GROM,
      O => rx_output_n0060_2_XORG
    );
  rx_output_n0060_2_CYINIT_347 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_49,
      O => rx_output_n0060_2_CYINIT
    );
  rx_output_n0060_4_LOGIC_ZERO_348 : X_ZERO
    port map (
      O => rx_output_n0060_4_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_52_349 : X_MUX2
    port map (
      IA => rx_output_n0060_4_LOGIC_ZERO,
      IB => rx_output_n0060_4_CYINIT,
      SEL => rx_output_n0060_4_FROM,
      O => rx_output_Madd_n0060_inst_cy_52
    );
  rx_output_Madd_n0060_inst_sum_52 : X_XOR2
    port map (
      I0 => rx_output_n0060_4_CYINIT,
      I1 => rx_output_n0060_4_FROM,
      O => rx_output_n0060_4_XORF
    );
  rx_output_n0060_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_4_FROM
    );
  rx_output_n0060_4_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(5),
      O => rx_output_n0060_4_GROM
    );
  rx_output_n0060_4_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_4_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_53
    );
  rx_output_n0060_4_XUSED : X_BUF
    port map (
      I => rx_output_n0060_4_XORF,
      O => rx_output_n0060(4)
    );
  rx_output_n0060_4_YUSED : X_BUF
    port map (
      I => rx_output_n0060_4_XORG,
      O => rx_output_n0060(5)
    );
  rx_output_Madd_n0060_inst_cy_53_350 : X_MUX2
    port map (
      IA => rx_output_n0060_4_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_52,
      SEL => rx_output_n0060_4_GROM,
      O => rx_output_n0060_4_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_53 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_52,
      I1 => rx_output_n0060_4_GROM,
      O => rx_output_n0060_4_XORG
    );
  rx_output_n0060_4_CYINIT_351 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_51,
      O => rx_output_n0060_4_CYINIT
    );
  rx_input_memio_dout_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_5_FFY_RST,
      O => rx_input_memio_dout(4)
    );
  rx_input_memio_dout_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_5_FFY_RST
    );
  rx_output_n0060_6_LOGIC_ZERO_352 : X_ZERO
    port map (
      O => rx_output_n0060_6_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_54_353 : X_MUX2
    port map (
      IA => rx_output_n0060_6_LOGIC_ZERO,
      IB => rx_output_n0060_6_CYINIT,
      SEL => rx_output_n0060_6_FROM,
      O => rx_output_Madd_n0060_inst_cy_54
    );
  rx_output_Madd_n0060_inst_sum_54 : X_XOR2
    port map (
      I0 => rx_output_n0060_6_CYINIT,
      I1 => rx_output_n0060_6_FROM,
      O => rx_output_n0060_6_XORF
    );
  rx_output_n0060_6_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_6_FROM
    );
  rx_output_n0060_6_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(7),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_6_GROM
    );
  rx_output_n0060_6_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_6_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_55
    );
  rx_output_n0060_6_XUSED : X_BUF
    port map (
      I => rx_output_n0060_6_XORF,
      O => rx_output_n0060(6)
    );
  rx_output_n0060_6_YUSED : X_BUF
    port map (
      I => rx_output_n0060_6_XORG,
      O => rx_output_n0060(7)
    );
  rx_output_Madd_n0060_inst_cy_55_354 : X_MUX2
    port map (
      IA => rx_output_n0060_6_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_54,
      SEL => rx_output_n0060_6_GROM,
      O => rx_output_n0060_6_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_55 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_54,
      I1 => rx_output_n0060_6_GROM,
      O => rx_output_n0060_6_XORG
    );
  rx_output_n0060_6_CYINIT_355 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_53,
      O => rx_output_n0060_6_CYINIT
    );
  rx_output_n0060_8_LOGIC_ZERO_356 : X_ZERO
    port map (
      O => rx_output_n0060_8_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_56_357 : X_MUX2
    port map (
      IA => rx_output_n0060_8_LOGIC_ZERO,
      IB => rx_output_n0060_8_CYINIT,
      SEL => rx_output_n0060_8_FROM,
      O => rx_output_Madd_n0060_inst_cy_56
    );
  rx_output_Madd_n0060_inst_sum_56 : X_XOR2
    port map (
      I0 => rx_output_n0060_8_CYINIT,
      I1 => rx_output_n0060_8_FROM,
      O => rx_output_n0060_8_XORF
    );
  rx_output_n0060_8_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_8_FROM
    );
  rx_output_n0060_8_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(9),
      O => rx_output_n0060_8_GROM
    );
  rx_output_n0060_8_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_8_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_57
    );
  rx_output_n0060_8_XUSED : X_BUF
    port map (
      I => rx_output_n0060_8_XORF,
      O => rx_output_n0060(8)
    );
  rx_output_n0060_8_YUSED : X_BUF
    port map (
      I => rx_output_n0060_8_XORG,
      O => rx_output_n0060(9)
    );
  rx_output_Madd_n0060_inst_cy_57_358 : X_MUX2
    port map (
      IA => rx_output_n0060_8_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_56,
      SEL => rx_output_n0060_8_GROM,
      O => rx_output_n0060_8_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_57 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_56,
      I1 => rx_output_n0060_8_GROM,
      O => rx_output_n0060_8_XORG
    );
  rx_output_n0060_8_CYINIT_359 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_55,
      O => rx_output_n0060_8_CYINIT
    );
  rx_output_n0060_10_LOGIC_ZERO_360 : X_ZERO
    port map (
      O => rx_output_n0060_10_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_58_361 : X_MUX2
    port map (
      IA => rx_output_n0060_10_LOGIC_ZERO,
      IB => rx_output_n0060_10_CYINIT,
      SEL => rx_output_n0060_10_FROM,
      O => rx_output_Madd_n0060_inst_cy_58
    );
  rx_output_Madd_n0060_inst_sum_58 : X_XOR2
    port map (
      I0 => rx_output_n0060_10_CYINIT,
      I1 => rx_output_n0060_10_FROM,
      O => rx_output_n0060_10_XORF
    );
  rx_output_n0060_10_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(10),
      ADR3 => VCC,
      O => rx_output_n0060_10_FROM
    );
  rx_output_n0060_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(11),
      O => rx_output_n0060_10_GROM
    );
  rx_output_n0060_10_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_10_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_59
    );
  rx_output_n0060_10_XUSED : X_BUF
    port map (
      I => rx_output_n0060_10_XORF,
      O => rx_output_n0060(10)
    );
  rx_output_n0060_10_YUSED : X_BUF
    port map (
      I => rx_output_n0060_10_XORG,
      O => rx_output_n0060(11)
    );
  rx_output_Madd_n0060_inst_cy_59_362 : X_MUX2
    port map (
      IA => rx_output_n0060_10_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_58,
      SEL => rx_output_n0060_10_GROM,
      O => rx_output_n0060_10_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_59 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_58,
      I1 => rx_output_n0060_10_GROM,
      O => rx_output_n0060_10_XORG
    );
  rx_output_n0060_10_CYINIT_363 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_57,
      O => rx_output_n0060_10_CYINIT
    );
  rx_output_n0060_12_LOGIC_ZERO_364 : X_ZERO
    port map (
      O => rx_output_n0060_12_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_60_365 : X_MUX2
    port map (
      IA => rx_output_n0060_12_LOGIC_ZERO,
      IB => rx_output_n0060_12_CYINIT,
      SEL => rx_output_n0060_12_FROM,
      O => rx_output_Madd_n0060_inst_cy_60
    );
  rx_output_Madd_n0060_inst_sum_60 : X_XOR2
    port map (
      I0 => rx_output_n0060_12_CYINIT,
      I1 => rx_output_n0060_12_FROM,
      O => rx_output_n0060_12_XORF
    );
  rx_output_n0060_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_12_FROM
    );
  rx_output_n0060_12_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(13),
      ADR3 => VCC,
      O => rx_output_n0060_12_GROM
    );
  rx_output_n0060_12_COUTUSED : X_BUF
    port map (
      I => rx_output_n0060_12_CYMUXG,
      O => rx_output_Madd_n0060_inst_cy_61
    );
  rx_output_n0060_12_XUSED : X_BUF
    port map (
      I => rx_output_n0060_12_XORF,
      O => rx_output_n0060(12)
    );
  rx_output_n0060_12_YUSED : X_BUF
    port map (
      I => rx_output_n0060_12_XORG,
      O => rx_output_n0060(13)
    );
  rx_output_Madd_n0060_inst_cy_61_366 : X_MUX2
    port map (
      IA => rx_output_n0060_12_LOGIC_ZERO,
      IB => rx_output_Madd_n0060_inst_cy_60,
      SEL => rx_output_n0060_12_GROM,
      O => rx_output_n0060_12_CYMUXG
    );
  rx_output_Madd_n0060_inst_sum_61 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_60,
      I1 => rx_output_n0060_12_GROM,
      O => rx_output_n0060_12_XORG
    );
  rx_output_n0060_12_CYINIT_367 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_59,
      O => rx_output_n0060_12_CYINIT
    );
  tx_output_FBBP_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(13),
      CE => txfbbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_13_FFX_RST,
      O => txfbbp(13)
    );
  txfbbp_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_13_FFX_RST
    );
  rx_output_n0060_14_LOGIC_ZERO_368 : X_ZERO
    port map (
      O => rx_output_n0060_14_LOGIC_ZERO
    );
  rx_output_Madd_n0060_inst_cy_62_369 : X_MUX2
    port map (
      IA => rx_output_n0060_14_LOGIC_ZERO,
      IB => rx_output_n0060_14_CYINIT,
      SEL => rx_output_n0060_14_FROM,
      O => rx_output_Madd_n0060_inst_cy_62
    );
  rx_output_Madd_n0060_inst_sum_62 : X_XOR2
    port map (
      I0 => rx_output_n0060_14_CYINIT,
      I1 => rx_output_n0060_14_FROM,
      O => rx_output_n0060_14_XORF
    );
  rx_output_n0060_14_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(14),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0060_14_FROM
    );
  rx_output_len_15_rt_370 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(15),
      O => rx_output_len_15_rt
    );
  rx_output_n0060_14_XUSED : X_BUF
    port map (
      I => rx_output_n0060_14_XORF,
      O => rx_output_n0060(14)
    );
  rx_output_n0060_14_YUSED : X_BUF
    port map (
      I => rx_output_n0060_14_XORG,
      O => rx_output_n0060(15)
    );
  rx_output_Madd_n0060_inst_sum_63 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0060_inst_cy_62,
      I1 => rx_output_len_15_rt,
      O => rx_output_n0060_14_XORG
    );
  rx_output_n0060_14_CYINIT_371 : X_BUF
    port map (
      I => rx_output_Madd_n0060_inst_cy_61,
      O => rx_output_n0060_14_CYINIT
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ONE_372 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ZERO_373 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_177_374 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(9),
      ADR1 => rx_input_memio_addrchk_datal(8),
      ADR2 => rx_input_memio_addrchk_macaddrl(9),
      ADR3 => rx_input_memio_addrchk_macaddrl(8),
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(11),
      ADR1 => rx_input_memio_addrchk_macaddrl(10),
      ADR2 => rx_input_memio_addrchk_datal(11),
      ADR3 => rx_input_memio_addrchk_datal(10),
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_375 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_4_LOGIC_ZERO_376 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_4_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_179_377 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_4_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_4_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(12),
      ADR1 => rx_input_memio_addrchk_macaddrl(13),
      ADR2 => rx_input_memio_addrchk_datal(13),
      ADR3 => rx_input_memio_addrchk_macaddrl(12),
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(14),
      ADR1 => rx_input_memio_addrchk_macaddrl(15),
      ADR2 => rx_input_memio_addrchk_datal(15),
      ADR3 => rx_input_memio_addrchk_datal(14),
      O => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_4_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_4_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(4)
    );
  rx_input_memio_addrchk_Mcompar_n0036_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_4_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0036_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_4_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_4_CYINIT_378 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0036_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_4_CYINIT
    );
  mac_control_rxcrcerr_cnt_0_LOGIC_ZERO_379 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_0_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_16_380 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_28,
      IB => mac_control_rxcrcerr_cnt_0_LOGIC_ZERO,
      SEL => mac_control_rxcrcerr_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_28,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(0),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_rxcrcerr_cnt_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_42,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(1),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_0_GROM
    );
  mac_control_rxcrcerr_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_0_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_17_381 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_42,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_rxcrcerr_cnt_0_GROM,
      O => mac_control_rxcrcerr_cnt_0_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_rxcrcerr_cnt_0_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(1)
    );
  mac_control_rxcrcerr_cnt_2_LOGIC_ZERO_382 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_2_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_18_383 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_2_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_2_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_2_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_2_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(2)
    );
  mac_control_rxcrcerr_cnt_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(2),
      O => mac_control_rxcrcerr_cnt_2_FROM
    );
  mac_control_rxcrcerr_cnt_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(3),
      O => mac_control_rxcrcerr_cnt_2_GROM
    );
  mac_control_rxcrcerr_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_2_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_19_384 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_rxcrcerr_cnt_2_GROM,
      O => mac_control_rxcrcerr_cnt_2_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_rxcrcerr_cnt_2_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(3)
    );
  mac_control_rxcrcerr_cnt_2_CYINIT_385 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_rxcrcerr_cnt_2_CYINIT
    );
  mac_control_rxcrcerr_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(5),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(5)
    );
  mac_control_rxcrcerr_cnt_4_LOGIC_ZERO_386 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_4_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_20_387 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_4_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_4_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_4_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_4_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(4)
    );
  mac_control_rxcrcerr_cnt_4_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(4),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_4_FROM
    );
  mac_control_rxcrcerr_cnt_4_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxcrcerr_cnt(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_4_GROM
    );
  mac_control_rxcrcerr_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_4_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_21_388 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_rxcrcerr_cnt_4_GROM,
      O => mac_control_rxcrcerr_cnt_4_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_rxcrcerr_cnt_4_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(5)
    );
  mac_control_rxcrcerr_cnt_4_CYINIT_389 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_rxcrcerr_cnt_4_CYINIT
    );
  mac_control_rxcrcerr_cnt_6_LOGIC_ZERO_390 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_6_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_22_391 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_6_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_6_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_6_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_6_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(6)
    );
  mac_control_rxcrcerr_cnt_6_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(6),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_6_FROM
    );
  mac_control_rxcrcerr_cnt_6_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(7),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_6_GROM
    );
  mac_control_rxcrcerr_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_6_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_23_392 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_rxcrcerr_cnt_6_GROM,
      O => mac_control_rxcrcerr_cnt_6_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_rxcrcerr_cnt_6_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(7)
    );
  mac_control_rxcrcerr_cnt_6_CYINIT_393 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_rxcrcerr_cnt_6_CYINIT
    );
  mac_control_rxcrcerr_cnt_8_LOGIC_ZERO_394 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_8_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_24_395 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_8_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_8_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_8_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_8_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(8)
    );
  mac_control_rxcrcerr_cnt_8_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(8),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_8_FROM
    );
  mac_control_rxcrcerr_cnt_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(9),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_8_GROM
    );
  mac_control_rxcrcerr_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_8_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_25_396 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_rxcrcerr_cnt_8_GROM,
      O => mac_control_rxcrcerr_cnt_8_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_rxcrcerr_cnt_8_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(9)
    );
  mac_control_rxcrcerr_cnt_8_CYINIT_397 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_rxcrcerr_cnt_8_CYINIT
    );
  mac_control_rxcrcerr_cnt_10_LOGIC_ZERO_398 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_10_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_26_399 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_10_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_10_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_10_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_10_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(10)
    );
  mac_control_rxcrcerr_cnt_10_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(10),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_10_FROM
    );
  mac_control_rxcrcerr_cnt_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(11),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_10_GROM
    );
  mac_control_rxcrcerr_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_10_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_27_400 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_rxcrcerr_cnt_10_GROM,
      O => mac_control_rxcrcerr_cnt_10_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_rxcrcerr_cnt_10_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(11)
    );
  mac_control_rxcrcerr_cnt_10_CYINIT_401 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_rxcrcerr_cnt_10_CYINIT
    );
  mac_control_rxcrcerr_cnt_12_LOGIC_ZERO_402 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_12_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_28_403 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_12_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_12_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_12_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_12_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(12)
    );
  mac_control_rxcrcerr_cnt_12_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(12),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_12_FROM
    );
  mac_control_rxcrcerr_cnt_12_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxcrcerr_cnt(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_12_GROM
    );
  mac_control_rxcrcerr_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_12_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_29_404 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_rxcrcerr_cnt_12_GROM,
      O => mac_control_rxcrcerr_cnt_12_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_rxcrcerr_cnt_12_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(13)
    );
  mac_control_rxcrcerr_cnt_12_CYINIT_405 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_rxcrcerr_cnt_12_CYINIT
    );
  mac_control_rxcrcerr_cnt_14_LOGIC_ZERO_406 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_14_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_30_407 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_14_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_14_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_14_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_14_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(14)
    );
  mac_control_rxcrcerr_cnt_14_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(14),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_14_FROM
    );
  mac_control_rxcrcerr_cnt_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(15),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_14_GROM
    );
  mac_control_rxcrcerr_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_14_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_31_408 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_rxcrcerr_cnt_14_GROM,
      O => mac_control_rxcrcerr_cnt_14_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_rxcrcerr_cnt_14_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(15)
    );
  mac_control_rxcrcerr_cnt_14_CYINIT_409 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_rxcrcerr_cnt_14_CYINIT
    );
  mac_control_rxcrcerr_cnt_16_LOGIC_ZERO_410 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_16_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_32_411 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_16_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_16_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_16_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_16_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(16)
    );
  mac_control_rxcrcerr_cnt_16_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxcrcerr_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_16_FROM
    );
  mac_control_rxcrcerr_cnt_16_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(17),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_16_GROM
    );
  mac_control_rxcrcerr_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_16_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_33_412 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_rxcrcerr_cnt_16_GROM,
      O => mac_control_rxcrcerr_cnt_16_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_rxcrcerr_cnt_16_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(17)
    );
  mac_control_rxcrcerr_cnt_16_CYINIT_413 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_rxcrcerr_cnt_16_CYINIT
    );
  mac_control_rxcrcerr_cnt_18_LOGIC_ZERO_414 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_18_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_34_415 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_18_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_18_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_18_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_18_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(18)
    );
  mac_control_rxcrcerr_cnt_18_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(18),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_18_FROM
    );
  mac_control_rxcrcerr_cnt_18_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(19),
      O => mac_control_rxcrcerr_cnt_18_GROM
    );
  mac_control_rxcrcerr_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_18_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_35_416 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_rxcrcerr_cnt_18_GROM,
      O => mac_control_rxcrcerr_cnt_18_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_rxcrcerr_cnt_18_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(19)
    );
  mac_control_rxcrcerr_cnt_18_CYINIT_417 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_rxcrcerr_cnt_18_CYINIT
    );
  rx_input_memio_dout_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_5_FFX_RST,
      O => rx_input_memio_dout(5)
    );
  rx_input_memio_dout_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_5_FFX_RST
    );
  mac_control_rxcrcerr_cnt_20_LOGIC_ZERO_418 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_20_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_36_419 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_20_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_20_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_20_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_20_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(20)
    );
  mac_control_rxcrcerr_cnt_20_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(20),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_20_FROM
    );
  mac_control_rxcrcerr_cnt_20_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(21),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_20_GROM
    );
  mac_control_rxcrcerr_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_20_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_37_420 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_rxcrcerr_cnt_20_GROM,
      O => mac_control_rxcrcerr_cnt_20_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_rxcrcerr_cnt_20_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(21)
    );
  mac_control_rxcrcerr_cnt_20_CYINIT_421 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_rxcrcerr_cnt_20_CYINIT
    );
  mac_control_rxcrcerr_cnt_22_LOGIC_ZERO_422 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_22_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_38_423 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_22_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_22_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_22_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_22_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(22)
    );
  mac_control_rxcrcerr_cnt_22_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(22),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_22_FROM
    );
  mac_control_rxcrcerr_cnt_22_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(23),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_22_GROM
    );
  mac_control_rxcrcerr_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_22_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_39_424 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_rxcrcerr_cnt_22_GROM,
      O => mac_control_rxcrcerr_cnt_22_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_rxcrcerr_cnt_22_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(23)
    );
  mac_control_rxcrcerr_cnt_22_CYINIT_425 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_rxcrcerr_cnt_22_CYINIT
    );
  mac_control_rxcrcerr_cnt_24_LOGIC_ZERO_426 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_24_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_40_427 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_24_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_24_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_24_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_24_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(24)
    );
  mac_control_rxcrcerr_cnt_24_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(24),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_24_FROM
    );
  mac_control_rxcrcerr_cnt_24_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(25),
      O => mac_control_rxcrcerr_cnt_24_GROM
    );
  mac_control_rxcrcerr_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_24_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_41_428 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_rxcrcerr_cnt_24_GROM,
      O => mac_control_rxcrcerr_cnt_24_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_rxcrcerr_cnt_24_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(25)
    );
  mac_control_rxcrcerr_cnt_24_CYINIT_429 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_rxcrcerr_cnt_24_CYINIT
    );
  mac_control_rxcrcerr_cnt_26_LOGIC_ZERO_430 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_26_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_42_431 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_26_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_26_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_26_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_26_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(26)
    );
  mac_control_rxcrcerr_cnt_26_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(26),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_26_FROM
    );
  mac_control_rxcrcerr_cnt_26_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(27),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_26_GROM
    );
  mac_control_rxcrcerr_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_26_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_43_432 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_rxcrcerr_cnt_26_GROM,
      O => mac_control_rxcrcerr_cnt_26_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_rxcrcerr_cnt_26_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(27)
    );
  mac_control_rxcrcerr_cnt_26_CYINIT_433 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_rxcrcerr_cnt_26_CYINIT
    );
  mac_control_rxcrcerr_cnt_28_LOGIC_ZERO_434 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_28_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_44_435 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_28_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_28_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_28_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_28_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(28)
    );
  mac_control_rxcrcerr_cnt_28_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxcrcerr_cnt(28),
      O => mac_control_rxcrcerr_cnt_28_FROM
    );
  mac_control_rxcrcerr_cnt_28_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(29),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_28_GROM
    );
  mac_control_rxcrcerr_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_28_CYMUXG,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_45_436 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_rxcrcerr_cnt_28_GROM,
      O => mac_control_rxcrcerr_cnt_28_CYMUXG
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_rxcrcerr_cnt_28_GROM,
      O => mac_control_rxcrcerr_cnt_n0000(29)
    );
  mac_control_rxcrcerr_cnt_28_CYINIT_437 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_rxcrcerr_cnt_28_CYINIT
    );
  mac_control_rxcrcerr_cnt_30_LOGIC_ZERO_438 : X_ZERO
    port map (
      O => mac_control_rxcrcerr_cnt_30_LOGIC_ZERO
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_46_439 : X_MUX2
    port map (
      IA => mac_control_rxcrcerr_cnt_30_LOGIC_ZERO,
      IB => mac_control_rxcrcerr_cnt_30_CYINIT,
      SEL => mac_control_rxcrcerr_cnt_30_FROM,
      O => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_30_CYINIT,
      I1 => mac_control_rxcrcerr_cnt_30_FROM,
      O => mac_control_rxcrcerr_cnt_n0000(30)
    );
  mac_control_rxcrcerr_cnt_30_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(30),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_30_FROM
    );
  mac_control_rxcrcerr_cnt_31_rt_440 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxcrcerr_cnt(31),
      ADR3 => VCC,
      O => mac_control_rxcrcerr_cnt_31_rt
    );
  mac_control_rxcrcerr_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_rxcrcerr_cnt_31_rt,
      O => mac_control_rxcrcerr_cnt_n0000(31)
    );
  mac_control_rxcrcerr_cnt_30_CYINIT_441 : X_BUF
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_rxcrcerr_cnt_30_CYINIT
    );
  rx_input_memio_bp_0_LOGIC_ONE_442 : X_ONE
    port map (
      O => rx_input_memio_bp_0_LOGIC_ONE
    );
  rx_input_memio_Msub_n0043_inst_cy_221_443 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_0,
      IB => rx_input_memio_bp_0_CYINIT,
      SEL => rx_input_memio_bp_0_FROM,
      O => rx_input_memio_Msub_n0043_inst_cy_221
    );
  rx_input_memio_Msub_n0043_inst_sum_187 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_0_CYINIT,
      I1 => rx_input_memio_bp_0_FROM,
      O => rx_input_memio_n0043(0)
    );
  rx_input_memio_bp_0_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_0,
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_70,
      ADR3 => VCC,
      O => rx_input_memio_bp_0_FROM
    );
  rx_input_memio_Msub_n0043_inst_lut2_1341 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_71,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_134
    );
  rx_input_memio_bp_0_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_0_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_222
    );
  rx_input_memio_Msub_n0043_inst_cy_222_444 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_71,
      IB => rx_input_memio_Msub_n0043_inst_cy_221,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_134,
      O => rx_input_memio_bp_0_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_188 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_221,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_134,
      O => rx_input_memio_n0043(1)
    );
  rx_input_memio_bp_0_CYINIT_445 : X_BUF
    port map (
      I => rx_input_memio_bp_0_LOGIC_ONE,
      O => rx_input_memio_bp_0_CYINIT
    );
  rx_input_memio_bp_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_2_FFY_RST
    );
  rx_input_memio_bp_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(3),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_2_FFY_RST,
      O => rx_input_memio_bp(3)
    );
  rx_input_memio_Msub_n0043_inst_cy_223_446 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_72,
      IB => rx_input_memio_bp_2_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_135,
      O => rx_input_memio_Msub_n0043_inst_cy_223
    );
  rx_input_memio_Msub_n0043_inst_sum_189 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_2_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_135,
      O => rx_input_memio_n0043(2)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1351 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_72,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_135
    );
  rx_input_memio_Msub_n0043_inst_lut2_1361 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_73,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_136
    );
  rx_input_memio_bp_2_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_2_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_224
    );
  rx_input_memio_Msub_n0043_inst_cy_224_447 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_73,
      IB => rx_input_memio_Msub_n0043_inst_cy_223,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_136,
      O => rx_input_memio_bp_2_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_190 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_223,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_136,
      O => rx_input_memio_n0043(3)
    );
  rx_input_memio_bp_2_CYINIT_448 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_222,
      O => rx_input_memio_bp_2_CYINIT
    );
  rx_input_memio_bp_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_4_FFY_RST
    );
  rx_input_memio_bp_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(5),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_4_FFY_RST,
      O => rx_input_memio_bp(5)
    );
  rx_input_memio_Msub_n0043_inst_cy_225_449 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_74,
      IB => rx_input_memio_bp_4_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_137,
      O => rx_input_memio_Msub_n0043_inst_cy_225
    );
  rx_input_memio_Msub_n0043_inst_sum_191 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_4_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_137,
      O => rx_input_memio_n0043(4)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1371 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_74,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_137
    );
  rx_input_memio_Msub_n0043_inst_lut2_1381 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_75,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_138
    );
  rx_input_memio_bp_4_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_4_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_226
    );
  rx_input_memio_Msub_n0043_inst_cy_226_450 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_75,
      IB => rx_input_memio_Msub_n0043_inst_cy_225,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_138,
      O => rx_input_memio_bp_4_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_192 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_225,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_138,
      O => rx_input_memio_n0043(5)
    );
  rx_input_memio_bp_4_CYINIT_451 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_224,
      O => rx_input_memio_bp_4_CYINIT
    );
  rx_input_memio_bp_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_6_FFY_RST
    );
  rx_input_memio_bp_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(7),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_6_FFY_RST,
      O => rx_input_memio_bp(7)
    );
  rx_input_memio_Msub_n0043_inst_cy_227_452 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_76,
      IB => rx_input_memio_bp_6_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_139,
      O => rx_input_memio_Msub_n0043_inst_cy_227
    );
  rx_input_memio_Msub_n0043_inst_sum_193 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_6_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_139,
      O => rx_input_memio_n0043(6)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1391 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_76,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_139
    );
  rx_input_memio_Msub_n0043_inst_lut2_1401 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_77,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_140
    );
  rx_input_memio_bp_6_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_6_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_228
    );
  rx_input_memio_Msub_n0043_inst_cy_228_453 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_77,
      IB => rx_input_memio_Msub_n0043_inst_cy_227,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_140,
      O => rx_input_memio_bp_6_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_194 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_227,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_140,
      O => rx_input_memio_n0043(7)
    );
  rx_input_memio_bp_6_CYINIT_454 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_226,
      O => rx_input_memio_bp_6_CYINIT
    );
  rx_input_memio_bp_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_8_FFY_RST
    );
  rx_input_memio_bp_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(9),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_8_FFY_RST,
      O => rx_input_memio_bp(9)
    );
  rx_input_memio_Msub_n0043_inst_cy_229_455 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_78,
      IB => rx_input_memio_bp_8_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_141,
      O => rx_input_memio_Msub_n0043_inst_cy_229
    );
  rx_input_memio_Msub_n0043_inst_sum_195 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_8_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_141,
      O => rx_input_memio_n0043(8)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1411 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_78,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_141
    );
  rx_input_memio_Msub_n0043_inst_lut2_1421 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_79,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_142
    );
  rx_input_memio_bp_8_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_8_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_230
    );
  rx_input_memio_Msub_n0043_inst_cy_230_456 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_79,
      IB => rx_input_memio_Msub_n0043_inst_cy_229,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_142,
      O => rx_input_memio_bp_8_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_196 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_229,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_142,
      O => rx_input_memio_n0043(9)
    );
  rx_input_memio_bp_8_CYINIT_457 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_228,
      O => rx_input_memio_bp_8_CYINIT
    );
  tx_output_FBBP_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(15),
      CE => txfbbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_15_FFX_RST,
      O => txfbbp(15)
    );
  txfbbp_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_15_FFX_RST
    );
  rx_input_memio_bp_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_10_FFY_RST
    );
  rx_input_memio_bp_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(11),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_10_FFY_RST,
      O => rx_input_memio_bp(11)
    );
  rx_input_memio_Msub_n0043_inst_cy_231_458 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_80,
      IB => rx_input_memio_bp_10_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_143,
      O => rx_input_memio_Msub_n0043_inst_cy_231
    );
  rx_input_memio_Msub_n0043_inst_sum_197 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_10_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_143,
      O => rx_input_memio_n0043(10)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1431 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_80,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_143
    );
  rx_input_memio_Msub_n0043_inst_lut2_1441 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_81,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_144
    );
  rx_input_memio_bp_10_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_10_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_232
    );
  rx_input_memio_Msub_n0043_inst_cy_232_459 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_81,
      IB => rx_input_memio_Msub_n0043_inst_cy_231,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_144,
      O => rx_input_memio_bp_10_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_198 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_231,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_144,
      O => rx_input_memio_n0043(11)
    );
  rx_input_memio_bp_10_CYINIT_460 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_230,
      O => rx_input_memio_bp_10_CYINIT
    );
  rx_input_memio_bp_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_12_FFY_RST
    );
  rx_input_memio_bp_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(13),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_12_FFY_RST,
      O => rx_input_memio_bp(13)
    );
  rx_input_memio_Msub_n0043_inst_cy_233_461 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_82,
      IB => rx_input_memio_bp_12_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_145,
      O => rx_input_memio_Msub_n0043_inst_cy_233
    );
  rx_input_memio_Msub_n0043_inst_sum_199 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_12_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_145,
      O => rx_input_memio_n0043(12)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1451 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_82,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_145
    );
  rx_input_memio_Msub_n0043_inst_lut2_1461 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_83,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_146
    );
  rx_input_memio_bp_12_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bp_12_CYMUXG,
      O => rx_input_memio_Msub_n0043_inst_cy_234
    );
  rx_input_memio_Msub_n0043_inst_cy_234_462 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_83,
      IB => rx_input_memio_Msub_n0043_inst_cy_233,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_146,
      O => rx_input_memio_bp_12_CYMUXG
    );
  rx_input_memio_Msub_n0043_inst_sum_200 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_233,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_146,
      O => rx_input_memio_n0043(13)
    );
  rx_input_memio_bp_12_CYINIT_463 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_232,
      O => rx_input_memio_bp_12_CYINIT
    );
  rx_input_memio_bp_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_14_FFY_RST
    );
  rx_input_memio_bp_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(15),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_14_FFY_RST,
      O => rx_input_memio_bp(15)
    );
  rx_input_memio_Msub_n0043_inst_cy_235_464 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_84,
      IB => rx_input_memio_bp_14_CYINIT,
      SEL => rx_input_memio_Msub_n0043_inst_lut2_147,
      O => rx_input_memio_Msub_n0043_inst_cy_235
    );
  rx_input_memio_Msub_n0043_inst_sum_201 : X_XOR2
    port map (
      I0 => rx_input_memio_bp_14_CYINIT,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_147,
      O => rx_input_memio_n0043(14)
    );
  rx_input_memio_Msub_n0043_inst_lut2_1471 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_84,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_147
    );
  rx_input_memio_Msub_n0043_inst_lut2_1481 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_macnt_85,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0043_inst_lut2_148
    );
  rx_input_memio_Msub_n0043_inst_sum_202 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0043_inst_cy_235,
      I1 => rx_input_memio_Msub_n0043_inst_lut2_148,
      O => rx_input_memio_n0043(15)
    );
  rx_input_memio_bp_14_CYINIT_465 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0043_inst_cy_234,
      O => rx_input_memio_bp_14_CYINIT
    );
  mac_control_rxoferr_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(1),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(1)
    );
  mac_control_rxoferr_cnt_0_LOGIC_ZERO_466 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_0_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_16_467 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_16,
      IB => mac_control_rxoferr_cnt_0_LOGIC_ZERO,
      SEL => mac_control_rxoferr_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_16,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(0),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_rxoferr_cnt_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_24,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(1),
      O => mac_control_rxoferr_cnt_0_GROM
    );
  mac_control_rxoferr_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_0_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_17_468 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_24,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_rxoferr_cnt_0_GROM,
      O => mac_control_rxoferr_cnt_0_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_rxoferr_cnt_0_GROM,
      O => mac_control_rxoferr_cnt_n0000(1)
    );
  mac_control_rxoferr_cnt_2_LOGIC_ZERO_469 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_2_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_18_470 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_2_CYINIT,
      SEL => mac_control_rxoferr_cnt_2_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_2_CYINIT,
      I1 => mac_control_rxoferr_cnt_2_FROM,
      O => mac_control_rxoferr_cnt_n0000(2)
    );
  mac_control_rxoferr_cnt_2_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(2),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_2_FROM
    );
  mac_control_rxoferr_cnt_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(3),
      O => mac_control_rxoferr_cnt_2_GROM
    );
  mac_control_rxoferr_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_2_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_19_471 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_rxoferr_cnt_2_GROM,
      O => mac_control_rxoferr_cnt_2_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_rxoferr_cnt_2_GROM,
      O => mac_control_rxoferr_cnt_n0000(3)
    );
  mac_control_rxoferr_cnt_2_CYINIT_472 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_rxoferr_cnt_2_CYINIT
    );
  mac_control_rxoferr_cnt_4_LOGIC_ZERO_473 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_4_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_20_474 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_4_CYINIT,
      SEL => mac_control_rxoferr_cnt_4_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_4_CYINIT,
      I1 => mac_control_rxoferr_cnt_4_FROM,
      O => mac_control_rxoferr_cnt_n0000(4)
    );
  mac_control_rxoferr_cnt_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxoferr_cnt(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_4_FROM
    );
  mac_control_rxoferr_cnt_4_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(5),
      O => mac_control_rxoferr_cnt_4_GROM
    );
  mac_control_rxoferr_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_4_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_21_475 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_rxoferr_cnt_4_GROM,
      O => mac_control_rxoferr_cnt_4_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_rxoferr_cnt_4_GROM,
      O => mac_control_rxoferr_cnt_n0000(5)
    );
  mac_control_rxoferr_cnt_4_CYINIT_476 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_rxoferr_cnt_4_CYINIT
    );
  mac_control_rxoferr_cnt_6_LOGIC_ZERO_477 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_6_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_22_478 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_6_CYINIT,
      SEL => mac_control_rxoferr_cnt_6_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_6_CYINIT,
      I1 => mac_control_rxoferr_cnt_6_FROM,
      O => mac_control_rxoferr_cnt_n0000(6)
    );
  mac_control_rxoferr_cnt_6_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(6),
      O => mac_control_rxoferr_cnt_6_FROM
    );
  mac_control_rxoferr_cnt_6_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(7),
      O => mac_control_rxoferr_cnt_6_GROM
    );
  mac_control_rxoferr_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_6_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_23_479 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_rxoferr_cnt_6_GROM,
      O => mac_control_rxoferr_cnt_6_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_rxoferr_cnt_6_GROM,
      O => mac_control_rxoferr_cnt_n0000(7)
    );
  mac_control_rxoferr_cnt_6_CYINIT_480 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_rxoferr_cnt_6_CYINIT
    );
  mac_control_rxoferr_cnt_8_LOGIC_ZERO_481 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_8_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_24_482 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_8_CYINIT,
      SEL => mac_control_rxoferr_cnt_8_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_8_CYINIT,
      I1 => mac_control_rxoferr_cnt_8_FROM,
      O => mac_control_rxoferr_cnt_n0000(8)
    );
  mac_control_rxoferr_cnt_8_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxoferr_cnt(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_8_FROM
    );
  mac_control_rxoferr_cnt_8_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(9),
      O => mac_control_rxoferr_cnt_8_GROM
    );
  mac_control_rxoferr_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_8_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_25_483 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_rxoferr_cnt_8_GROM,
      O => mac_control_rxoferr_cnt_8_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_rxoferr_cnt_8_GROM,
      O => mac_control_rxoferr_cnt_n0000(9)
    );
  mac_control_rxoferr_cnt_8_CYINIT_484 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_rxoferr_cnt_8_CYINIT
    );
  mac_control_rxoferr_cnt_10_LOGIC_ZERO_485 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_10_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_26_486 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_10_CYINIT,
      SEL => mac_control_rxoferr_cnt_10_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_10_CYINIT,
      I1 => mac_control_rxoferr_cnt_10_FROM,
      O => mac_control_rxoferr_cnt_n0000(10)
    );
  mac_control_rxoferr_cnt_10_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(10),
      O => mac_control_rxoferr_cnt_10_FROM
    );
  mac_control_rxoferr_cnt_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(11),
      O => mac_control_rxoferr_cnt_10_GROM
    );
  mac_control_rxoferr_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_10_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_27_487 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_rxoferr_cnt_10_GROM,
      O => mac_control_rxoferr_cnt_10_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_rxoferr_cnt_10_GROM,
      O => mac_control_rxoferr_cnt_n0000(11)
    );
  mac_control_rxoferr_cnt_10_CYINIT_488 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_rxoferr_cnt_10_CYINIT
    );
  mac_control_rxoferr_cnt_12_LOGIC_ZERO_489 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_12_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_28_490 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_12_CYINIT,
      SEL => mac_control_rxoferr_cnt_12_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_12_CYINIT,
      I1 => mac_control_rxoferr_cnt_12_FROM,
      O => mac_control_rxoferr_cnt_n0000(12)
    );
  mac_control_rxoferr_cnt_12_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(12),
      O => mac_control_rxoferr_cnt_12_FROM
    );
  mac_control_rxoferr_cnt_12_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(13),
      O => mac_control_rxoferr_cnt_12_GROM
    );
  mac_control_rxoferr_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_12_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_29_491 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_rxoferr_cnt_12_GROM,
      O => mac_control_rxoferr_cnt_12_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_rxoferr_cnt_12_GROM,
      O => mac_control_rxoferr_cnt_n0000(13)
    );
  mac_control_rxoferr_cnt_12_CYINIT_492 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_rxoferr_cnt_12_CYINIT
    );
  mac_control_rxoferr_cnt_14_LOGIC_ZERO_493 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_14_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_30_494 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_14_CYINIT,
      SEL => mac_control_rxoferr_cnt_14_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_14_CYINIT,
      I1 => mac_control_rxoferr_cnt_14_FROM,
      O => mac_control_rxoferr_cnt_n0000(14)
    );
  mac_control_rxoferr_cnt_14_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(14),
      O => mac_control_rxoferr_cnt_14_FROM
    );
  mac_control_rxoferr_cnt_14_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(15),
      O => mac_control_rxoferr_cnt_14_GROM
    );
  mac_control_rxoferr_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_14_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_31_495 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_rxoferr_cnt_14_GROM,
      O => mac_control_rxoferr_cnt_14_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_rxoferr_cnt_14_GROM,
      O => mac_control_rxoferr_cnt_n0000(15)
    );
  mac_control_rxoferr_cnt_14_CYINIT_496 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_rxoferr_cnt_14_CYINIT
    );
  rx_input_memio_dout_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_9_FFY_RST,
      O => rx_input_memio_dout(8)
    );
  rx_input_memio_dout_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_9_FFY_RST
    );
  mac_control_rxoferr_cnt_16_LOGIC_ZERO_497 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_16_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_32_498 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_16_CYINIT,
      SEL => mac_control_rxoferr_cnt_16_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_16_CYINIT,
      I1 => mac_control_rxoferr_cnt_16_FROM,
      O => mac_control_rxoferr_cnt_n0000(16)
    );
  mac_control_rxoferr_cnt_16_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(16),
      O => mac_control_rxoferr_cnt_16_FROM
    );
  mac_control_rxoferr_cnt_16_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(17),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_16_GROM
    );
  mac_control_rxoferr_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_16_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_33_499 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_rxoferr_cnt_16_GROM,
      O => mac_control_rxoferr_cnt_16_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_rxoferr_cnt_16_GROM,
      O => mac_control_rxoferr_cnt_n0000(17)
    );
  mac_control_rxoferr_cnt_16_CYINIT_500 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_rxoferr_cnt_16_CYINIT
    );
  addr3ext_7_LOGIC_ZERO_501 : X_ZERO
    port map (
      O => addr3ext_7_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_109_502 : X_MUX2
    port map (
      IA => addr3ext_7_LOGIC_ZERO,
      IB => addr3ext_7_CYINIT,
      SEL => rx_output_macnt_inst_lut3_7,
      O => rx_output_macnt_inst_cy_109
    );
  rx_output_macnt_inst_sum_102_503 : X_XOR2
    port map (
      I0 => addr3ext_7_CYINIT,
      I1 => rx_output_macnt_inst_lut3_7,
      O => rx_output_macnt_inst_sum_102
    );
  rx_output_macnt_inst_lut3_71 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => addr3ext(7),
      ADR1 => rx_output_cs_FFd19,
      ADR2 => rx_output_bp(7),
      ADR3 => VCC,
      O => rx_output_macnt_inst_lut3_7
    );
  rx_output_macnt_inst_lut3_81 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_bp(8),
      ADR2 => addr3ext(8),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_8
    );
  addr3ext_7_COUTUSED : X_BUF
    port map (
      I => addr3ext_7_CYMUXG,
      O => rx_output_macnt_inst_cy_110
    );
  rx_output_macnt_inst_cy_110_504 : X_MUX2
    port map (
      IA => addr3ext_7_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_109,
      SEL => rx_output_macnt_inst_lut3_8,
      O => addr3ext_7_CYMUXG
    );
  rx_output_macnt_inst_sum_103_505 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_109,
      I1 => rx_output_macnt_inst_lut3_8,
      O => rx_output_macnt_inst_sum_103
    );
  addr3ext_7_CYINIT_506 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_108,
      O => addr3ext_7_CYINIT
    );
  addr3ext_9_LOGIC_ZERO_507 : X_ZERO
    port map (
      O => addr3ext_9_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_111_508 : X_MUX2
    port map (
      IA => addr3ext_9_LOGIC_ZERO,
      IB => addr3ext_9_CYINIT,
      SEL => rx_output_macnt_inst_lut3_9,
      O => rx_output_macnt_inst_cy_111
    );
  rx_output_macnt_inst_sum_104_509 : X_XOR2
    port map (
      I0 => addr3ext_9_CYINIT,
      I1 => rx_output_macnt_inst_lut3_9,
      O => rx_output_macnt_inst_sum_104
    );
  rx_output_macnt_inst_lut3_91 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(9),
      ADR2 => rx_output_bp(9),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_9
    );
  rx_output_macnt_inst_lut3_101 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_bp(10),
      ADR2 => addr3ext(10),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_10
    );
  addr3ext_9_COUTUSED : X_BUF
    port map (
      I => addr3ext_9_CYMUXG,
      O => rx_output_macnt_inst_cy_112
    );
  rx_output_macnt_inst_cy_112_510 : X_MUX2
    port map (
      IA => addr3ext_9_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_111,
      SEL => rx_output_macnt_inst_lut3_10,
      O => addr3ext_9_CYMUXG
    );
  rx_output_macnt_inst_sum_105_511 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_111,
      I1 => rx_output_macnt_inst_lut3_10,
      O => rx_output_macnt_inst_sum_105
    );
  addr3ext_9_CYINIT_512 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_110,
      O => addr3ext_9_CYINIT
    );
  rx_input_fifo_control_DATA_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(5),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_5_FFY_RST,
      O => rx_input_data(5)
    );
  rx_input_data_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_5_FFY_RST
    );
  addr3ext_11_LOGIC_ZERO_513 : X_ZERO
    port map (
      O => addr3ext_11_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_113_514 : X_MUX2
    port map (
      IA => addr3ext_11_LOGIC_ZERO,
      IB => addr3ext_11_CYINIT,
      SEL => rx_output_macnt_inst_lut3_11,
      O => rx_output_macnt_inst_cy_113
    );
  rx_output_macnt_inst_sum_106_515 : X_XOR2
    port map (
      I0 => addr3ext_11_CYINIT,
      I1 => rx_output_macnt_inst_lut3_11,
      O => rx_output_macnt_inst_sum_106
    );
  rx_output_macnt_inst_lut3_111 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(11),
      ADR2 => rx_output_bp(11),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_11
    );
  rx_output_macnt_inst_lut3_121 : X_LUT4
    generic map(
      INIT => X"D8D8"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => rx_output_bp(12),
      ADR2 => addr3ext(12),
      ADR3 => VCC,
      O => rx_output_macnt_inst_lut3_12
    );
  addr3ext_11_COUTUSED : X_BUF
    port map (
      I => addr3ext_11_CYMUXG,
      O => rx_output_macnt_inst_cy_114
    );
  rx_output_macnt_inst_cy_114_516 : X_MUX2
    port map (
      IA => addr3ext_11_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_113,
      SEL => rx_output_macnt_inst_lut3_12,
      O => addr3ext_11_CYMUXG
    );
  rx_output_macnt_inst_sum_107_517 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_113,
      I1 => rx_output_macnt_inst_lut3_12,
      O => rx_output_macnt_inst_sum_107
    );
  addr3ext_11_CYINIT_518 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_112,
      O => addr3ext_11_CYINIT
    );
  addr3ext_13_LOGIC_ZERO_519 : X_ZERO
    port map (
      O => addr3ext_13_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_115_520 : X_MUX2
    port map (
      IA => addr3ext_13_LOGIC_ZERO,
      IB => addr3ext_13_CYINIT,
      SEL => rx_output_macnt_inst_lut3_13,
      O => rx_output_macnt_inst_cy_115
    );
  rx_output_macnt_inst_sum_108_521 : X_XOR2
    port map (
      I0 => addr3ext_13_CYINIT,
      I1 => rx_output_macnt_inst_lut3_13,
      O => rx_output_macnt_inst_sum_108
    );
  rx_output_macnt_inst_lut3_131 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(13),
      ADR2 => rx_output_bp(13),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_13
    );
  rx_output_macnt_inst_lut3_141 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => addr3ext(14),
      ADR1 => rx_output_cs_FFd19,
      ADR2 => rx_output_bp(14),
      ADR3 => VCC,
      O => rx_output_macnt_inst_lut3_14
    );
  addr3ext_13_COUTUSED : X_BUF
    port map (
      I => addr3ext_13_CYMUXG,
      O => rx_output_macnt_inst_cy_116
    );
  rx_output_macnt_inst_cy_116_522 : X_MUX2
    port map (
      IA => addr3ext_13_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_115,
      SEL => rx_output_macnt_inst_lut3_14,
      O => addr3ext_13_CYMUXG
    );
  rx_output_macnt_inst_sum_109_523 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_115,
      I1 => rx_output_macnt_inst_lut3_14,
      O => rx_output_macnt_inst_sum_109
    );
  addr3ext_13_CYINIT_524 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_114,
      O => addr3ext_13_CYINIT
    );
  rx_output_macnt_inst_sum_110_525 : X_XOR2
    port map (
      I0 => addr3ext_15_CYINIT,
      I1 => rx_output_macnt_inst_lut3_15,
      O => rx_output_macnt_inst_sum_110
    );
  rx_output_macnt_inst_lut3_151 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(15),
      ADR2 => rx_output_bp(15),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_15
    );
  addr3ext_15_CYINIT_526 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_116,
      O => addr3ext_15_CYINIT
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE_527 : X_ONE
    port map (
      O => rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO_528 : X_ZERO
    port map (
      O => rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_151_529 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE,
      SEL => rx_fifocheck_diff_0_rt,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_151
    );
  rx_fifocheck_diff_0_rt_530 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_fifocheck_diff(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_diff_0_rt
    );
  rx_fifocheck_BEL_2 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_fifocheck_diff(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_SIG_21
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_152_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_152
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_152_531 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_151,
      SEL => rx_fifocheck_SIG_21,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE_532 : X_ONE
    port map (
      O => rx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_153_533 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut4_8,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_153
    );
  rx_fifocheck_Mcompar_n0003_inst_lut4_81 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(2),
      ADR1 => rx_fifocheck_diff(4),
      ADR2 => rx_fifocheck_diff(1),
      ADR3 => rx_fifocheck_diff(3),
      O => rx_fifocheck_Mcompar_n0003_inst_lut4_8
    );
  rx_fifocheck_Mcompar_n0003_inst_lut4_91 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(4),
      ADR1 => rx_fifocheck_diff(1),
      ADR2 => rx_fifocheck_diff(3),
      ADR3 => rx_fifocheck_diff(2),
      O => rx_fifocheck_Mcompar_n0003_inst_lut4_9
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_154_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_154
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_154_534 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_153,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut4_9,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT_535 : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_152,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT
    );
  tx_output_cs_FFd4_536 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd4_FFX_RST,
      O => tx_output_cs_FFd4
    );
  tx_output_cs_FFd4_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd4_FFX_RST
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE_537 : X_ONE
    port map (
      O => rx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_155_538 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut4_10,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_155
    );
  rx_fifocheck_Mcompar_n0003_inst_lut4_101 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(6),
      ADR1 => rx_fifocheck_diff(5),
      ADR2 => rx_fifocheck_diff(8),
      ADR3 => rx_fifocheck_diff(7),
      O => rx_fifocheck_Mcompar_n0003_inst_lut4_10
    );
  rx_fifocheck_Mcompar_n0003_inst_lut4_111 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => rx_fifocheck_diff(9),
      ADR1 => rx_fifocheck_diff(11),
      ADR2 => rx_fifocheck_diff(10),
      ADR3 => rx_fifocheck_diff(12),
      O => rx_fifocheck_Mcompar_n0003_inst_lut4_11
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_156_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_156
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_156_539 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_155,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut4_11,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT_540 : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_154,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO_541 : X_ZERO
    port map (
      O => rx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_157_542 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT,
      SEL => rx_fifocheck_diff_13_rt,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_157
    );
  rx_fifocheck_diff_13_rt_543 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_diff(13),
      O => rx_fifocheck_diff_13_rt
    );
  rx_fifocheck_BEL_3 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_fifocheck_diff(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_SIG_22
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_158_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_158
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_158_544 : X_MUX2
    port map (
      IA => rx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_157,
      SEL => rx_fifocheck_SIG_22,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT_545 : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_156,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT
    );
  rx_fifocheck_n0003_LOGIC_ONE_546 : X_ONE
    port map (
      O => rx_fifocheck_n0003_LOGIC_ONE
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_159_547 : X_MUX2
    port map (
      IA => rx_fifocheck_n0003_LOGIC_ONE,
      IB => rx_fifocheck_n0003_CYINIT,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut3_32,
      O => rx_fifocheck_Mcompar_n0003_inst_cy_159
    );
  rx_fifocheck_Mcompar_n0003_inst_lut3_321 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_fifocheck_diff(14),
      ADR2 => VCC,
      ADR3 => rx_fifocheck_diff(15),
      O => rx_fifocheck_Mcompar_n0003_inst_lut3_32
    );
  rx_fifocheck_Mcompar_n0003_inst_lut3_331 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_fifocheck_diff(15),
      ADR2 => VCC,
      ADR3 => rx_fifocheck_diff(14),
      O => rx_fifocheck_Mcompar_n0003_inst_lut3_33
    );
  rx_fifocheck_n0003_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_n0003_CYMUXG,
      O => rx_fifocheck_n0003
    );
  rx_fifocheck_Mcompar_n0003_inst_cy_160 : X_MUX2
    port map (
      IA => rx_fifocheck_n0003_LOGIC_ONE,
      IB => rx_fifocheck_Mcompar_n0003_inst_cy_159,
      SEL => rx_fifocheck_Mcompar_n0003_inst_lut3_33,
      O => rx_fifocheck_n0003_CYMUXG
    );
  rx_fifocheck_n0003_CYINIT_548 : X_BUF
    port map (
      I => rx_fifocheck_Mcompar_n0003_inst_cy_158,
      O => rx_fifocheck_n0003_CYINIT
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE_549 : X_ONE
    port map (
      O => tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO_550 : X_ZERO
    port map (
      O => tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_151_551 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ONE,
      SEL => tx_fifocheck_diff_0_rt,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_151
    );
  tx_fifocheck_diff_0_rt_552 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_fifocheck_diff(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_diff_0_rt
    );
  tx_fifocheck_BEL_4 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => tx_fifocheck_diff(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_SIG_23
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_152_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_152
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_152_553 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_152_LOGIC_ZERO,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_151,
      SEL => tx_fifocheck_SIG_23,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_152_CYMUXG
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE_554 : X_ONE
    port map (
      O => tx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_153_555 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut4_8,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_153
    );
  tx_fifocheck_Mcompar_n0003_inst_lut4_81 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(4),
      ADR1 => tx_fifocheck_diff(2),
      ADR2 => tx_fifocheck_diff(3),
      ADR3 => tx_fifocheck_diff(1),
      O => tx_fifocheck_Mcompar_n0003_inst_lut4_8
    );
  tx_fifocheck_Mcompar_n0003_inst_lut4_91 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(3),
      ADR1 => tx_fifocheck_diff(2),
      ADR2 => tx_fifocheck_diff(1),
      ADR3 => tx_fifocheck_diff(4),
      O => tx_fifocheck_Mcompar_n0003_inst_lut4_9
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_154_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_154
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_154_556 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_154_LOGIC_ONE,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_153,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut4_9,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_154_CYMUXG
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT_557 : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_152,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_154_CYINIT
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE_558 : X_ONE
    port map (
      O => tx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_155_559 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut4_10,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_155
    );
  tx_fifocheck_Mcompar_n0003_inst_lut4_101 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(8),
      ADR1 => tx_fifocheck_diff(5),
      ADR2 => tx_fifocheck_diff(7),
      ADR3 => tx_fifocheck_diff(6),
      O => tx_fifocheck_Mcompar_n0003_inst_lut4_10
    );
  tx_fifocheck_Mcompar_n0003_inst_lut4_111 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(11),
      ADR1 => tx_fifocheck_diff(9),
      ADR2 => tx_fifocheck_diff(10),
      ADR3 => tx_fifocheck_diff(12),
      O => tx_fifocheck_Mcompar_n0003_inst_lut4_11
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_156_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_156
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_156_560 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_156_LOGIC_ONE,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_155,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut4_11,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_156_CYMUXG
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT_561 : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_154,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_156_CYINIT
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO_562 : X_ZERO
    port map (
      O => tx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_157_563 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT,
      SEL => tx_fifocheck_diff_13_rt,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_157
    );
  tx_fifocheck_diff_13_rt_564 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_fifocheck_diff(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_diff_13_rt
    );
  tx_fifocheck_BEL_5 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_fifocheck_diff(13),
      ADR3 => VCC,
      O => tx_fifocheck_SIG_24
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_158_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_158
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_158_565 : X_MUX2
    port map (
      IA => tx_fifocheck_Mcompar_n0003_inst_cy_158_LOGIC_ZERO,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_157,
      SEL => tx_fifocheck_SIG_24,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_158_CYMUXG
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT_566 : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_156,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_158_CYINIT
    );
  tx_fifocheck_n0003_LOGIC_ONE_567 : X_ONE
    port map (
      O => tx_fifocheck_n0003_LOGIC_ONE
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_159_568 : X_MUX2
    port map (
      IA => tx_fifocheck_n0003_LOGIC_ONE,
      IB => tx_fifocheck_n0003_CYINIT,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut3_32,
      O => tx_fifocheck_Mcompar_n0003_inst_cy_159
    );
  tx_fifocheck_Mcompar_n0003_inst_lut3_321 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_fifocheck_diff(15),
      ADR2 => VCC,
      ADR3 => tx_fifocheck_diff(14),
      O => tx_fifocheck_Mcompar_n0003_inst_lut3_32
    );
  tx_fifocheck_Mcompar_n0003_inst_lut3_331 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_fifocheck_diff(15),
      ADR3 => tx_fifocheck_diff(14),
      O => tx_fifocheck_Mcompar_n0003_inst_lut3_33
    );
  tx_fifocheck_n0003_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_n0003_CYMUXG,
      O => tx_fifocheck_n0003
    );
  tx_fifocheck_Mcompar_n0003_inst_cy_160 : X_MUX2
    port map (
      IA => tx_fifocheck_n0003_LOGIC_ONE,
      IB => tx_fifocheck_Mcompar_n0003_inst_cy_159,
      SEL => tx_fifocheck_Mcompar_n0003_inst_lut3_33,
      O => tx_fifocheck_n0003_CYMUXG
    );
  tx_fifocheck_n0003_CYINIT_569 : X_BUF
    port map (
      I => tx_fifocheck_Mcompar_n0003_inst_cy_158,
      O => tx_fifocheck_n0003_CYINIT
    );
  mac_control_phyrstcnt_110_LOGIC_ONE_570 : X_ONE
    port map (
      O => mac_control_phyrstcnt_110_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_294_571 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_16,
      IB => mac_control_phyrstcnt_110_LOGIC_ONE,
      SEL => mac_control_N53144_rt,
      O => mac_control_phyrstcnt_inst_cy_294
    );
  mac_control_N53144_rt_572 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_16,
      ADR1 => VCC,
      ADR2 => mac_control_N53144,
      ADR3 => VCC,
      O => mac_control_N53144_rt
    );
  mac_control_phyrstcnt_inst_lut3_1921 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_9,
      ADR1 => VCC,
      ADR2 => mac_control_N53144,
      ADR3 => mac_control_phyrstcnt_110,
      O => mac_control_phyrstcnt_inst_lut3_192
    );
  mac_control_phyrstcnt_110_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_110_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_295
    );
  mac_control_phyrstcnt_inst_cy_295_573 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_9,
      IB => mac_control_phyrstcnt_inst_cy_294,
      SEL => mac_control_phyrstcnt_inst_lut3_192,
      O => mac_control_phyrstcnt_110_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_257_574 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_294,
      I1 => mac_control_phyrstcnt_inst_lut3_192,
      O => mac_control_phyrstcnt_inst_sum_257
    );
  mac_control_phyrstcnt_111_LOGIC_ONE_575 : X_ONE
    port map (
      O => mac_control_phyrstcnt_111_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_296_576 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_111_LOGIC_ONE,
      IB => mac_control_phyrstcnt_111_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_193,
      O => mac_control_phyrstcnt_inst_cy_296
    );
  mac_control_phyrstcnt_inst_sum_258_577 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_111_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_193,
      O => mac_control_phyrstcnt_inst_sum_258
    );
  mac_control_phyrstcnt_inst_lut3_1931 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_111,
      ADR1 => mac_control_N53144,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_193
    );
  mac_control_phyrstcnt_inst_lut3_1941 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N53144,
      ADR2 => mac_control_phyrstcnt_112,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_194
    );
  mac_control_phyrstcnt_111_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_111_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_297
    );
  mac_control_phyrstcnt_inst_cy_297_578 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_111_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_296,
      SEL => mac_control_phyrstcnt_inst_lut3_194,
      O => mac_control_phyrstcnt_111_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_259_579 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_296,
      I1 => mac_control_phyrstcnt_inst_lut3_194,
      O => mac_control_phyrstcnt_inst_sum_259
    );
  mac_control_phyrstcnt_111_CYINIT_580 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_295,
      O => mac_control_phyrstcnt_111_CYINIT
    );
  mac_control_phyrstcnt_113_LOGIC_ONE_581 : X_ONE
    port map (
      O => mac_control_phyrstcnt_113_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_298_582 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_113_LOGIC_ONE,
      IB => mac_control_phyrstcnt_113_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_195,
      O => mac_control_phyrstcnt_inst_cy_298
    );
  mac_control_phyrstcnt_inst_sum_260_583 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_113_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_195,
      O => mac_control_phyrstcnt_inst_sum_260
    );
  mac_control_phyrstcnt_inst_lut3_1951 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => mac_control_phyrstcnt_113,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_195
    );
  mac_control_phyrstcnt_inst_lut3_1961 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_114,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_196
    );
  mac_control_phyrstcnt_113_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_113_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_299
    );
  mac_control_phyrstcnt_inst_cy_299_584 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_113_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_298,
      SEL => mac_control_phyrstcnt_inst_lut3_196,
      O => mac_control_phyrstcnt_113_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_261_585 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_298,
      I1 => mac_control_phyrstcnt_inst_lut3_196,
      O => mac_control_phyrstcnt_inst_sum_261
    );
  mac_control_phyrstcnt_113_CYINIT_586 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_297,
      O => mac_control_phyrstcnt_113_CYINIT
    );
  mac_control_phyrstcnt_115_LOGIC_ONE_587 : X_ONE
    port map (
      O => mac_control_phyrstcnt_115_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_300_588 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_115_LOGIC_ONE,
      IB => mac_control_phyrstcnt_115_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_197,
      O => mac_control_phyrstcnt_inst_cy_300
    );
  mac_control_phyrstcnt_inst_sum_262_589 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_115_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_197,
      O => mac_control_phyrstcnt_inst_sum_262
    );
  mac_control_phyrstcnt_inst_lut3_1971 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_115,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_N53144,
      O => mac_control_phyrstcnt_inst_lut3_197
    );
  mac_control_phyrstcnt_inst_lut3_1981 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_116,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_198
    );
  mac_control_phyrstcnt_115_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_115_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_301
    );
  mac_control_phyrstcnt_inst_cy_301_590 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_115_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_300,
      SEL => mac_control_phyrstcnt_inst_lut3_198,
      O => mac_control_phyrstcnt_115_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_263_591 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_300,
      I1 => mac_control_phyrstcnt_inst_lut3_198,
      O => mac_control_phyrstcnt_inst_sum_263
    );
  mac_control_phyrstcnt_115_CYINIT_592 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_299,
      O => mac_control_phyrstcnt_115_CYINIT
    );
  mac_control_phyrstcnt_117_LOGIC_ONE_593 : X_ONE
    port map (
      O => mac_control_phyrstcnt_117_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_302_594 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_117_LOGIC_ONE,
      IB => mac_control_phyrstcnt_117_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_199,
      O => mac_control_phyrstcnt_inst_cy_302
    );
  mac_control_phyrstcnt_inst_sum_264_595 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_117_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_199,
      O => mac_control_phyrstcnt_inst_sum_264
    );
  mac_control_phyrstcnt_inst_lut3_1991 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_117,
      O => mac_control_phyrstcnt_inst_lut3_199
    );
  mac_control_phyrstcnt_inst_lut3_2001 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_118,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_200
    );
  mac_control_phyrstcnt_117_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_117_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_303
    );
  mac_control_phyrstcnt_inst_cy_303_596 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_117_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_302,
      SEL => mac_control_phyrstcnt_inst_lut3_200,
      O => mac_control_phyrstcnt_117_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_265_597 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_302,
      I1 => mac_control_phyrstcnt_inst_lut3_200,
      O => mac_control_phyrstcnt_inst_sum_265
    );
  mac_control_phyrstcnt_117_CYINIT_598 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_301,
      O => mac_control_phyrstcnt_117_CYINIT
    );
  mac_control_phyrstcnt_119_LOGIC_ONE_599 : X_ONE
    port map (
      O => mac_control_phyrstcnt_119_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_304_600 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_119_LOGIC_ONE,
      IB => mac_control_phyrstcnt_119_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_201,
      O => mac_control_phyrstcnt_inst_cy_304
    );
  mac_control_phyrstcnt_inst_sum_266_601 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_119_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_201,
      O => mac_control_phyrstcnt_inst_sum_266
    );
  mac_control_phyrstcnt_inst_lut3_2011 : X_LUT4
    generic map(
      INIT => X"BBBB"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => mac_control_phyrstcnt_119,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_201
    );
  mac_control_phyrstcnt_inst_lut3_2021 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_120,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_202
    );
  mac_control_phyrstcnt_119_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_119_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_305
    );
  mac_control_phyrstcnt_inst_cy_305_602 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_119_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_304,
      SEL => mac_control_phyrstcnt_inst_lut3_202,
      O => mac_control_phyrstcnt_119_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_267_603 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_304,
      I1 => mac_control_phyrstcnt_inst_lut3_202,
      O => mac_control_phyrstcnt_inst_sum_267
    );
  mac_control_phyrstcnt_119_CYINIT_604 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_303,
      O => mac_control_phyrstcnt_119_CYINIT
    );
  mac_control_phyrstcnt_121_LOGIC_ONE_605 : X_ONE
    port map (
      O => mac_control_phyrstcnt_121_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_306_606 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_121_LOGIC_ONE,
      IB => mac_control_phyrstcnt_121_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_203,
      O => mac_control_phyrstcnt_inst_cy_306
    );
  mac_control_phyrstcnt_inst_sum_268_607 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_121_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_203,
      O => mac_control_phyrstcnt_inst_sum_268
    );
  mac_control_phyrstcnt_inst_lut3_2031 : X_LUT4
    generic map(
      INIT => X"FF33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyrstcnt_121,
      ADR2 => VCC,
      ADR3 => mac_control_N53144,
      O => mac_control_phyrstcnt_inst_lut3_203
    );
  mac_control_phyrstcnt_inst_lut3_2041 : X_LUT4
    generic map(
      INIT => X"FF0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_122,
      ADR3 => mac_control_N53144,
      O => mac_control_phyrstcnt_inst_lut3_204
    );
  mac_control_phyrstcnt_121_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_121_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_307
    );
  mac_control_phyrstcnt_inst_cy_307_608 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_121_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_306,
      SEL => mac_control_phyrstcnt_inst_lut3_204,
      O => mac_control_phyrstcnt_121_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_269_609 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_306,
      I1 => mac_control_phyrstcnt_inst_lut3_204,
      O => mac_control_phyrstcnt_inst_sum_269
    );
  mac_control_phyrstcnt_121_CYINIT_610 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_305,
      O => mac_control_phyrstcnt_121_CYINIT
    );
  mac_control_phyrstcnt_123_LOGIC_ONE_611 : X_ONE
    port map (
      O => mac_control_phyrstcnt_123_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_308_612 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_123_LOGIC_ONE,
      IB => mac_control_phyrstcnt_123_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_205,
      O => mac_control_phyrstcnt_inst_cy_308
    );
  mac_control_phyrstcnt_inst_sum_270_613 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_123_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_205,
      O => mac_control_phyrstcnt_inst_sum_270
    );
  mac_control_phyrstcnt_inst_lut3_2051 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_123,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_205
    );
  mac_control_phyrstcnt_inst_lut3_2061 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_124,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_206
    );
  mac_control_phyrstcnt_123_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_123_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_309
    );
  mac_control_phyrstcnt_inst_cy_309_614 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_123_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_308,
      SEL => mac_control_phyrstcnt_inst_lut3_206,
      O => mac_control_phyrstcnt_123_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_271_615 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_308,
      I1 => mac_control_phyrstcnt_inst_lut3_206,
      O => mac_control_phyrstcnt_inst_sum_271
    );
  mac_control_phyrstcnt_123_CYINIT_616 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_307,
      O => mac_control_phyrstcnt_123_CYINIT
    );
  mac_control_phyrstcnt_125_LOGIC_ONE_617 : X_ONE
    port map (
      O => mac_control_phyrstcnt_125_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_310_618 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_125_LOGIC_ONE,
      IB => mac_control_phyrstcnt_125_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_207,
      O => mac_control_phyrstcnt_inst_cy_310
    );
  mac_control_phyrstcnt_inst_sum_272_619 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_125_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_207,
      O => mac_control_phyrstcnt_inst_sum_272
    );
  mac_control_phyrstcnt_inst_lut3_2071 : X_LUT4
    generic map(
      INIT => X"F3F3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyrstcnt_125,
      ADR2 => mac_control_N53144,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_207
    );
  mac_control_phyrstcnt_inst_lut3_2081 : X_LUT4
    generic map(
      INIT => X"F3F3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyrstcnt_126,
      ADR2 => mac_control_N53144,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_208
    );
  mac_control_phyrstcnt_125_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_125_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_311
    );
  mac_control_phyrstcnt_inst_cy_311_620 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_125_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_310,
      SEL => mac_control_phyrstcnt_inst_lut3_208,
      O => mac_control_phyrstcnt_125_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_273_621 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_310,
      I1 => mac_control_phyrstcnt_inst_lut3_208,
      O => mac_control_phyrstcnt_inst_sum_273
    );
  mac_control_phyrstcnt_125_CYINIT_622 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_309,
      O => mac_control_phyrstcnt_125_CYINIT
    );
  mac_control_phyrstcnt_127_LOGIC_ONE_623 : X_ONE
    port map (
      O => mac_control_phyrstcnt_127_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_312_624 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_127_LOGIC_ONE,
      IB => mac_control_phyrstcnt_127_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_209,
      O => mac_control_phyrstcnt_inst_cy_312
    );
  mac_control_phyrstcnt_inst_sum_274_625 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_127_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_209,
      O => mac_control_phyrstcnt_inst_sum_274
    );
  mac_control_phyrstcnt_inst_lut3_2091 : X_LUT4
    generic map(
      INIT => X"F5F5"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_127,
      ADR1 => VCC,
      ADR2 => mac_control_N53144,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_209
    );
  mac_control_phyrstcnt_inst_lut3_2101 : X_LUT4
    generic map(
      INIT => X"F3F3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyrstcnt_128,
      ADR2 => mac_control_N53144,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_210
    );
  mac_control_phyrstcnt_127_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_127_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_313
    );
  mac_control_phyrstcnt_inst_cy_313_626 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_127_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_312,
      SEL => mac_control_phyrstcnt_inst_lut3_210,
      O => mac_control_phyrstcnt_127_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_275_627 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_312,
      I1 => mac_control_phyrstcnt_inst_lut3_210,
      O => mac_control_phyrstcnt_inst_sum_275
    );
  mac_control_phyrstcnt_127_CYINIT_628 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_311,
      O => mac_control_phyrstcnt_127_CYINIT
    );
  mac_control_phyrstcnt_129_LOGIC_ONE_629 : X_ONE
    port map (
      O => mac_control_phyrstcnt_129_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_314_630 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_129_LOGIC_ONE,
      IB => mac_control_phyrstcnt_129_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_211,
      O => mac_control_phyrstcnt_inst_cy_314
    );
  mac_control_phyrstcnt_inst_sum_276_631 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_129_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_211,
      O => mac_control_phyrstcnt_inst_sum_276
    );
  mac_control_phyrstcnt_inst_lut3_2111 : X_LUT4
    generic map(
      INIT => X"F5F5"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_129,
      ADR1 => VCC,
      ADR2 => mac_control_N53144,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_211
    );
  mac_control_phyrstcnt_inst_lut3_2121 : X_LUT4
    generic map(
      INIT => X"AAFF"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_phyrstcnt_130,
      O => mac_control_phyrstcnt_inst_lut3_212
    );
  mac_control_phyrstcnt_129_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_129_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_315
    );
  mac_control_phyrstcnt_inst_cy_315_632 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_129_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_314,
      SEL => mac_control_phyrstcnt_inst_lut3_212,
      O => mac_control_phyrstcnt_129_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_277_633 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_314,
      I1 => mac_control_phyrstcnt_inst_lut3_212,
      O => mac_control_phyrstcnt_inst_sum_277
    );
  mac_control_phyrstcnt_129_CYINIT_634 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_313,
      O => mac_control_phyrstcnt_129_CYINIT
    );
  mac_control_phyrstcnt_131_LOGIC_ONE_635 : X_ONE
    port map (
      O => mac_control_phyrstcnt_131_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_316_636 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_131_LOGIC_ONE,
      IB => mac_control_phyrstcnt_131_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_213,
      O => mac_control_phyrstcnt_inst_cy_316
    );
  mac_control_phyrstcnt_inst_sum_278_637 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_131_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_213,
      O => mac_control_phyrstcnt_inst_sum_278
    );
  mac_control_phyrstcnt_inst_lut3_2131 : X_LUT4
    generic map(
      INIT => X"BBBB"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => mac_control_phyrstcnt_131,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_213
    );
  mac_control_phyrstcnt_inst_lut3_2141 : X_LUT4
    generic map(
      INIT => X"AFAF"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_132,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_214
    );
  mac_control_phyrstcnt_131_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_131_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_317
    );
  mac_control_phyrstcnt_inst_cy_317_638 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_131_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_316,
      SEL => mac_control_phyrstcnt_inst_lut3_214,
      O => mac_control_phyrstcnt_131_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_279_639 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_316,
      I1 => mac_control_phyrstcnt_inst_lut3_214,
      O => mac_control_phyrstcnt_inst_sum_279
    );
  mac_control_phyrstcnt_131_CYINIT_640 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_315,
      O => mac_control_phyrstcnt_131_CYINIT
    );
  mac_control_phyrstcnt_133_LOGIC_ONE_641 : X_ONE
    port map (
      O => mac_control_phyrstcnt_133_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_318_642 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_133_LOGIC_ONE,
      IB => mac_control_phyrstcnt_133_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_215,
      O => mac_control_phyrstcnt_inst_cy_318
    );
  mac_control_phyrstcnt_inst_sum_280_643 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_133_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_215,
      O => mac_control_phyrstcnt_inst_sum_280
    );
  mac_control_phyrstcnt_inst_lut3_2151 : X_LUT4
    generic map(
      INIT => X"FF33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyrstcnt_133,
      ADR2 => VCC,
      ADR3 => mac_control_N53144,
      O => mac_control_phyrstcnt_inst_lut3_215
    );
  mac_control_phyrstcnt_inst_lut3_2161 : X_LUT4
    generic map(
      INIT => X"FF0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_phyrstcnt_134,
      ADR3 => mac_control_N53144,
      O => mac_control_phyrstcnt_inst_lut3_216
    );
  mac_control_phyrstcnt_133_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_133_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_319
    );
  mac_control_phyrstcnt_inst_cy_319_644 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_133_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_318,
      SEL => mac_control_phyrstcnt_inst_lut3_216,
      O => mac_control_phyrstcnt_133_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_281_645 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_318,
      I1 => mac_control_phyrstcnt_inst_lut3_216,
      O => mac_control_phyrstcnt_inst_sum_281
    );
  mac_control_phyrstcnt_133_CYINIT_646 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_317,
      O => mac_control_phyrstcnt_133_CYINIT
    );
  mac_control_phyrstcnt_135_LOGIC_ONE_647 : X_ONE
    port map (
      O => mac_control_phyrstcnt_135_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_320_648 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_135_LOGIC_ONE,
      IB => mac_control_phyrstcnt_135_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_217,
      O => mac_control_phyrstcnt_inst_cy_320
    );
  mac_control_phyrstcnt_inst_sum_282_649 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_135_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_217,
      O => mac_control_phyrstcnt_inst_sum_282
    );
  mac_control_phyrstcnt_inst_lut3_2171 : X_LUT4
    generic map(
      INIT => X"BBBB"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => mac_control_phyrstcnt_135,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_217
    );
  mac_control_phyrstcnt_inst_lut3_2181 : X_LUT4
    generic map(
      INIT => X"BBBB"
    )
    port map (
      ADR0 => mac_control_N53144,
      ADR1 => mac_control_phyrstcnt_136,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_218
    );
  mac_control_phyrstcnt_135_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_135_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_321
    );
  mac_control_phyrstcnt_inst_cy_321_650 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_135_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_320,
      SEL => mac_control_phyrstcnt_inst_lut3_218,
      O => mac_control_phyrstcnt_135_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_283_651 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_320,
      I1 => mac_control_phyrstcnt_inst_lut3_218,
      O => mac_control_phyrstcnt_inst_sum_283
    );
  mac_control_phyrstcnt_135_CYINIT_652 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_319,
      O => mac_control_phyrstcnt_135_CYINIT
    );
  mac_control_phyrstcnt_137_LOGIC_ONE_653 : X_ONE
    port map (
      O => mac_control_phyrstcnt_137_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_322_654 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_137_LOGIC_ONE,
      IB => mac_control_phyrstcnt_137_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_219,
      O => mac_control_phyrstcnt_inst_cy_322
    );
  mac_control_phyrstcnt_inst_sum_284_655 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_137_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_219,
      O => mac_control_phyrstcnt_inst_sum_284
    );
  mac_control_phyrstcnt_inst_lut3_2191 : X_LUT4
    generic map(
      INIT => X"F3F3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyrstcnt_137,
      ADR2 => mac_control_N53144,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_219
    );
  mac_control_phyrstcnt_inst_lut3_2201 : X_LUT4
    generic map(
      INIT => X"F0FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_N53144,
      ADR3 => mac_control_phyrstcnt_138,
      O => mac_control_phyrstcnt_inst_lut3_220
    );
  mac_control_phyrstcnt_137_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_137_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_323
    );
  mac_control_phyrstcnt_inst_cy_323_656 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_137_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_322,
      SEL => mac_control_phyrstcnt_inst_lut3_220,
      O => mac_control_phyrstcnt_137_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_285_657 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_322,
      I1 => mac_control_phyrstcnt_inst_lut3_220,
      O => mac_control_phyrstcnt_inst_sum_285
    );
  mac_control_phyrstcnt_137_CYINIT_658 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_321,
      O => mac_control_phyrstcnt_137_CYINIT
    );
  mac_control_phyrstcnt_139_LOGIC_ONE_659 : X_ONE
    port map (
      O => mac_control_phyrstcnt_139_LOGIC_ONE
    );
  mac_control_phyrstcnt_inst_cy_324_660 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_139_LOGIC_ONE,
      IB => mac_control_phyrstcnt_139_CYINIT,
      SEL => mac_control_phyrstcnt_inst_lut3_221,
      O => mac_control_phyrstcnt_inst_cy_324
    );
  mac_control_phyrstcnt_inst_sum_286_661 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_139_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_221,
      O => mac_control_phyrstcnt_inst_sum_286
    );
  mac_control_phyrstcnt_inst_lut3_2211 : X_LUT4
    generic map(
      INIT => X"F5F5"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_139,
      ADR1 => VCC,
      ADR2 => mac_control_N53144,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_221
    );
  mac_control_phyrstcnt_inst_lut3_2221 : X_LUT4
    generic map(
      INIT => X"F3F3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyrstcnt_140,
      ADR2 => mac_control_N53144,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_222
    );
  mac_control_phyrstcnt_139_COUTUSED : X_BUF
    port map (
      I => mac_control_phyrstcnt_139_CYMUXG,
      O => mac_control_phyrstcnt_inst_cy_325
    );
  mac_control_phyrstcnt_inst_cy_325_662 : X_MUX2
    port map (
      IA => mac_control_phyrstcnt_139_LOGIC_ONE,
      IB => mac_control_phyrstcnt_inst_cy_324,
      SEL => mac_control_phyrstcnt_inst_lut3_222,
      O => mac_control_phyrstcnt_139_CYMUXG
    );
  mac_control_phyrstcnt_inst_sum_287_663 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_inst_cy_324,
      I1 => mac_control_phyrstcnt_inst_lut3_222,
      O => mac_control_phyrstcnt_inst_sum_287
    );
  mac_control_phyrstcnt_139_CYINIT_664 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_323,
      O => mac_control_phyrstcnt_139_CYINIT
    );
  rx_input_fifo_control_DATA_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(6),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_6_FFY_RST,
      O => rx_input_data(6)
    );
  rx_input_data_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_6_FFY_RST
    );
  mac_control_phyrstcnt_inst_sum_288_665 : X_XOR2
    port map (
      I0 => mac_control_phyrstcnt_141_CYINIT,
      I1 => mac_control_phyrstcnt_inst_lut3_223,
      O => mac_control_phyrstcnt_inst_sum_288
    );
  mac_control_phyrstcnt_inst_lut3_2231 : X_LUT4
    generic map(
      INIT => X"F3F3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phyrstcnt_141,
      ADR2 => mac_control_N53144,
      ADR3 => VCC,
      O => mac_control_phyrstcnt_inst_lut3_223
    );
  mac_control_phyrstcnt_141_CYINIT_666 : X_BUF
    port map (
      I => mac_control_phyrstcnt_inst_cy_325,
      O => mac_control_phyrstcnt_141_CYINIT
    );
  rx_input_memio_macnt_70_LOGIC_ZERO_667 : X_ZERO
    port map (
      O => rx_input_memio_macnt_70_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_253_668 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_2,
      IB => rx_input_memio_macnt_70_LOGIC_ZERO,
      SEL => rx_input_memio_cs_FFd16_1_rt,
      O => rx_input_memio_macnt_inst_cy_253
    );
  rx_input_memio_cs_FFd16_1_rt_669 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_2,
      ADR1 => VCC,
      ADR2 => rx_input_memio_cs_FFd16_1,
      ADR3 => VCC,
      O => rx_input_memio_cs_FFd16_1_rt
    );
  rx_input_memio_macnt_inst_lut3_561 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_11,
      ADR1 => rx_input_memio_bp(0),
      ADR2 => rx_input_memio_macnt_70,
      ADR3 => rx_input_memio_cs_FFd16_1,
      O => rx_input_memio_macnt_inst_lut3_56
    );
  rx_input_memio_macnt_70_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_70_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_254
    );
  rx_input_memio_macnt_inst_cy_254_670 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_11,
      IB => rx_input_memio_macnt_inst_cy_253,
      SEL => rx_input_memio_macnt_inst_lut3_56,
      O => rx_input_memio_macnt_70_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_219_671 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_253,
      I1 => rx_input_memio_macnt_inst_lut3_56,
      O => rx_input_memio_macnt_inst_sum_219
    );
  rx_input_memio_macnt_71_LOGIC_ZERO_672 : X_ZERO
    port map (
      O => rx_input_memio_macnt_71_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_255_673 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_71_LOGIC_ZERO,
      IB => rx_input_memio_macnt_71_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_57,
      O => rx_input_memio_macnt_inst_cy_255
    );
  rx_input_memio_macnt_inst_sum_220_674 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_71_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_57,
      O => rx_input_memio_macnt_inst_sum_220
    );
  rx_input_memio_macnt_inst_lut3_571 : X_LUT4
    generic map(
      INIT => X"F3C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd16_2,
      ADR2 => rx_input_memio_bp(1),
      ADR3 => rx_input_memio_macnt_71,
      O => rx_input_memio_macnt_inst_lut3_57
    );
  rx_input_memio_macnt_inst_lut3_581 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16_2,
      ADR1 => rx_input_memio_bp(2),
      ADR2 => VCC,
      ADR3 => rx_input_memio_macnt_72,
      O => rx_input_memio_macnt_inst_lut3_58
    );
  rx_input_memio_macnt_71_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_71_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_256
    );
  rx_input_memio_macnt_71_YUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_71_XORG,
      O => rx_input_memio_macnt_inst_sum_221
    );
  rx_input_memio_macnt_inst_cy_256_675 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_71_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_255,
      SEL => rx_input_memio_macnt_inst_lut3_58,
      O => rx_input_memio_macnt_71_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_221_676 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_255,
      I1 => rx_input_memio_macnt_inst_lut3_58,
      O => rx_input_memio_macnt_71_XORG
    );
  rx_input_memio_macnt_71_CYINIT_677 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_254,
      O => rx_input_memio_macnt_71_CYINIT
    );
  rx_input_memio_macnt_73_LOGIC_ZERO_678 : X_ZERO
    port map (
      O => rx_input_memio_macnt_73_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_257_679 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_73_LOGIC_ZERO,
      IB => rx_input_memio_macnt_73_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_59,
      O => rx_input_memio_macnt_inst_cy_257
    );
  rx_input_memio_macnt_inst_sum_222_680 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_73_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_59,
      O => rx_input_memio_macnt_inst_sum_222
    );
  rx_input_memio_macnt_inst_lut3_591 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => rx_input_memio_macnt_73,
      ADR1 => rx_input_memio_cs_FFd16_2,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bp(3),
      O => rx_input_memio_macnt_inst_lut3_59
    );
  rx_input_memio_macnt_inst_lut3_601 : X_LUT4
    generic map(
      INIT => X"D8D8"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16_2,
      ADR1 => rx_input_memio_bp(4),
      ADR2 => rx_input_memio_macnt_74,
      ADR3 => VCC,
      O => rx_input_memio_macnt_inst_lut3_60
    );
  rx_input_memio_macnt_73_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_73_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_258
    );
  rx_input_memio_macnt_inst_cy_258_681 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_73_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_257,
      SEL => rx_input_memio_macnt_inst_lut3_60,
      O => rx_input_memio_macnt_73_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_223_682 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_257,
      I1 => rx_input_memio_macnt_inst_lut3_60,
      O => rx_input_memio_macnt_inst_sum_223
    );
  rx_input_memio_macnt_73_CYINIT_683 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_256,
      O => rx_input_memio_macnt_73_CYINIT
    );
  mac_control_rxoferr_cnt_18_LOGIC_ZERO_684 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_18_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_34_685 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_18_CYINIT,
      SEL => mac_control_rxoferr_cnt_18_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_18_CYINIT,
      I1 => mac_control_rxoferr_cnt_18_FROM,
      O => mac_control_rxoferr_cnt_n0000(18)
    );
  mac_control_rxoferr_cnt_18_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(18),
      O => mac_control_rxoferr_cnt_18_FROM
    );
  mac_control_rxoferr_cnt_18_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(19),
      O => mac_control_rxoferr_cnt_18_GROM
    );
  mac_control_rxoferr_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_18_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_35_686 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_rxoferr_cnt_18_GROM,
      O => mac_control_rxoferr_cnt_18_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_rxoferr_cnt_18_GROM,
      O => mac_control_rxoferr_cnt_n0000(19)
    );
  mac_control_rxoferr_cnt_18_CYINIT_687 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_rxoferr_cnt_18_CYINIT
    );
  rx_input_memio_dout_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_n0044,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_7_FFX_RST,
      O => rx_input_memio_dout(7)
    );
  rx_input_memio_dout_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_7_FFX_RST
    );
  mac_control_rxoferr_cnt_20_LOGIC_ZERO_688 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_20_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_36_689 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_20_CYINIT,
      SEL => mac_control_rxoferr_cnt_20_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_20_CYINIT,
      I1 => mac_control_rxoferr_cnt_20_FROM,
      O => mac_control_rxoferr_cnt_n0000(20)
    );
  mac_control_rxoferr_cnt_20_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(20),
      O => mac_control_rxoferr_cnt_20_FROM
    );
  mac_control_rxoferr_cnt_20_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(21),
      O => mac_control_rxoferr_cnt_20_GROM
    );
  mac_control_rxoferr_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_20_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_37_690 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_rxoferr_cnt_20_GROM,
      O => mac_control_rxoferr_cnt_20_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_rxoferr_cnt_20_GROM,
      O => mac_control_rxoferr_cnt_n0000(21)
    );
  mac_control_rxoferr_cnt_20_CYINIT_691 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_rxoferr_cnt_20_CYINIT
    );
  mac_control_rxoferr_cnt_22_LOGIC_ZERO_692 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_22_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_38_693 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_22_CYINIT,
      SEL => mac_control_rxoferr_cnt_22_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_22_CYINIT,
      I1 => mac_control_rxoferr_cnt_22_FROM,
      O => mac_control_rxoferr_cnt_n0000(22)
    );
  mac_control_rxoferr_cnt_22_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(22),
      O => mac_control_rxoferr_cnt_22_FROM
    );
  mac_control_rxoferr_cnt_22_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(23),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_22_GROM
    );
  mac_control_rxoferr_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_22_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_39_694 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_rxoferr_cnt_22_GROM,
      O => mac_control_rxoferr_cnt_22_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_rxoferr_cnt_22_GROM,
      O => mac_control_rxoferr_cnt_n0000(23)
    );
  mac_control_rxoferr_cnt_22_CYINIT_695 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_rxoferr_cnt_22_CYINIT
    );
  mac_control_rxoferr_cnt_24_LOGIC_ZERO_696 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_24_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_40_697 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_24_CYINIT,
      SEL => mac_control_rxoferr_cnt_24_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_24_CYINIT,
      I1 => mac_control_rxoferr_cnt_24_FROM,
      O => mac_control_rxoferr_cnt_n0000(24)
    );
  mac_control_rxoferr_cnt_24_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(24),
      O => mac_control_rxoferr_cnt_24_FROM
    );
  mac_control_rxoferr_cnt_24_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxoferr_cnt(25),
      ADR3 => VCC,
      O => mac_control_rxoferr_cnt_24_GROM
    );
  mac_control_rxoferr_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_24_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_41_698 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_rxoferr_cnt_24_GROM,
      O => mac_control_rxoferr_cnt_24_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_rxoferr_cnt_24_GROM,
      O => mac_control_rxoferr_cnt_n0000(25)
    );
  mac_control_rxoferr_cnt_24_CYINIT_699 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_rxoferr_cnt_24_CYINIT
    );
  mac_control_rxoferr_cnt_26_LOGIC_ZERO_700 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_26_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_42_701 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_26_CYINIT,
      SEL => mac_control_rxoferr_cnt_26_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_26_CYINIT,
      I1 => mac_control_rxoferr_cnt_26_FROM,
      O => mac_control_rxoferr_cnt_n0000(26)
    );
  mac_control_rxoferr_cnt_26_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(26),
      O => mac_control_rxoferr_cnt_26_FROM
    );
  mac_control_rxoferr_cnt_26_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(27),
      O => mac_control_rxoferr_cnt_26_GROM
    );
  mac_control_rxoferr_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_26_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_43_702 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_rxoferr_cnt_26_GROM,
      O => mac_control_rxoferr_cnt_26_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_rxoferr_cnt_26_GROM,
      O => mac_control_rxoferr_cnt_n0000(27)
    );
  mac_control_rxoferr_cnt_26_CYINIT_703 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_rxoferr_cnt_26_CYINIT
    );
  mac_control_rxoferr_cnt_28_LOGIC_ZERO_704 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_28_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_44_705 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_28_CYINIT,
      SEL => mac_control_rxoferr_cnt_28_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_28_CYINIT,
      I1 => mac_control_rxoferr_cnt_28_FROM,
      O => mac_control_rxoferr_cnt_n0000(28)
    );
  mac_control_rxoferr_cnt_28_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(28),
      O => mac_control_rxoferr_cnt_28_FROM
    );
  mac_control_rxoferr_cnt_28_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(29),
      O => mac_control_rxoferr_cnt_28_GROM
    );
  mac_control_rxoferr_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_28_CYMUXG,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_45_706 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_rxoferr_cnt_28_GROM,
      O => mac_control_rxoferr_cnt_28_CYMUXG
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_rxoferr_cnt_28_GROM,
      O => mac_control_rxoferr_cnt_n0000(29)
    );
  mac_control_rxoferr_cnt_28_CYINIT_707 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_rxoferr_cnt_28_CYINIT
    );
  mac_control_rxoferr_cnt_30_LOGIC_ZERO_708 : X_ZERO
    port map (
      O => mac_control_rxoferr_cnt_30_LOGIC_ZERO
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_cy_46_709 : X_MUX2
    port map (
      IA => mac_control_rxoferr_cnt_30_LOGIC_ZERO,
      IB => mac_control_rxoferr_cnt_30_CYINIT,
      SEL => mac_control_rxoferr_cnt_30_FROM,
      O => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_30_CYINIT,
      I1 => mac_control_rxoferr_cnt_30_FROM,
      O => mac_control_rxoferr_cnt_n0000(30)
    );
  mac_control_rxoferr_cnt_30_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(30),
      O => mac_control_rxoferr_cnt_30_FROM
    );
  mac_control_rxoferr_cnt_31_rt_710 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxoferr_cnt(31),
      O => mac_control_rxoferr_cnt_31_rt
    );
  mac_control_rxoferr_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_rxoferr_cnt_31_rt,
      O => mac_control_rxoferr_cnt_n0000(31)
    );
  mac_control_rxoferr_cnt_30_CYINIT_711 : X_BUF
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_rxoferr_cnt_30_CYINIT
    );
  mac_control_ledrx_cnt_154_LOGIC_ONE_712 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_154_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_340_713 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_22,
      IB => mac_control_ledrx_cnt_154_LOGIC_ONE,
      SEL => mac_control_ledrx_rst_rt,
      O => mac_control_ledrx_cnt_inst_cy_340
    );
  mac_control_ledrx_rst_rt_714 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_22,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_rst,
      ADR3 => VCC,
      O => mac_control_ledrx_rst_rt
    );
  mac_control_ledrx_cnt_inst_lut3_2361 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_14,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_rst,
      ADR3 => mac_control_ledrx_cnt_154,
      O => mac_control_ledrx_cnt_inst_lut3_236
    );
  mac_control_ledrx_cnt_154_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_154_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_341
    );
  mac_control_ledrx_cnt_inst_cy_341_715 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_14,
      IB => mac_control_ledrx_cnt_inst_cy_340,
      SEL => mac_control_ledrx_cnt_inst_lut3_236,
      O => mac_control_ledrx_cnt_154_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_301_716 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_340,
      I1 => mac_control_ledrx_cnt_inst_lut3_236,
      O => mac_control_ledrx_cnt_inst_sum_301
    );
  mac_control_ledrx_cnt_155_LOGIC_ONE_717 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_155_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_342_718 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_155_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_155_CYINIT,
      SEL => mac_control_ledrx_cnt_inst_lut3_237,
      O => mac_control_ledrx_cnt_inst_cy_342
    );
  mac_control_ledrx_cnt_inst_sum_302_719 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_155_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_237,
      O => mac_control_ledrx_cnt_inst_sum_302
    );
  mac_control_ledrx_cnt_inst_lut3_2371 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledrx_cnt_155,
      ADR2 => mac_control_ledrx_rst,
      ADR3 => VCC,
      O => mac_control_ledrx_cnt_inst_lut3_237
    );
  mac_control_ledrx_cnt_inst_lut3_2381 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_rst,
      ADR3 => mac_control_ledrx_cnt_156,
      O => mac_control_ledrx_cnt_inst_lut3_238
    );
  mac_control_ledrx_cnt_155_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_155_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_343
    );
  mac_control_ledrx_cnt_inst_cy_343_720 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_155_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_inst_cy_342,
      SEL => mac_control_ledrx_cnt_inst_lut3_238,
      O => mac_control_ledrx_cnt_155_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_303_721 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_342,
      I1 => mac_control_ledrx_cnt_inst_lut3_238,
      O => mac_control_ledrx_cnt_inst_sum_303
    );
  mac_control_ledrx_cnt_155_CYINIT_722 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_341,
      O => mac_control_ledrx_cnt_155_CYINIT
    );
  mac_control_ledrx_cnt_157_LOGIC_ONE_723 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_157_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_344_724 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_157_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_157_CYINIT,
      SEL => mac_control_ledrx_cnt_inst_lut3_239,
      O => mac_control_ledrx_cnt_inst_cy_344
    );
  mac_control_ledrx_cnt_inst_sum_304_725 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_157_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_239,
      O => mac_control_ledrx_cnt_inst_sum_304
    );
  mac_control_ledrx_cnt_inst_lut3_2391 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_ledrx_rst,
      ADR1 => mac_control_ledrx_cnt_157,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledrx_cnt_inst_lut3_239
    );
  mac_control_ledrx_cnt_inst_lut3_2401 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_ledrx_rst,
      ADR1 => mac_control_ledrx_cnt_158,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledrx_cnt_inst_lut3_240
    );
  mac_control_ledrx_cnt_157_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_157_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_345
    );
  mac_control_ledrx_cnt_inst_cy_345_726 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_157_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_inst_cy_344,
      SEL => mac_control_ledrx_cnt_inst_lut3_240,
      O => mac_control_ledrx_cnt_157_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_305_727 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_344,
      I1 => mac_control_ledrx_cnt_inst_lut3_240,
      O => mac_control_ledrx_cnt_inst_sum_305
    );
  mac_control_ledrx_cnt_157_CYINIT_728 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_343,
      O => mac_control_ledrx_cnt_157_CYINIT
    );
  mac_control_ledrx_cnt_159_LOGIC_ONE_729 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_159_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_346_730 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_159_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_159_CYINIT,
      SEL => mac_control_ledrx_cnt_inst_lut3_241,
      O => mac_control_ledrx_cnt_inst_cy_346
    );
  mac_control_ledrx_cnt_inst_sum_306_731 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_159_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_241,
      O => mac_control_ledrx_cnt_inst_sum_306
    );
  mac_control_ledrx_cnt_inst_lut3_2411 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_cnt_159,
      ADR3 => mac_control_ledrx_rst,
      O => mac_control_ledrx_cnt_inst_lut3_241
    );
  mac_control_ledrx_cnt_inst_lut3_2421 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => mac_control_ledrx_rst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_ledrx_cnt_160,
      O => mac_control_ledrx_cnt_inst_lut3_242
    );
  mac_control_ledrx_cnt_159_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_159_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_347
    );
  mac_control_ledrx_cnt_inst_cy_347_732 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_159_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_inst_cy_346,
      SEL => mac_control_ledrx_cnt_inst_lut3_242,
      O => mac_control_ledrx_cnt_159_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_307_733 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_346,
      I1 => mac_control_ledrx_cnt_inst_lut3_242,
      O => mac_control_ledrx_cnt_inst_sum_307
    );
  mac_control_ledrx_cnt_159_CYINIT_734 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_345,
      O => mac_control_ledrx_cnt_159_CYINIT
    );
  mac_control_ledrx_cnt_161_LOGIC_ONE_735 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_161_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_348_736 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_161_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_161_CYINIT,
      SEL => mac_control_ledrx_cnt_inst_lut3_243,
      O => mac_control_ledrx_cnt_inst_cy_348
    );
  mac_control_ledrx_cnt_inst_sum_308_737 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_161_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_243,
      O => mac_control_ledrx_cnt_inst_sum_308
    );
  mac_control_ledrx_cnt_inst_lut3_2431 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => mac_control_ledrx_cnt_161,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_ledrx_rst,
      O => mac_control_ledrx_cnt_inst_lut3_243
    );
  mac_control_ledrx_cnt_inst_lut3_2441 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_cnt_162,
      ADR3 => mac_control_ledrx_rst,
      O => mac_control_ledrx_cnt_inst_lut3_244
    );
  mac_control_ledrx_cnt_161_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_161_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_349
    );
  mac_control_ledrx_cnt_inst_cy_349_738 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_161_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_inst_cy_348,
      SEL => mac_control_ledrx_cnt_inst_lut3_244,
      O => mac_control_ledrx_cnt_161_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_309_739 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_348,
      I1 => mac_control_ledrx_cnt_inst_lut3_244,
      O => mac_control_ledrx_cnt_inst_sum_309
    );
  mac_control_ledrx_cnt_161_CYINIT_740 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_347,
      O => mac_control_ledrx_cnt_161_CYINIT
    );
  rx_input_memio_dout_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_9_FFX_RST,
      O => rx_input_memio_dout(9)
    );
  rx_input_memio_dout_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_9_FFX_RST
    );
  mac_control_ledrx_cnt_163_LOGIC_ONE_741 : X_ONE
    port map (
      O => mac_control_ledrx_cnt_163_LOGIC_ONE
    );
  mac_control_ledrx_cnt_inst_cy_350_742 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_163_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_163_CYINIT,
      SEL => mac_control_ledrx_cnt_inst_lut3_245,
      O => mac_control_ledrx_cnt_inst_cy_350
    );
  mac_control_ledrx_cnt_inst_sum_310_743 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_163_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_245,
      O => mac_control_ledrx_cnt_inst_sum_310
    );
  mac_control_ledrx_cnt_inst_lut3_2451 : X_LUT4
    generic map(
      INIT => X"0033"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledrx_rst,
      ADR2 => VCC,
      ADR3 => mac_control_ledrx_cnt_163,
      O => mac_control_ledrx_cnt_inst_lut3_245
    );
  mac_control_ledrx_cnt_inst_lut3_2461 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledrx_rst,
      ADR3 => mac_control_ledrx_cnt_164,
      O => mac_control_ledrx_cnt_inst_lut3_246
    );
  mac_control_ledrx_cnt_163_COUTUSED : X_BUF
    port map (
      I => mac_control_ledrx_cnt_163_CYMUXG,
      O => mac_control_ledrx_cnt_inst_cy_351
    );
  mac_control_ledrx_cnt_inst_cy_351_744 : X_MUX2
    port map (
      IA => mac_control_ledrx_cnt_163_LOGIC_ONE,
      IB => mac_control_ledrx_cnt_inst_cy_350,
      SEL => mac_control_ledrx_cnt_inst_lut3_246,
      O => mac_control_ledrx_cnt_163_CYMUXG
    );
  mac_control_ledrx_cnt_inst_sum_311_745 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_inst_cy_350,
      I1 => mac_control_ledrx_cnt_inst_lut3_246,
      O => mac_control_ledrx_cnt_inst_sum_311
    );
  mac_control_ledrx_cnt_163_CYINIT_746 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_349,
      O => mac_control_ledrx_cnt_163_CYINIT
    );
  mac_control_ledrx_cnt_inst_sum_312_747 : X_XOR2
    port map (
      I0 => mac_control_ledrx_cnt_165_CYINIT,
      I1 => mac_control_ledrx_cnt_inst_lut3_247,
      O => mac_control_ledrx_cnt_inst_sum_312
    );
  mac_control_ledrx_cnt_inst_lut3_2471 : X_LUT4
    generic map(
      INIT => X"1111"
    )
    port map (
      ADR0 => mac_control_ledrx_rst,
      ADR1 => mac_control_ledrx_cnt_165,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledrx_cnt_inst_lut3_247
    );
  mac_control_ledrx_cnt_165_CYINIT_748 : X_BUF
    port map (
      I => mac_control_ledrx_cnt_inst_cy_351,
      O => mac_control_ledrx_cnt_165_CYINIT
    );
  tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ONE_749 : X_ONE
    port map (
      O => tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ONE
    );
  tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ZERO_750 : X_ZERO
    port map (
      O => tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ZERO
    );
  tx_output_Mcompar_n0035_inst_cy_194_751 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ONE,
      SEL => tx_output_bcntl_1_rt,
      O => tx_output_Mcompar_n0035_inst_cy_194
    );
  tx_output_bcntl_1_rt_752 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => tx_output_bcntl(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_output_bcntl_1_rt
    );
  tx_output_BEL_0 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_bcntl(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_output_SIG_19
    );
  tx_output_Mcompar_n0035_inst_cy_195_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_195_CYMUXG,
      O => tx_output_Mcompar_n0035_inst_cy_195
    );
  tx_output_Mcompar_n0035_inst_cy_195_753 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_195_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0035_inst_cy_194,
      SEL => tx_output_SIG_19,
      O => tx_output_Mcompar_n0035_inst_cy_195_CYMUXG
    );
  tx_output_Mcompar_n0035_inst_cy_197_LOGIC_ONE_754 : X_ONE
    port map (
      O => tx_output_Mcompar_n0035_inst_cy_197_LOGIC_ONE
    );
  tx_output_Mcompar_n0035_inst_cy_196_755 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_197_LOGIC_ONE,
      IB => tx_output_Mcompar_n0035_inst_cy_197_CYINIT,
      SEL => tx_output_Mcompar_n0035_inst_lut1_61_O,
      O => tx_output_Mcompar_n0035_inst_cy_196
    );
  tx_output_Mcompar_n0035_inst_lut1_61 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_bcntl(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_output_Mcompar_n0035_inst_lut1_61_O
    );
  tx_output_Mcompar_n0035_inst_lut1_71 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_bcntl(2),
      ADR3 => VCC,
      O => tx_output_Mcompar_n0035_inst_lut1_71_O
    );
  tx_output_Mcompar_n0035_inst_cy_197_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_197_CYMUXG,
      O => tx_output_Mcompar_n0035_inst_cy_197
    );
  tx_output_Mcompar_n0035_inst_cy_197_756 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_197_LOGIC_ONE,
      IB => tx_output_Mcompar_n0035_inst_cy_196,
      SEL => tx_output_Mcompar_n0035_inst_lut1_71_O,
      O => tx_output_Mcompar_n0035_inst_cy_197_CYMUXG
    );
  tx_output_Mcompar_n0035_inst_cy_197_CYINIT_757 : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_195,
      O => tx_output_Mcompar_n0035_inst_cy_197_CYINIT
    );
  tx_output_Mcompar_n0035_inst_cy_199_LOGIC_ZERO_758 : X_ZERO
    port map (
      O => tx_output_Mcompar_n0035_inst_cy_199_LOGIC_ZERO
    );
  tx_output_Mcompar_n0035_inst_cy_198_759 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_199_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0035_inst_cy_199_CYINIT,
      SEL => tx_output_bcntl_3_rt,
      O => tx_output_Mcompar_n0035_inst_cy_198
    );
  tx_output_bcntl_3_rt_760 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_bcntl(3),
      O => tx_output_bcntl_3_rt
    );
  tx_output_BEL_1 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_bcntl(3),
      O => tx_output_SIG_20
    );
  tx_output_Mcompar_n0035_inst_cy_199_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_199_CYMUXG,
      O => tx_output_Mcompar_n0035_inst_cy_199
    );
  tx_output_Mcompar_n0035_inst_cy_199_761 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_199_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0035_inst_cy_198,
      SEL => tx_output_SIG_20,
      O => tx_output_Mcompar_n0035_inst_cy_199_CYMUXG
    );
  tx_output_Mcompar_n0035_inst_cy_199_CYINIT_762 : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_197,
      O => tx_output_Mcompar_n0035_inst_cy_199_CYINIT
    );
  tx_output_Mcompar_n0035_inst_cy_201_LOGIC_ONE_763 : X_ONE
    port map (
      O => tx_output_Mcompar_n0035_inst_cy_201_LOGIC_ONE
    );
  tx_output_Mcompar_n0035_inst_cy_200_764 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_201_LOGIC_ONE,
      IB => tx_output_Mcompar_n0035_inst_cy_201_CYINIT,
      SEL => tx_output_Mcompar_n0035_inst_lut4_161_O,
      O => tx_output_Mcompar_n0035_inst_cy_200
    );
  tx_output_Mcompar_n0035_inst_lut4_161 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcntl(4),
      ADR1 => tx_output_bcntl(6),
      ADR2 => tx_output_bcntl(5),
      ADR3 => tx_output_bcntl(7),
      O => tx_output_Mcompar_n0035_inst_lut4_161_O
    );
  tx_output_Mcompar_n0035_inst_lut4_171 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcntl(7),
      ADR1 => tx_output_bcntl(5),
      ADR2 => tx_output_bcntl(4),
      ADR3 => tx_output_bcntl(6),
      O => tx_output_Mcompar_n0035_inst_lut4_171_O
    );
  tx_output_Mcompar_n0035_inst_cy_201_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_201_CYMUXG,
      O => tx_output_Mcompar_n0035_inst_cy_201
    );
  tx_output_Mcompar_n0035_inst_cy_201_765 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0035_inst_cy_201_LOGIC_ONE,
      IB => tx_output_Mcompar_n0035_inst_cy_200,
      SEL => tx_output_Mcompar_n0035_inst_lut4_171_O,
      O => tx_output_Mcompar_n0035_inst_cy_201_CYMUXG
    );
  tx_output_Mcompar_n0035_inst_cy_201_CYINIT_766 : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_199,
      O => tx_output_Mcompar_n0035_inst_cy_201_CYINIT
    );
  tx_output_n0035_LOGIC_ONE_767 : X_ONE
    port map (
      O => tx_output_n0035_LOGIC_ONE
    );
  tx_output_Mcompar_n0035_inst_cy_202_768 : X_MUX2
    port map (
      IA => tx_output_n0035_LOGIC_ONE,
      IB => tx_output_n0035_CYINIT,
      SEL => tx_output_Mcompar_n0035_inst_lut4_18,
      O => tx_output_Mcompar_n0035_inst_cy_202
    );
  tx_output_Mcompar_n0035_inst_lut4_181 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcntl(10),
      ADR1 => tx_output_bcntl(9),
      ADR2 => tx_output_bcntl(8),
      ADR3 => tx_output_bcntl(11),
      O => tx_output_Mcompar_n0035_inst_lut4_18
    );
  tx_output_Mcompar_n0035_inst_lut4_191 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_bcntl(13),
      ADR1 => tx_output_bcntl(14),
      ADR2 => tx_output_bcntl(15),
      ADR3 => tx_output_bcntl(12),
      O => tx_output_Mcompar_n0035_inst_lut4_19
    );
  tx_output_n0035_COUTUSED : X_BUF
    port map (
      I => tx_output_n0035_CYMUXG,
      O => tx_output_n0035
    );
  tx_output_Mcompar_n0035_inst_cy_203 : X_MUX2
    port map (
      IA => tx_output_n0035_LOGIC_ONE,
      IB => tx_output_Mcompar_n0035_inst_cy_202,
      SEL => tx_output_Mcompar_n0035_inst_lut4_19,
      O => tx_output_n0035_CYMUXG
    );
  tx_output_n0035_CYINIT_769 : X_BUF
    port map (
      I => tx_output_Mcompar_n0035_inst_cy_201,
      O => tx_output_n0035_CYINIT
    );
  mac_control_rxphyerr_cnt_0_LOGIC_ZERO_770 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_0_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_16_771 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_24,
      IB => mac_control_rxphyerr_cnt_0_LOGIC_ZERO,
      SEL => mac_control_rxphyerr_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_24,
      ADR1 => mac_control_rxphyerr_cnt(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_rxphyerr_cnt_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_37,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(1),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_0_GROM
    );
  mac_control_rxphyerr_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_0_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_17_772 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_37,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_rxphyerr_cnt_0_GROM,
      O => mac_control_rxphyerr_cnt_0_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_rxphyerr_cnt_0_GROM,
      O => mac_control_rxphyerr_cnt_n0000(1)
    );
  mac_control_rxphyerr_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(3),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(3)
    );
  mac_control_rxphyerr_cnt_2_LOGIC_ZERO_773 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_2_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_18_774 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_2_CYINIT,
      SEL => mac_control_rxphyerr_cnt_2_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_2_CYINIT,
      I1 => mac_control_rxphyerr_cnt_2_FROM,
      O => mac_control_rxphyerr_cnt_n0000(2)
    );
  mac_control_rxphyerr_cnt_2_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_2_FROM
    );
  mac_control_rxphyerr_cnt_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxphyerr_cnt(3),
      O => mac_control_rxphyerr_cnt_2_GROM
    );
  mac_control_rxphyerr_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_2_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_19_775 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_rxphyerr_cnt_2_GROM,
      O => mac_control_rxphyerr_cnt_2_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_rxphyerr_cnt_2_GROM,
      O => mac_control_rxphyerr_cnt_n0000(3)
    );
  mac_control_rxphyerr_cnt_2_CYINIT_776 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_rxphyerr_cnt_2_CYINIT
    );
  mac_control_rxphyerr_cnt_4_LOGIC_ZERO_777 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_4_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_20_778 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_4_CYINIT,
      SEL => mac_control_rxphyerr_cnt_4_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_4_CYINIT,
      I1 => mac_control_rxphyerr_cnt_4_FROM,
      O => mac_control_rxphyerr_cnt_n0000(4)
    );
  mac_control_rxphyerr_cnt_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_4_FROM
    );
  mac_control_rxphyerr_cnt_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(5),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_4_GROM
    );
  mac_control_rxphyerr_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_4_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_21_779 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_rxphyerr_cnt_4_GROM,
      O => mac_control_rxphyerr_cnt_4_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_rxphyerr_cnt_4_GROM,
      O => mac_control_rxphyerr_cnt_n0000(5)
    );
  mac_control_rxphyerr_cnt_4_CYINIT_780 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_rxphyerr_cnt_4_CYINIT
    );
  mac_control_rxphyerr_cnt_6_LOGIC_ZERO_781 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_6_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_22_782 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_6_CYINIT,
      SEL => mac_control_rxphyerr_cnt_6_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_6_CYINIT,
      I1 => mac_control_rxphyerr_cnt_6_FROM,
      O => mac_control_rxphyerr_cnt_n0000(6)
    );
  mac_control_rxphyerr_cnt_6_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_6_FROM
    );
  mac_control_rxphyerr_cnt_6_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(7),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_6_GROM
    );
  mac_control_rxphyerr_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_6_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_23_783 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_rxphyerr_cnt_6_GROM,
      O => mac_control_rxphyerr_cnt_6_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_rxphyerr_cnt_6_GROM,
      O => mac_control_rxphyerr_cnt_n0000(7)
    );
  mac_control_rxphyerr_cnt_6_CYINIT_784 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_rxphyerr_cnt_6_CYINIT
    );
  mac_control_rxphyerr_cnt_8_LOGIC_ZERO_785 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_8_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_24_786 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_8_CYINIT,
      SEL => mac_control_rxphyerr_cnt_8_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_8_CYINIT,
      I1 => mac_control_rxphyerr_cnt_8_FROM,
      O => mac_control_rxphyerr_cnt_n0000(8)
    );
  mac_control_rxphyerr_cnt_8_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_8_FROM
    );
  mac_control_rxphyerr_cnt_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(9),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_8_GROM
    );
  mac_control_rxphyerr_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_8_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_25_787 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_rxphyerr_cnt_8_GROM,
      O => mac_control_rxphyerr_cnt_8_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_rxphyerr_cnt_8_GROM,
      O => mac_control_rxphyerr_cnt_n0000(9)
    );
  mac_control_rxphyerr_cnt_8_CYINIT_788 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_rxphyerr_cnt_8_CYINIT
    );
  mac_control_rxphyerr_cnt_10_LOGIC_ZERO_789 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_10_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_26_790 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_10_CYINIT,
      SEL => mac_control_rxphyerr_cnt_10_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_10_CYINIT,
      I1 => mac_control_rxphyerr_cnt_10_FROM,
      O => mac_control_rxphyerr_cnt_n0000(10)
    );
  mac_control_rxphyerr_cnt_10_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_10_FROM
    );
  mac_control_rxphyerr_cnt_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(11),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_10_GROM
    );
  mac_control_rxphyerr_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_10_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_27_791 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_rxphyerr_cnt_10_GROM,
      O => mac_control_rxphyerr_cnt_10_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_rxphyerr_cnt_10_GROM,
      O => mac_control_rxphyerr_cnt_n0000(11)
    );
  mac_control_rxphyerr_cnt_10_CYINIT_792 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_rxphyerr_cnt_10_CYINIT
    );
  mac_control_rxphyerr_cnt_12_LOGIC_ZERO_793 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_12_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_28_794 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_12_CYINIT,
      SEL => mac_control_rxphyerr_cnt_12_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_12_CYINIT,
      I1 => mac_control_rxphyerr_cnt_12_FROM,
      O => mac_control_rxphyerr_cnt_n0000(12)
    );
  mac_control_rxphyerr_cnt_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_12_FROM
    );
  mac_control_rxphyerr_cnt_12_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(13),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_12_GROM
    );
  mac_control_rxphyerr_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_12_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_29_795 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_rxphyerr_cnt_12_GROM,
      O => mac_control_rxphyerr_cnt_12_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_rxphyerr_cnt_12_GROM,
      O => mac_control_rxphyerr_cnt_n0000(13)
    );
  mac_control_rxphyerr_cnt_12_CYINIT_796 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_rxphyerr_cnt_12_CYINIT
    );
  mac_control_rxphyerr_cnt_14_LOGIC_ZERO_797 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_14_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_30_798 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_14_CYINIT,
      SEL => mac_control_rxphyerr_cnt_14_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_14_CYINIT,
      I1 => mac_control_rxphyerr_cnt_14_FROM,
      O => mac_control_rxphyerr_cnt_n0000(14)
    );
  mac_control_rxphyerr_cnt_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_14_FROM
    );
  mac_control_rxphyerr_cnt_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(15),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_14_GROM
    );
  mac_control_rxphyerr_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_14_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_31_799 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_rxphyerr_cnt_14_GROM,
      O => mac_control_rxphyerr_cnt_14_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_rxphyerr_cnt_14_GROM,
      O => mac_control_rxphyerr_cnt_n0000(15)
    );
  mac_control_rxphyerr_cnt_14_CYINIT_800 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_rxphyerr_cnt_14_CYINIT
    );
  mac_control_rxphyerr_cnt_16_LOGIC_ZERO_801 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_16_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_32_802 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_16_CYINIT,
      SEL => mac_control_rxphyerr_cnt_16_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_16_CYINIT,
      I1 => mac_control_rxphyerr_cnt_16_FROM,
      O => mac_control_rxphyerr_cnt_n0000(16)
    );
  mac_control_rxphyerr_cnt_16_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_16_FROM
    );
  mac_control_rxphyerr_cnt_16_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(17),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_16_GROM
    );
  mac_control_rxphyerr_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_16_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_33_803 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_rxphyerr_cnt_16_GROM,
      O => mac_control_rxphyerr_cnt_16_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_rxphyerr_cnt_16_GROM,
      O => mac_control_rxphyerr_cnt_n0000(17)
    );
  mac_control_rxphyerr_cnt_16_CYINIT_804 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_rxphyerr_cnt_16_CYINIT
    );
  mac_control_rxphyerr_cnt_18_LOGIC_ZERO_805 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_18_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_34_806 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_18_CYINIT,
      SEL => mac_control_rxphyerr_cnt_18_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_18_CYINIT,
      I1 => mac_control_rxphyerr_cnt_18_FROM,
      O => mac_control_rxphyerr_cnt_n0000(18)
    );
  mac_control_rxphyerr_cnt_18_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_18_FROM
    );
  mac_control_rxphyerr_cnt_18_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(19),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_18_GROM
    );
  mac_control_rxphyerr_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_18_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_35_807 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_rxphyerr_cnt_18_GROM,
      O => mac_control_rxphyerr_cnt_18_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_rxphyerr_cnt_18_GROM,
      O => mac_control_rxphyerr_cnt_n0000(19)
    );
  mac_control_rxphyerr_cnt_18_CYINIT_808 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_rxphyerr_cnt_18_CYINIT
    );
  mac_control_rxphyerr_cnt_20_LOGIC_ZERO_809 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_20_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_36_810 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_20_CYINIT,
      SEL => mac_control_rxphyerr_cnt_20_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_20_CYINIT,
      I1 => mac_control_rxphyerr_cnt_20_FROM,
      O => mac_control_rxphyerr_cnt_n0000(20)
    );
  mac_control_rxphyerr_cnt_20_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cnt(20),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_20_FROM
    );
  mac_control_rxphyerr_cnt_20_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(21),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_20_GROM
    );
  mac_control_rxphyerr_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_20_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_37_811 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_rxphyerr_cnt_20_GROM,
      O => mac_control_rxphyerr_cnt_20_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_rxphyerr_cnt_20_GROM,
      O => mac_control_rxphyerr_cnt_n0000(21)
    );
  mac_control_rxphyerr_cnt_20_CYINIT_812 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_rxphyerr_cnt_20_CYINIT
    );
  rx_output_cs_FFd5_813 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd5_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd5_FFX_RST,
      O => rx_output_cs_FFd5
    );
  rx_output_cs_FFd5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd5_FFX_RST
    );
  mac_control_rxphyerr_cnt_22_LOGIC_ZERO_814 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_22_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_38_815 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_22_CYINIT,
      SEL => mac_control_rxphyerr_cnt_22_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_22_CYINIT,
      I1 => mac_control_rxphyerr_cnt_22_FROM,
      O => mac_control_rxphyerr_cnt_n0000(22)
    );
  mac_control_rxphyerr_cnt_22_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(22),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_22_FROM
    );
  mac_control_rxphyerr_cnt_22_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(23),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_22_GROM
    );
  mac_control_rxphyerr_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_22_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_39_816 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_rxphyerr_cnt_22_GROM,
      O => mac_control_rxphyerr_cnt_22_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_rxphyerr_cnt_22_GROM,
      O => mac_control_rxphyerr_cnt_n0000(23)
    );
  mac_control_rxphyerr_cnt_22_CYINIT_817 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_rxphyerr_cnt_22_CYINIT
    );
  mac_control_rxphyerr_cnt_24_LOGIC_ZERO_818 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_24_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_40_819 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_24_CYINIT,
      SEL => mac_control_rxphyerr_cnt_24_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_24_CYINIT,
      I1 => mac_control_rxphyerr_cnt_24_FROM,
      O => mac_control_rxphyerr_cnt_n0000(24)
    );
  mac_control_rxphyerr_cnt_24_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(24),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_24_FROM
    );
  mac_control_rxphyerr_cnt_24_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(25),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_24_GROM
    );
  mac_control_rxphyerr_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_24_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_41_820 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_rxphyerr_cnt_24_GROM,
      O => mac_control_rxphyerr_cnt_24_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_rxphyerr_cnt_24_GROM,
      O => mac_control_rxphyerr_cnt_n0000(25)
    );
  mac_control_rxphyerr_cnt_24_CYINIT_821 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_rxphyerr_cnt_24_CYINIT
    );
  mac_control_rxphyerr_cnt_26_LOGIC_ZERO_822 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_26_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_42_823 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_26_CYINIT,
      SEL => mac_control_rxphyerr_cnt_26_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_26_CYINIT,
      I1 => mac_control_rxphyerr_cnt_26_FROM,
      O => mac_control_rxphyerr_cnt_n0000(26)
    );
  mac_control_rxphyerr_cnt_26_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(26),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_26_FROM
    );
  mac_control_rxphyerr_cnt_26_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(27),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_26_GROM
    );
  mac_control_rxphyerr_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_26_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_43_824 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_rxphyerr_cnt_26_GROM,
      O => mac_control_rxphyerr_cnt_26_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_rxphyerr_cnt_26_GROM,
      O => mac_control_rxphyerr_cnt_n0000(27)
    );
  mac_control_rxphyerr_cnt_26_CYINIT_825 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_rxphyerr_cnt_26_CYINIT
    );
  mac_control_rxphyerr_cnt_28_LOGIC_ZERO_826 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_28_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_44_827 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_28_CYINIT,
      SEL => mac_control_rxphyerr_cnt_28_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_28_CYINIT,
      I1 => mac_control_rxphyerr_cnt_28_FROM,
      O => mac_control_rxphyerr_cnt_n0000(28)
    );
  mac_control_rxphyerr_cnt_28_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(28),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_28_FROM
    );
  mac_control_rxphyerr_cnt_28_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(29),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_28_GROM
    );
  mac_control_rxphyerr_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_28_CYMUXG,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_45_828 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_rxphyerr_cnt_28_GROM,
      O => mac_control_rxphyerr_cnt_28_CYMUXG
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_rxphyerr_cnt_28_GROM,
      O => mac_control_rxphyerr_cnt_n0000(29)
    );
  mac_control_rxphyerr_cnt_28_CYINIT_829 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_rxphyerr_cnt_28_CYINIT
    );
  mac_control_rxphyerr_cnt_30_LOGIC_ZERO_830 : X_ZERO
    port map (
      O => mac_control_rxphyerr_cnt_30_LOGIC_ZERO
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_46_831 : X_MUX2
    port map (
      IA => mac_control_rxphyerr_cnt_30_LOGIC_ZERO,
      IB => mac_control_rxphyerr_cnt_30_CYINIT,
      SEL => mac_control_rxphyerr_cnt_30_FROM,
      O => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_30_CYINIT,
      I1 => mac_control_rxphyerr_cnt_30_FROM,
      O => mac_control_rxphyerr_cnt_n0000(30)
    );
  mac_control_rxphyerr_cnt_30_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxphyerr_cnt(30),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_30_FROM
    );
  mac_control_rxphyerr_cnt_31_rt_832 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxphyerr_cnt(31),
      ADR3 => VCC,
      O => mac_control_rxphyerr_cnt_31_rt
    );
  mac_control_rxphyerr_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_rxphyerr_cnt_31_rt,
      O => mac_control_rxphyerr_cnt_n0000(31)
    );
  mac_control_rxphyerr_cnt_30_CYINIT_833 : X_BUF
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_rxphyerr_cnt_30_CYINIT
    );
  mac_control_rxfifowerr_cnt_0_LOGIC_ZERO_834 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_0_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_16_835 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_29,
      IB => mac_control_rxfifowerr_cnt_0_LOGIC_ZERO,
      SEL => mac_control_rxfifowerr_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_29,
      ADR1 => mac_control_rxfifowerr_cnt(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_rxfifowerr_cnt_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_43,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(1),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_0_GROM
    );
  mac_control_rxfifowerr_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_0_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_17_836 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_43,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_rxfifowerr_cnt_0_GROM,
      O => mac_control_rxfifowerr_cnt_0_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_rxfifowerr_cnt_0_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(1)
    );
  mac_control_rxfifowerr_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(3),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(3)
    );
  mac_control_rxfifowerr_cnt_2_LOGIC_ZERO_837 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_2_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_18_838 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_2_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_2_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_2_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_2_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(2)
    );
  mac_control_rxfifowerr_cnt_2_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_2_FROM
    );
  mac_control_rxfifowerr_cnt_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(3),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_2_GROM
    );
  mac_control_rxfifowerr_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_2_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_19_839 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_rxfifowerr_cnt_2_GROM,
      O => mac_control_rxfifowerr_cnt_2_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_rxfifowerr_cnt_2_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(3)
    );
  mac_control_rxfifowerr_cnt_2_CYINIT_840 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_rxfifowerr_cnt_2_CYINIT
    );
  mac_control_rxfifowerr_cnt_4_LOGIC_ZERO_841 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_4_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_20_842 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_4_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_4_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_4_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_4_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(4)
    );
  mac_control_rxfifowerr_cnt_4_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_4_FROM
    );
  mac_control_rxfifowerr_cnt_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(5),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_4_GROM
    );
  mac_control_rxfifowerr_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_4_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_21_843 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_rxfifowerr_cnt_4_GROM,
      O => mac_control_rxfifowerr_cnt_4_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_rxfifowerr_cnt_4_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(5)
    );
  mac_control_rxfifowerr_cnt_4_CYINIT_844 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_rxfifowerr_cnt_4_CYINIT
    );
  mac_control_rxfifowerr_cnt_6_LOGIC_ZERO_845 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_6_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_22_846 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_6_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_6_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_6_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_6_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(6)
    );
  mac_control_rxfifowerr_cnt_6_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_6_FROM
    );
  mac_control_rxfifowerr_cnt_6_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(7),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_6_GROM
    );
  mac_control_rxfifowerr_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_6_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_23_847 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_rxfifowerr_cnt_6_GROM,
      O => mac_control_rxfifowerr_cnt_6_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_rxfifowerr_cnt_6_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(7)
    );
  mac_control_rxfifowerr_cnt_6_CYINIT_848 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_rxfifowerr_cnt_6_CYINIT
    );
  mac_control_rxfifowerr_cnt_8_LOGIC_ZERO_849 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_8_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_24_850 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_8_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_8_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_8_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_8_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(8)
    );
  mac_control_rxfifowerr_cnt_8_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_8_FROM
    );
  mac_control_rxfifowerr_cnt_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(9),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_8_GROM
    );
  mac_control_rxfifowerr_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_8_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_25_851 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_rxfifowerr_cnt_8_GROM,
      O => mac_control_rxfifowerr_cnt_8_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_rxfifowerr_cnt_8_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(9)
    );
  mac_control_rxfifowerr_cnt_8_CYINIT_852 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_rxfifowerr_cnt_8_CYINIT
    );
  mac_control_rxfifowerr_cnt_10_LOGIC_ZERO_853 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_10_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_26_854 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_10_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_10_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_10_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_10_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(10)
    );
  mac_control_rxfifowerr_cnt_10_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_10_FROM
    );
  mac_control_rxfifowerr_cnt_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(11),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_10_GROM
    );
  mac_control_rxfifowerr_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_10_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_27_855 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_rxfifowerr_cnt_10_GROM,
      O => mac_control_rxfifowerr_cnt_10_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_rxfifowerr_cnt_10_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(11)
    );
  mac_control_rxfifowerr_cnt_10_CYINIT_856 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_rxfifowerr_cnt_10_CYINIT
    );
  mac_control_rxfifowerr_cnt_12_LOGIC_ZERO_857 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_12_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_28_858 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_12_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_12_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_12_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_12_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(12)
    );
  mac_control_rxfifowerr_cnt_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_12_FROM
    );
  mac_control_rxfifowerr_cnt_12_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(13),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_12_GROM
    );
  mac_control_rxfifowerr_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_12_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_29_859 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_rxfifowerr_cnt_12_GROM,
      O => mac_control_rxfifowerr_cnt_12_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_rxfifowerr_cnt_12_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(13)
    );
  mac_control_rxfifowerr_cnt_12_CYINIT_860 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_rxfifowerr_cnt_12_CYINIT
    );
  mac_control_rxfifowerr_cnt_14_LOGIC_ZERO_861 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_14_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_30_862 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_14_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_14_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_14_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_14_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(14)
    );
  mac_control_rxfifowerr_cnt_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_14_FROM
    );
  mac_control_rxfifowerr_cnt_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(15),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_14_GROM
    );
  mac_control_rxfifowerr_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_14_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_31_863 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_rxfifowerr_cnt_14_GROM,
      O => mac_control_rxfifowerr_cnt_14_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_rxfifowerr_cnt_14_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(15)
    );
  mac_control_rxfifowerr_cnt_14_CYINIT_864 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_rxfifowerr_cnt_14_CYINIT
    );
  mac_control_rxfifowerr_cnt_16_LOGIC_ZERO_865 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_16_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_32_866 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_16_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_16_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_16_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_16_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(16)
    );
  mac_control_rxfifowerr_cnt_16_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_16_FROM
    );
  mac_control_rxfifowerr_cnt_16_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(17),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_16_GROM
    );
  mac_control_rxfifowerr_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_16_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_33_867 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_rxfifowerr_cnt_16_GROM,
      O => mac_control_rxfifowerr_cnt_16_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_rxfifowerr_cnt_16_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(17)
    );
  mac_control_rxfifowerr_cnt_16_CYINIT_868 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_rxfifowerr_cnt_16_CYINIT
    );
  mac_control_rxfifowerr_cnt_18_LOGIC_ZERO_869 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_18_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_34_870 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_18_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_18_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_18_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_18_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(18)
    );
  mac_control_rxfifowerr_cnt_18_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(18),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_18_FROM
    );
  mac_control_rxfifowerr_cnt_18_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(19),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_18_GROM
    );
  mac_control_rxfifowerr_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_18_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_35_871 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_rxfifowerr_cnt_18_GROM,
      O => mac_control_rxfifowerr_cnt_18_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_rxfifowerr_cnt_18_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(19)
    );
  mac_control_rxfifowerr_cnt_18_CYINIT_872 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_rxfifowerr_cnt_18_CYINIT
    );
  rx_input_fifo_control_DATA_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(0),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_0_FFY_RST,
      O => rx_input_data(0)
    );
  rx_input_data_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_0_FFY_RST
    );
  mac_control_rxfifowerr_cnt_20_LOGIC_ZERO_873 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_20_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_36_874 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_20_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_20_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_20_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_20_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(20)
    );
  mac_control_rxfifowerr_cnt_20_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(20),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_20_FROM
    );
  mac_control_rxfifowerr_cnt_20_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(21),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_20_GROM
    );
  mac_control_rxfifowerr_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_20_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_37_875 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_rxfifowerr_cnt_20_GROM,
      O => mac_control_rxfifowerr_cnt_20_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_rxfifowerr_cnt_20_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(21)
    );
  mac_control_rxfifowerr_cnt_20_CYINIT_876 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_rxfifowerr_cnt_20_CYINIT
    );
  mac_control_rxfifowerr_cnt_22_LOGIC_ZERO_877 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_22_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_38_878 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_22_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_22_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_22_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_22_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(22)
    );
  mac_control_rxfifowerr_cnt_22_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(22),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_22_FROM
    );
  mac_control_rxfifowerr_cnt_22_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(23),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_22_GROM
    );
  mac_control_rxfifowerr_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_22_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_39_879 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_rxfifowerr_cnt_22_GROM,
      O => mac_control_rxfifowerr_cnt_22_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_rxfifowerr_cnt_22_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(23)
    );
  mac_control_rxfifowerr_cnt_22_CYINIT_880 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_rxfifowerr_cnt_22_CYINIT
    );
  mac_control_rxfifowerr_cnt_24_LOGIC_ZERO_881 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_24_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_40_882 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_24_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_24_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_24_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_24_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(24)
    );
  mac_control_rxfifowerr_cnt_24_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(24),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_24_FROM
    );
  mac_control_rxfifowerr_cnt_24_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(25),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_24_GROM
    );
  mac_control_rxfifowerr_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_24_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_41_883 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_rxfifowerr_cnt_24_GROM,
      O => mac_control_rxfifowerr_cnt_24_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_rxfifowerr_cnt_24_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(25)
    );
  mac_control_rxfifowerr_cnt_24_CYINIT_884 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_rxfifowerr_cnt_24_CYINIT
    );
  mac_control_rxfifowerr_cnt_26_LOGIC_ZERO_885 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_26_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_42_886 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_26_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_26_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_26_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_26_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(26)
    );
  mac_control_rxfifowerr_cnt_26_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(26),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_26_FROM
    );
  mac_control_rxfifowerr_cnt_26_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(27),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_26_GROM
    );
  mac_control_rxfifowerr_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_26_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_43_887 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_rxfifowerr_cnt_26_GROM,
      O => mac_control_rxfifowerr_cnt_26_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_rxfifowerr_cnt_26_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(27)
    );
  mac_control_rxfifowerr_cnt_26_CYINIT_888 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_rxfifowerr_cnt_26_CYINIT
    );
  mac_control_rxfifowerr_cnt_28_LOGIC_ZERO_889 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_28_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_44_890 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_28_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_28_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_28_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_28_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(28)
    );
  mac_control_rxfifowerr_cnt_28_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxfifowerr_cnt(28),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_28_FROM
    );
  mac_control_rxfifowerr_cnt_28_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(29),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_28_GROM
    );
  mac_control_rxfifowerr_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_28_CYMUXG,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_45_891 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_rxfifowerr_cnt_28_GROM,
      O => mac_control_rxfifowerr_cnt_28_CYMUXG
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_rxfifowerr_cnt_28_GROM,
      O => mac_control_rxfifowerr_cnt_n0000(29)
    );
  mac_control_rxfifowerr_cnt_28_CYINIT_892 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_rxfifowerr_cnt_28_CYINIT
    );
  mac_control_rxfifowerr_cnt_30_LOGIC_ZERO_893 : X_ZERO
    port map (
      O => mac_control_rxfifowerr_cnt_30_LOGIC_ZERO
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_46_894 : X_MUX2
    port map (
      IA => mac_control_rxfifowerr_cnt_30_LOGIC_ZERO,
      IB => mac_control_rxfifowerr_cnt_30_CYINIT,
      SEL => mac_control_rxfifowerr_cnt_30_FROM,
      O => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_30_CYINIT,
      I1 => mac_control_rxfifowerr_cnt_30_FROM,
      O => mac_control_rxfifowerr_cnt_n0000(30)
    );
  mac_control_rxfifowerr_cnt_30_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cnt(30),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_30_FROM
    );
  mac_control_rxfifowerr_cnt_31_rt_895 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxfifowerr_cnt(31),
      ADR3 => VCC,
      O => mac_control_rxfifowerr_cnt_31_rt
    );
  mac_control_rxfifowerr_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_rxfifowerr_cnt_31_rt,
      O => mac_control_rxfifowerr_cnt_n0000(31)
    );
  mac_control_rxfifowerr_cnt_30_CYINIT_896 : X_BUF
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_rxfifowerr_cnt_30_CYINIT
    );
  mac_control_txfifowerr_cnt_0_LOGIC_ZERO_897 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_0_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_16_898 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_15,
      IB => mac_control_txfifowerr_cnt_0_LOGIC_ZERO,
      SEL => mac_control_txfifowerr_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"3333"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_15,
      ADR1 => mac_control_txfifowerr_cnt(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_txfifowerr_cnt_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_25,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(1),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_0_GROM
    );
  mac_control_txfifowerr_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_0_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_17_899 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_25,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_txfifowerr_cnt_0_GROM,
      O => mac_control_txfifowerr_cnt_0_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_txfifowerr_cnt_0_GROM,
      O => mac_control_txfifowerr_cnt_n0000(1)
    );
  mac_control_txfifowerr_cnt_2_LOGIC_ZERO_900 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_2_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_18_901 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_2_CYINIT,
      SEL => mac_control_txfifowerr_cnt_2_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_2_CYINIT,
      I1 => mac_control_txfifowerr_cnt_2_FROM,
      O => mac_control_txfifowerr_cnt_n0000(2)
    );
  mac_control_txfifowerr_cnt_2_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_2_FROM
    );
  mac_control_txfifowerr_cnt_2_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(3),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_2_GROM
    );
  mac_control_txfifowerr_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_2_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_19_902 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_2_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_txfifowerr_cnt_2_GROM,
      O => mac_control_txfifowerr_cnt_2_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_txfifowerr_cnt_2_GROM,
      O => mac_control_txfifowerr_cnt_n0000(3)
    );
  mac_control_txfifowerr_cnt_2_CYINIT_903 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_txfifowerr_cnt_2_CYINIT
    );
  mac_control_txfifowerr_cnt_4_LOGIC_ZERO_904 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_4_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_20_905 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_4_CYINIT,
      SEL => mac_control_txfifowerr_cnt_4_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_4_CYINIT,
      I1 => mac_control_txfifowerr_cnt_4_FROM,
      O => mac_control_txfifowerr_cnt_n0000(4)
    );
  mac_control_txfifowerr_cnt_4_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_4_FROM
    );
  mac_control_txfifowerr_cnt_4_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(5),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_4_GROM
    );
  mac_control_txfifowerr_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_4_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_21_906 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_4_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_txfifowerr_cnt_4_GROM,
      O => mac_control_txfifowerr_cnt_4_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_txfifowerr_cnt_4_GROM,
      O => mac_control_txfifowerr_cnt_n0000(5)
    );
  mac_control_txfifowerr_cnt_4_CYINIT_907 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_txfifowerr_cnt_4_CYINIT
    );
  mac_control_txfifowerr_cnt_6_LOGIC_ZERO_908 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_6_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_22_909 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_6_CYINIT,
      SEL => mac_control_txfifowerr_cnt_6_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_6_CYINIT,
      I1 => mac_control_txfifowerr_cnt_6_FROM,
      O => mac_control_txfifowerr_cnt_n0000(6)
    );
  mac_control_txfifowerr_cnt_6_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_6_FROM
    );
  mac_control_txfifowerr_cnt_6_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(7),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_6_GROM
    );
  mac_control_txfifowerr_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_6_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_23_910 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_6_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_txfifowerr_cnt_6_GROM,
      O => mac_control_txfifowerr_cnt_6_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_txfifowerr_cnt_6_GROM,
      O => mac_control_txfifowerr_cnt_n0000(7)
    );
  mac_control_txfifowerr_cnt_6_CYINIT_911 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_txfifowerr_cnt_6_CYINIT
    );
  mac_control_txfifowerr_cnt_8_LOGIC_ZERO_912 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_8_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_24_913 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_8_CYINIT,
      SEL => mac_control_txfifowerr_cnt_8_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_8_CYINIT,
      I1 => mac_control_txfifowerr_cnt_8_FROM,
      O => mac_control_txfifowerr_cnt_n0000(8)
    );
  mac_control_txfifowerr_cnt_8_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_8_FROM
    );
  mac_control_txfifowerr_cnt_8_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_8_GROM
    );
  mac_control_txfifowerr_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_8_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_25_914 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_8_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_txfifowerr_cnt_8_GROM,
      O => mac_control_txfifowerr_cnt_8_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_txfifowerr_cnt_8_GROM,
      O => mac_control_txfifowerr_cnt_n0000(9)
    );
  mac_control_txfifowerr_cnt_8_CYINIT_915 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_txfifowerr_cnt_8_CYINIT
    );
  mac_control_txfifowerr_cnt_10_LOGIC_ZERO_916 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_10_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_26_917 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_10_CYINIT,
      SEL => mac_control_txfifowerr_cnt_10_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_10_CYINIT,
      I1 => mac_control_txfifowerr_cnt_10_FROM,
      O => mac_control_txfifowerr_cnt_n0000(10)
    );
  mac_control_txfifowerr_cnt_10_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_10_FROM
    );
  mac_control_txfifowerr_cnt_10_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(11),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_10_GROM
    );
  mac_control_txfifowerr_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_10_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_27_918 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_10_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_txfifowerr_cnt_10_GROM,
      O => mac_control_txfifowerr_cnt_10_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_txfifowerr_cnt_10_GROM,
      O => mac_control_txfifowerr_cnt_n0000(11)
    );
  mac_control_txfifowerr_cnt_10_CYINIT_919 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_txfifowerr_cnt_10_CYINIT
    );
  mac_control_txfifowerr_cnt_12_LOGIC_ZERO_920 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_12_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_28_921 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_12_CYINIT,
      SEL => mac_control_txfifowerr_cnt_12_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_12_CYINIT,
      I1 => mac_control_txfifowerr_cnt_12_FROM,
      O => mac_control_txfifowerr_cnt_n0000(12)
    );
  mac_control_txfifowerr_cnt_12_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_12_FROM
    );
  mac_control_txfifowerr_cnt_12_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(13),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_12_GROM
    );
  mac_control_txfifowerr_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_12_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_29_922 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_12_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_txfifowerr_cnt_12_GROM,
      O => mac_control_txfifowerr_cnt_12_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_txfifowerr_cnt_12_GROM,
      O => mac_control_txfifowerr_cnt_n0000(13)
    );
  mac_control_txfifowerr_cnt_12_CYINIT_923 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_txfifowerr_cnt_12_CYINIT
    );
  mac_control_txfifowerr_cnt_14_LOGIC_ZERO_924 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_14_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_30_925 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_14_CYINIT,
      SEL => mac_control_txfifowerr_cnt_14_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_14_CYINIT,
      I1 => mac_control_txfifowerr_cnt_14_FROM,
      O => mac_control_txfifowerr_cnt_n0000(14)
    );
  mac_control_txfifowerr_cnt_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_14_FROM
    );
  mac_control_txfifowerr_cnt_14_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(15),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_14_GROM
    );
  mac_control_txfifowerr_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_14_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_31_926 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_14_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_txfifowerr_cnt_14_GROM,
      O => mac_control_txfifowerr_cnt_14_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_txfifowerr_cnt_14_GROM,
      O => mac_control_txfifowerr_cnt_n0000(15)
    );
  mac_control_txfifowerr_cnt_14_CYINIT_927 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_txfifowerr_cnt_14_CYINIT
    );
  mac_control_txfifowerr_cnt_16_LOGIC_ZERO_928 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_16_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_32_929 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_16_CYINIT,
      SEL => mac_control_txfifowerr_cnt_16_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_16_CYINIT,
      I1 => mac_control_txfifowerr_cnt_16_FROM,
      O => mac_control_txfifowerr_cnt_n0000(16)
    );
  mac_control_txfifowerr_cnt_16_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(16),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_16_FROM
    );
  mac_control_txfifowerr_cnt_16_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(17),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_16_GROM
    );
  mac_control_txfifowerr_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_16_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_33_930 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_16_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_txfifowerr_cnt_16_GROM,
      O => mac_control_txfifowerr_cnt_16_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_txfifowerr_cnt_16_GROM,
      O => mac_control_txfifowerr_cnt_n0000(17)
    );
  mac_control_txfifowerr_cnt_16_CYINIT_931 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_txfifowerr_cnt_16_CYINIT
    );
  mac_control_txfifowerr_cnt_18_LOGIC_ZERO_932 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_18_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_34_933 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_18_CYINIT,
      SEL => mac_control_txfifowerr_cnt_18_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_18_CYINIT,
      I1 => mac_control_txfifowerr_cnt_18_FROM,
      O => mac_control_txfifowerr_cnt_n0000(18)
    );
  mac_control_txfifowerr_cnt_18_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_18_FROM
    );
  mac_control_txfifowerr_cnt_18_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(19),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_18_GROM
    );
  mac_control_txfifowerr_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_18_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_35_934 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_18_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_txfifowerr_cnt_18_GROM,
      O => mac_control_txfifowerr_cnt_18_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_txfifowerr_cnt_18_GROM,
      O => mac_control_txfifowerr_cnt_n0000(19)
    );
  mac_control_txfifowerr_cnt_18_CYINIT_935 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_txfifowerr_cnt_18_CYINIT
    );
  mac_control_txfifowerr_cnt_20_LOGIC_ZERO_936 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_20_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_36_937 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_20_CYINIT,
      SEL => mac_control_txfifowerr_cnt_20_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_20_CYINIT,
      I1 => mac_control_txfifowerr_cnt_20_FROM,
      O => mac_control_txfifowerr_cnt_n0000(20)
    );
  mac_control_txfifowerr_cnt_20_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(20),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_20_FROM
    );
  mac_control_txfifowerr_cnt_20_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(21),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_20_GROM
    );
  mac_control_txfifowerr_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_20_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_37_938 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_20_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_txfifowerr_cnt_20_GROM,
      O => mac_control_txfifowerr_cnt_20_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_txfifowerr_cnt_20_GROM,
      O => mac_control_txfifowerr_cnt_n0000(21)
    );
  mac_control_txfifowerr_cnt_20_CYINIT_939 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_txfifowerr_cnt_20_CYINIT
    );
  mac_control_txfifowerr_cnt_22_LOGIC_ZERO_940 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_22_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_38_941 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_22_CYINIT,
      SEL => mac_control_txfifowerr_cnt_22_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_22_CYINIT,
      I1 => mac_control_txfifowerr_cnt_22_FROM,
      O => mac_control_txfifowerr_cnt_n0000(22)
    );
  mac_control_txfifowerr_cnt_22_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(22),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_22_FROM
    );
  mac_control_txfifowerr_cnt_22_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txfifowerr_cnt(23),
      O => mac_control_txfifowerr_cnt_22_GROM
    );
  mac_control_txfifowerr_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_22_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_39_942 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_22_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_txfifowerr_cnt_22_GROM,
      O => mac_control_txfifowerr_cnt_22_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_txfifowerr_cnt_22_GROM,
      O => mac_control_txfifowerr_cnt_n0000(23)
    );
  mac_control_txfifowerr_cnt_22_CYINIT_943 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_txfifowerr_cnt_22_CYINIT
    );
  mac_control_txfifowerr_cnt_24_LOGIC_ZERO_944 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_24_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_40_945 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_24_CYINIT,
      SEL => mac_control_txfifowerr_cnt_24_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_24_CYINIT,
      I1 => mac_control_txfifowerr_cnt_24_FROM,
      O => mac_control_txfifowerr_cnt_n0000(24)
    );
  mac_control_txfifowerr_cnt_24_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txfifowerr_cnt(24),
      O => mac_control_txfifowerr_cnt_24_FROM
    );
  mac_control_txfifowerr_cnt_24_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(25),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_24_GROM
    );
  mac_control_txfifowerr_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_24_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_41_946 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_24_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_txfifowerr_cnt_24_GROM,
      O => mac_control_txfifowerr_cnt_24_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_txfifowerr_cnt_24_GROM,
      O => mac_control_txfifowerr_cnt_n0000(25)
    );
  mac_control_txfifowerr_cnt_24_CYINIT_947 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_txfifowerr_cnt_24_CYINIT
    );
  mac_control_txfifowerr_cnt_26_LOGIC_ZERO_948 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_26_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_42_949 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_26_CYINIT,
      SEL => mac_control_txfifowerr_cnt_26_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_26_CYINIT,
      I1 => mac_control_txfifowerr_cnt_26_FROM,
      O => mac_control_txfifowerr_cnt_n0000(26)
    );
  mac_control_txfifowerr_cnt_26_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(26),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_26_FROM
    );
  mac_control_txfifowerr_cnt_26_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txfifowerr_cnt(27),
      O => mac_control_txfifowerr_cnt_26_GROM
    );
  mac_control_txfifowerr_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_26_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_43_950 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_26_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_txfifowerr_cnt_26_GROM,
      O => mac_control_txfifowerr_cnt_26_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_txfifowerr_cnt_26_GROM,
      O => mac_control_txfifowerr_cnt_n0000(27)
    );
  mac_control_txfifowerr_cnt_26_CYINIT_951 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_txfifowerr_cnt_26_CYINIT
    );
  mac_control_txfifowerr_cnt_28_LOGIC_ZERO_952 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_28_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_44_953 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_28_CYINIT,
      SEL => mac_control_txfifowerr_cnt_28_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_28_CYINIT,
      I1 => mac_control_txfifowerr_cnt_28_FROM,
      O => mac_control_txfifowerr_cnt_n0000(28)
    );
  mac_control_txfifowerr_cnt_28_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(28),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_28_FROM
    );
  mac_control_txfifowerr_cnt_28_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txfifowerr_cnt(29),
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_28_GROM
    );
  mac_control_txfifowerr_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_28_CYMUXG,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_45_954 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_28_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_txfifowerr_cnt_28_GROM,
      O => mac_control_txfifowerr_cnt_28_CYMUXG
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_txfifowerr_cnt_28_GROM,
      O => mac_control_txfifowerr_cnt_n0000(29)
    );
  mac_control_txfifowerr_cnt_28_CYINIT_955 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_txfifowerr_cnt_28_CYINIT
    );
  mac_control_txfifowerr_cnt_30_LOGIC_ZERO_956 : X_ZERO
    port map (
      O => mac_control_txfifowerr_cnt_30_LOGIC_ZERO
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_46_957 : X_MUX2
    port map (
      IA => mac_control_txfifowerr_cnt_30_LOGIC_ZERO,
      IB => mac_control_txfifowerr_cnt_30_CYINIT,
      SEL => mac_control_txfifowerr_cnt_30_FROM,
      O => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_30_CYINIT,
      I1 => mac_control_txfifowerr_cnt_30_FROM,
      O => mac_control_txfifowerr_cnt_n0000(30)
    );
  mac_control_txfifowerr_cnt_30_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txfifowerr_cnt(30),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_30_FROM
    );
  mac_control_txfifowerr_cnt_31_rt_958 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cnt(31),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txfifowerr_cnt_31_rt
    );
  mac_control_txfifowerr_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_txfifowerr_cnt_31_rt,
      O => mac_control_txfifowerr_cnt_n0000(31)
    );
  mac_control_txfifowerr_cnt_30_CYINIT_959 : X_BUF
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_txfifowerr_cnt_30_CYINIT
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ONE_960 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ZERO_961 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_177_962 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(25),
      ADR1 => rx_input_memio_addrchk_macaddrl(24),
      ADR2 => rx_input_memio_addrchk_datal(24),
      ADR3 => rx_input_memio_addrchk_datal(25),
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(27),
      ADR1 => rx_input_memio_addrchk_macaddrl(27),
      ADR2 => rx_input_memio_addrchk_macaddrl(26),
      ADR3 => rx_input_memio_addrchk_datal(26),
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_963 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_2_LOGIC_ZERO_964 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_2_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_179_965 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_2_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_2_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(29),
      ADR1 => rx_input_memio_addrchk_datal(28),
      ADR2 => rx_input_memio_addrchk_macaddrl(28),
      ADR3 => rx_input_memio_addrchk_datal(29),
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(30),
      ADR1 => rx_input_memio_addrchk_datal(31),
      ADR2 => rx_input_memio_addrchk_macaddrl(31),
      ADR3 => rx_input_memio_addrchk_datal(30),
      O => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_2_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_2_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(2)
    );
  rx_input_memio_addrchk_Mcompar_n0042_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_2_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0042_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_2_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_2_CYINIT_966 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0042_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_2_CYINIT
    );
  rx_output_bp_0_LOGIC_ONE_967 : X_ONE
    port map (
      O => rx_output_bp_0_LOGIC_ONE
    );
  rx_output_Madd_lbp_inst_cy_86_968 : X_MUX2
    port map (
      IA => rx_output_lenr(2),
      IB => rx_output_bp_0_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_79,
      O => rx_output_Madd_lbp_inst_cy_86
    );
  rx_output_Madd_lbp_inst_sum_79 : X_XOR2
    port map (
      I0 => rx_output_bp_0_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_79,
      O => rx_output_lbp(0)
    );
  rx_output_Madd_lbp_inst_lut2_791 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_lenr(2),
      ADR1 => VCC,
      ADR2 => rx_output_bp(0),
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_79
    );
  rx_output_Madd_lbp_inst_lut2_801 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(1),
      O => rx_output_Madd_lbp_inst_lut2_80
    );
  rx_output_bp_0_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_0_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_87
    );
  rx_output_Madd_lbp_inst_cy_87_969 : X_MUX2
    port map (
      IA => rx_output_lenr(3),
      IB => rx_output_Madd_lbp_inst_cy_86,
      SEL => rx_output_Madd_lbp_inst_lut2_80,
      O => rx_output_bp_0_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_80 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_86,
      I1 => rx_output_Madd_lbp_inst_lut2_80,
      O => rx_output_lbp(1)
    );
  rx_output_bp_0_CYINIT_970 : X_BUF
    port map (
      I => rx_output_bp_0_LOGIC_ONE,
      O => rx_output_bp_0_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_88_971 : X_MUX2
    port map (
      IA => rx_output_lenr(4),
      IB => rx_output_bp_2_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_81,
      O => rx_output_Madd_lbp_inst_cy_88
    );
  rx_output_Madd_lbp_inst_sum_81 : X_XOR2
    port map (
      I0 => rx_output_bp_2_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_81,
      O => rx_output_lbp(2)
    );
  rx_output_Madd_lbp_inst_lut2_811 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(2),
      O => rx_output_Madd_lbp_inst_lut2_81
    );
  rx_output_Madd_lbp_inst_lut2_821 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_lenr(5),
      ADR1 => VCC,
      ADR2 => rx_output_bp(3),
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_82
    );
  rx_output_bp_2_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_2_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_89
    );
  rx_output_Madd_lbp_inst_cy_89_972 : X_MUX2
    port map (
      IA => rx_output_lenr(5),
      IB => rx_output_Madd_lbp_inst_cy_88,
      SEL => rx_output_Madd_lbp_inst_lut2_82,
      O => rx_output_bp_2_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_82 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_88,
      I1 => rx_output_Madd_lbp_inst_lut2_82,
      O => rx_output_lbp(3)
    );
  rx_output_bp_2_CYINIT_973 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_87,
      O => rx_output_bp_2_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_90_974 : X_MUX2
    port map (
      IA => rx_output_lenr(6),
      IB => rx_output_bp_4_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_83,
      O => rx_output_Madd_lbp_inst_cy_90
    );
  rx_output_Madd_lbp_inst_sum_83 : X_XOR2
    port map (
      I0 => rx_output_bp_4_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_83,
      O => rx_output_lbp(4)
    );
  rx_output_Madd_lbp_inst_lut2_831 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_lenr(6),
      ADR1 => VCC,
      ADR2 => rx_output_bp(4),
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_83
    );
  rx_output_Madd_lbp_inst_lut2_841 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(7),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(5),
      O => rx_output_Madd_lbp_inst_lut2_84
    );
  rx_output_bp_4_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_4_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_91
    );
  rx_output_Madd_lbp_inst_cy_91_975 : X_MUX2
    port map (
      IA => rx_output_lenr(7),
      IB => rx_output_Madd_lbp_inst_cy_90,
      SEL => rx_output_Madd_lbp_inst_lut2_84,
      O => rx_output_bp_4_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_84 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_90,
      I1 => rx_output_Madd_lbp_inst_lut2_84,
      O => rx_output_lbp(5)
    );
  rx_output_bp_4_CYINIT_976 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_89,
      O => rx_output_bp_4_CYINIT
    );
  rx_input_fifo_control_DATA_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(1),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_1_FFY_RST,
      O => rx_input_data(1)
    );
  rx_input_data_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_1_FFY_RST
    );
  rx_output_Madd_lbp_inst_cy_92_977 : X_MUX2
    port map (
      IA => rx_output_lenr(8),
      IB => rx_output_bp_6_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_85,
      O => rx_output_Madd_lbp_inst_cy_92
    );
  rx_output_Madd_lbp_inst_sum_85 : X_XOR2
    port map (
      I0 => rx_output_bp_6_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_85,
      O => rx_output_lbp(6)
    );
  rx_output_Madd_lbp_inst_lut2_851 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(6),
      O => rx_output_Madd_lbp_inst_lut2_85
    );
  rx_output_Madd_lbp_inst_lut2_861 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(7),
      O => rx_output_Madd_lbp_inst_lut2_86
    );
  rx_output_bp_6_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_6_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_93
    );
  rx_output_Madd_lbp_inst_cy_93_978 : X_MUX2
    port map (
      IA => rx_output_lenr(9),
      IB => rx_output_Madd_lbp_inst_cy_92,
      SEL => rx_output_Madd_lbp_inst_lut2_86,
      O => rx_output_bp_6_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_86 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_92,
      I1 => rx_output_Madd_lbp_inst_lut2_86,
      O => rx_output_lbp(7)
    );
  rx_output_bp_6_CYINIT_979 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_91,
      O => rx_output_bp_6_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_94_980 : X_MUX2
    port map (
      IA => rx_output_lenr(10),
      IB => rx_output_bp_8_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_87,
      O => rx_output_Madd_lbp_inst_cy_94
    );
  rx_output_Madd_lbp_inst_sum_87 : X_XOR2
    port map (
      I0 => rx_output_bp_8_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_87,
      O => rx_output_lbp(8)
    );
  rx_output_Madd_lbp_inst_lut2_871 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_lenr(10),
      ADR1 => rx_output_bp(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_87
    );
  rx_output_Madd_lbp_inst_lut2_881 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_lenr(11),
      ADR1 => VCC,
      ADR2 => rx_output_bp(9),
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_88
    );
  rx_output_bp_8_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_8_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_95
    );
  rx_output_Madd_lbp_inst_cy_95_981 : X_MUX2
    port map (
      IA => rx_output_lenr(11),
      IB => rx_output_Madd_lbp_inst_cy_94,
      SEL => rx_output_Madd_lbp_inst_lut2_88,
      O => rx_output_bp_8_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_88 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_94,
      I1 => rx_output_Madd_lbp_inst_lut2_88,
      O => rx_output_lbp(9)
    );
  rx_output_bp_8_CYINIT_982 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_93,
      O => rx_output_bp_8_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_96_983 : X_MUX2
    port map (
      IA => rx_output_lenr(12),
      IB => rx_output_bp_10_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_89,
      O => rx_output_Madd_lbp_inst_cy_96
    );
  rx_output_Madd_lbp_inst_sum_89 : X_XOR2
    port map (
      I0 => rx_output_bp_10_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_89,
      O => rx_output_lbp(10)
    );
  rx_output_Madd_lbp_inst_lut2_891 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rx_output_lenr(12),
      ADR1 => VCC,
      ADR2 => rx_output_bp(10),
      ADR3 => VCC,
      O => rx_output_Madd_lbp_inst_lut2_89
    );
  rx_output_Madd_lbp_inst_lut2_901 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(11),
      O => rx_output_Madd_lbp_inst_lut2_90
    );
  rx_output_bp_10_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_10_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_97
    );
  rx_output_Madd_lbp_inst_cy_97_984 : X_MUX2
    port map (
      IA => rx_output_lenr(13),
      IB => rx_output_Madd_lbp_inst_cy_96,
      SEL => rx_output_Madd_lbp_inst_lut2_90,
      O => rx_output_bp_10_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_90 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_96,
      I1 => rx_output_Madd_lbp_inst_lut2_90,
      O => rx_output_lbp(11)
    );
  rx_output_bp_10_CYINIT_985 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_95,
      O => rx_output_bp_10_CYINIT
    );
  rx_output_Madd_lbp_inst_cy_98_986 : X_MUX2
    port map (
      IA => rx_output_lenr(14),
      IB => rx_output_bp_12_CYINIT,
      SEL => rx_output_Madd_lbp_inst_lut2_91,
      O => rx_output_Madd_lbp_inst_cy_98
    );
  rx_output_Madd_lbp_inst_sum_91 : X_XOR2
    port map (
      I0 => rx_output_bp_12_CYINIT,
      I1 => rx_output_Madd_lbp_inst_lut2_91,
      O => rx_output_lbp(12)
    );
  rx_output_Madd_lbp_inst_lut2_911 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(14),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(12),
      O => rx_output_Madd_lbp_inst_lut2_91
    );
  rx_output_Madd_lbp_inst_lut2_921 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_lenr(15),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(13),
      O => rx_output_Madd_lbp_inst_lut2_92
    );
  rx_output_bp_12_COUTUSED : X_BUF
    port map (
      I => rx_output_bp_12_CYMUXG,
      O => rx_output_Madd_lbp_inst_cy_99
    );
  rx_output_Madd_lbp_inst_cy_99_987 : X_MUX2
    port map (
      IA => rx_output_lenr(15),
      IB => rx_output_Madd_lbp_inst_cy_98,
      SEL => rx_output_Madd_lbp_inst_lut2_92,
      O => rx_output_bp_12_CYMUXG
    );
  rx_output_Madd_lbp_inst_sum_92 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_98,
      I1 => rx_output_Madd_lbp_inst_lut2_92,
      O => rx_output_lbp(13)
    );
  rx_output_bp_12_CYINIT_988 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_97,
      O => rx_output_bp_12_CYINIT
    );
  rx_output_bp_14_LOGIC_ZERO_989 : X_ZERO
    port map (
      O => rx_output_bp_14_LOGIC_ZERO
    );
  rx_output_Madd_lbp_inst_cy_100_990 : X_MUX2
    port map (
      IA => rx_output_bp_14_LOGIC_ZERO,
      IB => rx_output_bp_14_CYINIT,
      SEL => rx_output_bp_14_FROM,
      O => rx_output_Madd_lbp_inst_cy_100
    );
  rx_output_Madd_lbp_inst_sum_93 : X_XOR2
    port map (
      I0 => rx_output_bp_14_CYINIT,
      I1 => rx_output_bp_14_FROM,
      O => rx_output_lbp(14)
    );
  rx_output_bp_14_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_bp(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_bp_14_FROM
    );
  rx_output_bp_15_rt_991 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_bp(15),
      O => rx_output_bp_15_rt
    );
  rx_output_Madd_lbp_inst_sum_94 : X_XOR2
    port map (
      I0 => rx_output_Madd_lbp_inst_cy_100,
      I1 => rx_output_bp_15_rt,
      O => rx_output_lbp(15)
    );
  rx_output_bp_14_CYINIT_992 : X_BUF
    port map (
      I => rx_output_Madd_lbp_inst_cy_99,
      O => rx_output_bp_14_CYINIT
    );
  tx_output_bcnt_38_LOGIC_ONE_993 : X_ONE
    port map (
      O => tx_output_bcnt_38_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_204_994 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_17,
      IB => tx_output_bcnt_38_LOGIC_ONE,
      SEL => tx_output_cs_FFd12_rt,
      O => tx_output_bcnt_inst_cy_204
    );
  tx_output_cs_FFd12_rt_995 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_17,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd12,
      ADR3 => VCC,
      O => tx_output_cs_FFd12_rt
    );
  tx_output_bcnt_inst_lut3_401 : X_LUT4
    generic map(
      INIT => X"03CF"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_10,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_bcnt_38,
      ADR3 => q2(0),
      O => tx_output_bcnt_inst_lut3_40
    );
  tx_output_bcnt_38_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_38_CYMUXG,
      O => tx_output_bcnt_inst_cy_205
    );
  tx_output_bcnt_inst_cy_205_996 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_10,
      IB => tx_output_bcnt_inst_cy_204,
      SEL => tx_output_bcnt_inst_lut3_40,
      O => tx_output_bcnt_38_CYMUXG
    );
  tx_output_bcnt_inst_sum_171_997 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_204,
      I1 => tx_output_bcnt_inst_lut3_40,
      O => tx_output_bcnt_inst_sum_171
    );
  tx_output_bcnt_39_LOGIC_ONE_998 : X_ONE
    port map (
      O => tx_output_bcnt_39_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_206_999 : X_MUX2
    port map (
      IA => tx_output_bcnt_39_LOGIC_ONE,
      IB => tx_output_bcnt_39_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_41,
      O => tx_output_bcnt_inst_cy_206
    );
  tx_output_bcnt_inst_sum_172_1000 : X_XOR2
    port map (
      I0 => tx_output_bcnt_39_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_41,
      O => tx_output_bcnt_inst_sum_172
    );
  tx_output_bcnt_inst_lut3_411 : X_LUT4
    generic map(
      INIT => X"4747"
    )
    port map (
      ADR0 => q2(1),
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_bcnt_39,
      ADR3 => VCC,
      O => tx_output_bcnt_inst_lut3_41
    );
  tx_output_bcnt_inst_lut3_421 : X_LUT4
    generic map(
      INIT => X"03CF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_bcnt_40,
      ADR3 => q2(2),
      O => tx_output_bcnt_inst_lut3_42
    );
  tx_output_bcnt_39_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_39_CYMUXG,
      O => tx_output_bcnt_inst_cy_207
    );
  tx_output_bcnt_inst_cy_207_1001 : X_MUX2
    port map (
      IA => tx_output_bcnt_39_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_206,
      SEL => tx_output_bcnt_inst_lut3_42,
      O => tx_output_bcnt_39_CYMUXG
    );
  tx_output_bcnt_inst_sum_173_1002 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_206,
      I1 => tx_output_bcnt_inst_lut3_42,
      O => tx_output_bcnt_inst_sum_173
    );
  tx_output_bcnt_39_CYINIT_1003 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_205,
      O => tx_output_bcnt_39_CYINIT
    );
  tx_output_bcnt_41_LOGIC_ONE_1004 : X_ONE
    port map (
      O => tx_output_bcnt_41_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_208_1005 : X_MUX2
    port map (
      IA => tx_output_bcnt_41_LOGIC_ONE,
      IB => tx_output_bcnt_41_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_43,
      O => tx_output_bcnt_inst_cy_208
    );
  tx_output_bcnt_inst_sum_174_1006 : X_XOR2
    port map (
      I0 => tx_output_bcnt_41_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_43,
      O => tx_output_bcnt_inst_sum_174
    );
  tx_output_bcnt_inst_lut3_431 : X_LUT4
    generic map(
      INIT => X"4747"
    )
    port map (
      ADR0 => q2(3),
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_bcnt_41,
      ADR3 => VCC,
      O => tx_output_bcnt_inst_lut3_43
    );
  tx_output_bcnt_inst_lut3_441 : X_LUT4
    generic map(
      INIT => X"03CF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_bcnt_42,
      ADR3 => q2(4),
      O => tx_output_bcnt_inst_lut3_44
    );
  tx_output_bcnt_41_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_41_CYMUXG,
      O => tx_output_bcnt_inst_cy_209
    );
  tx_output_bcnt_inst_cy_209_1007 : X_MUX2
    port map (
      IA => tx_output_bcnt_41_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_208,
      SEL => tx_output_bcnt_inst_lut3_44,
      O => tx_output_bcnt_41_CYMUXG
    );
  tx_output_bcnt_inst_sum_175_1008 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_208,
      I1 => tx_output_bcnt_inst_lut3_44,
      O => tx_output_bcnt_inst_sum_175
    );
  tx_output_bcnt_41_CYINIT_1009 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_207,
      O => tx_output_bcnt_41_CYINIT
    );
  tx_output_bcnt_43_LOGIC_ONE_1010 : X_ONE
    port map (
      O => tx_output_bcnt_43_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_210_1011 : X_MUX2
    port map (
      IA => tx_output_bcnt_43_LOGIC_ONE,
      IB => tx_output_bcnt_43_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_45,
      O => tx_output_bcnt_inst_cy_210
    );
  tx_output_bcnt_inst_sum_176_1012 : X_XOR2
    port map (
      I0 => tx_output_bcnt_43_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_45,
      O => tx_output_bcnt_inst_sum_176
    );
  tx_output_bcnt_inst_lut3_451 : X_LUT4
    generic map(
      INIT => X"4747"
    )
    port map (
      ADR0 => q2(5),
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_bcnt_43,
      ADR3 => VCC,
      O => tx_output_bcnt_inst_lut3_45
    );
  tx_output_bcnt_inst_lut3_461 : X_LUT4
    generic map(
      INIT => X"0F33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_bcnt_44,
      ADR2 => q2(6),
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_46
    );
  tx_output_bcnt_43_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_43_CYMUXG,
      O => tx_output_bcnt_inst_cy_211
    );
  tx_output_bcnt_inst_cy_211_1013 : X_MUX2
    port map (
      IA => tx_output_bcnt_43_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_210,
      SEL => tx_output_bcnt_inst_lut3_46,
      O => tx_output_bcnt_43_CYMUXG
    );
  tx_output_bcnt_inst_sum_177_1014 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_210,
      I1 => tx_output_bcnt_inst_lut3_46,
      O => tx_output_bcnt_inst_sum_177
    );
  tx_output_bcnt_43_CYINIT_1015 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_209,
      O => tx_output_bcnt_43_CYINIT
    );
  tx_output_bcnt_45_LOGIC_ONE_1016 : X_ONE
    port map (
      O => tx_output_bcnt_45_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_212_1017 : X_MUX2
    port map (
      IA => tx_output_bcnt_45_LOGIC_ONE,
      IB => tx_output_bcnt_45_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_47,
      O => tx_output_bcnt_inst_cy_212
    );
  tx_output_bcnt_inst_sum_178_1018 : X_XOR2
    port map (
      I0 => tx_output_bcnt_45_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_47,
      O => tx_output_bcnt_inst_sum_178
    );
  tx_output_bcnt_inst_lut3_471 : X_LUT4
    generic map(
      INIT => X"550F"
    )
    port map (
      ADR0 => q2(7),
      ADR1 => VCC,
      ADR2 => tx_output_bcnt_45,
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_47
    );
  tx_output_bcnt_inst_lut3_481 : X_LUT4
    generic map(
      INIT => X"4747"
    )
    port map (
      ADR0 => q2(8),
      ADR1 => tx_output_cs_FFd12,
      ADR2 => tx_output_bcnt_46,
      ADR3 => VCC,
      O => tx_output_bcnt_inst_lut3_48
    );
  tx_output_bcnt_45_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_45_CYMUXG,
      O => tx_output_bcnt_inst_cy_213
    );
  tx_output_bcnt_inst_cy_213_1019 : X_MUX2
    port map (
      IA => tx_output_bcnt_45_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_212,
      SEL => tx_output_bcnt_inst_lut3_48,
      O => tx_output_bcnt_45_CYMUXG
    );
  tx_output_bcnt_inst_sum_179_1020 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_212,
      I1 => tx_output_bcnt_inst_lut3_48,
      O => tx_output_bcnt_inst_sum_179
    );
  tx_output_bcnt_45_CYINIT_1021 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_211,
      O => tx_output_bcnt_45_CYINIT
    );
  tx_output_bcnt_47_LOGIC_ONE_1022 : X_ONE
    port map (
      O => tx_output_bcnt_47_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_214_1023 : X_MUX2
    port map (
      IA => tx_output_bcnt_47_LOGIC_ONE,
      IB => tx_output_bcnt_47_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_49,
      O => tx_output_bcnt_inst_cy_214
    );
  tx_output_bcnt_inst_sum_180_1024 : X_XOR2
    port map (
      I0 => tx_output_bcnt_47_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_49,
      O => tx_output_bcnt_inst_sum_180
    );
  tx_output_bcnt_inst_lut3_491 : X_LUT4
    generic map(
      INIT => X"550F"
    )
    port map (
      ADR0 => q2(9),
      ADR1 => VCC,
      ADR2 => tx_output_bcnt_47,
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_49
    );
  tx_output_bcnt_inst_lut3_501 : X_LUT4
    generic map(
      INIT => X"0C3F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => q2(10),
      ADR3 => tx_output_bcnt_48,
      O => tx_output_bcnt_inst_lut3_50
    );
  tx_output_bcnt_47_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_47_CYMUXG,
      O => tx_output_bcnt_inst_cy_215
    );
  tx_output_bcnt_inst_cy_215_1025 : X_MUX2
    port map (
      IA => tx_output_bcnt_47_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_214,
      SEL => tx_output_bcnt_inst_lut3_50,
      O => tx_output_bcnt_47_CYMUXG
    );
  tx_output_bcnt_inst_sum_181_1026 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_214,
      I1 => tx_output_bcnt_inst_lut3_50,
      O => tx_output_bcnt_inst_sum_181
    );
  tx_output_bcnt_47_CYINIT_1027 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_213,
      O => tx_output_bcnt_47_CYINIT
    );
  tx_output_bcnt_49_LOGIC_ONE_1028 : X_ONE
    port map (
      O => tx_output_bcnt_49_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_216_1029 : X_MUX2
    port map (
      IA => tx_output_bcnt_49_LOGIC_ONE,
      IB => tx_output_bcnt_49_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_51,
      O => tx_output_bcnt_inst_cy_216
    );
  tx_output_bcnt_inst_sum_182_1030 : X_XOR2
    port map (
      I0 => tx_output_bcnt_49_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_51,
      O => tx_output_bcnt_inst_sum_182
    );
  tx_output_bcnt_inst_lut3_511 : X_LUT4
    generic map(
      INIT => X"0F33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_bcnt_49,
      ADR2 => q2(11),
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_51
    );
  tx_output_bcnt_inst_lut3_521 : X_LUT4
    generic map(
      INIT => X"0F55"
    )
    port map (
      ADR0 => tx_output_bcnt_50,
      ADR1 => VCC,
      ADR2 => q2(12),
      ADR3 => tx_output_cs_FFd12,
      O => tx_output_bcnt_inst_lut3_52
    );
  tx_output_bcnt_49_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_49_CYMUXG,
      O => tx_output_bcnt_inst_cy_217
    );
  tx_output_bcnt_inst_cy_217_1031 : X_MUX2
    port map (
      IA => tx_output_bcnt_49_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_216,
      SEL => tx_output_bcnt_inst_lut3_52,
      O => tx_output_bcnt_49_CYMUXG
    );
  tx_output_bcnt_inst_sum_183_1032 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_216,
      I1 => tx_output_bcnt_inst_lut3_52,
      O => tx_output_bcnt_inst_sum_183
    );
  tx_output_bcnt_49_CYINIT_1033 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_215,
      O => tx_output_bcnt_49_CYINIT
    );
  tx_output_bcnt_51_LOGIC_ONE_1034 : X_ONE
    port map (
      O => tx_output_bcnt_51_LOGIC_ONE
    );
  tx_output_bcnt_inst_cy_218_1035 : X_MUX2
    port map (
      IA => tx_output_bcnt_51_LOGIC_ONE,
      IB => tx_output_bcnt_51_CYINIT,
      SEL => tx_output_bcnt_inst_lut3_53,
      O => tx_output_bcnt_inst_cy_218
    );
  tx_output_bcnt_inst_sum_184_1036 : X_XOR2
    port map (
      I0 => tx_output_bcnt_51_CYINIT,
      I1 => tx_output_bcnt_inst_lut3_53,
      O => tx_output_bcnt_inst_sum_184
    );
  tx_output_bcnt_inst_lut3_531 : X_LUT4
    generic map(
      INIT => X"2727"
    )
    port map (
      ADR0 => tx_output_cs_FFd12,
      ADR1 => q2(13),
      ADR2 => tx_output_bcnt_51,
      ADR3 => VCC,
      O => tx_output_bcnt_inst_lut3_53
    );
  tx_output_bcnt_inst_lut3_541 : X_LUT4
    generic map(
      INIT => X"05F5"
    )
    port map (
      ADR0 => tx_output_bcnt_52,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd12,
      ADR3 => q2(14),
      O => tx_output_bcnt_inst_lut3_54
    );
  tx_output_bcnt_51_COUTUSED : X_BUF
    port map (
      I => tx_output_bcnt_51_CYMUXG,
      O => tx_output_bcnt_inst_cy_219
    );
  tx_output_bcnt_inst_cy_219_1037 : X_MUX2
    port map (
      IA => tx_output_bcnt_51_LOGIC_ONE,
      IB => tx_output_bcnt_inst_cy_218,
      SEL => tx_output_bcnt_inst_lut3_54,
      O => tx_output_bcnt_51_CYMUXG
    );
  tx_output_bcnt_inst_sum_185_1038 : X_XOR2
    port map (
      I0 => tx_output_bcnt_inst_cy_218,
      I1 => tx_output_bcnt_inst_lut3_54,
      O => tx_output_bcnt_inst_sum_185
    );
  tx_output_bcnt_51_CYINIT_1039 : X_BUF
    port map (
      I => tx_output_bcnt_inst_cy_217,
      O => tx_output_bcnt_51_CYINIT
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ONE_1040 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ZERO_1041 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_177_1042 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(17),
      ADR1 => rx_input_memio_addrchk_macaddrl(16),
      ADR2 => rx_input_memio_addrchk_macaddrl(17),
      ADR3 => rx_input_memio_addrchk_datal(16),
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(19),
      ADR1 => rx_input_memio_addrchk_macaddrl(18),
      ADR2 => rx_input_memio_addrchk_macaddrl(19),
      ADR3 => rx_input_memio_addrchk_datal(18),
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_1043 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_3_LOGIC_ZERO_1044 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_3_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_179_1045 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_3_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_3_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(21),
      ADR1 => rx_input_memio_addrchk_macaddrl(21),
      ADR2 => rx_input_memio_addrchk_datal(20),
      ADR3 => rx_input_memio_addrchk_macaddrl(20),
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(22),
      ADR1 => rx_input_memio_addrchk_macaddrl(22),
      ADR2 => rx_input_memio_addrchk_macaddrl(23),
      ADR3 => rx_input_memio_addrchk_datal(23),
      O => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_3_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_3_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(3)
    );
  rx_input_memio_addrchk_Mcompar_n0039_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_3_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0039_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_3_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_3_CYINIT_1046 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0039_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_3_CYINIT
    );
  rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ONE_1047 : X_ONE
    port map (
      O => rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ONE
    );
  rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ZERO_1048 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ZERO
    );
  rx_output_Mcompar_n0017_inst_cy_78_1049 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ONE,
      SEL => rx_output_Mcompar_n0017_inst_lut4_0,
      O => rx_output_Mcompar_n0017_inst_cy_78
    );
  rx_output_Mcompar_n0017_inst_lut4_01 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rxfbbp(0),
      ADR1 => rxfbbp(1),
      ADR2 => rxbp(0),
      ADR3 => rxbp(1),
      O => rx_output_Mcompar_n0017_inst_lut4_0
    );
  rx_output_Mcompar_n0017_inst_lut4_11 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rxfbbp(3),
      ADR1 => rxbp(3),
      ADR2 => rxfbbp(2),
      ADR3 => rxbp(2),
      O => rx_output_Mcompar_n0017_inst_lut4_1
    );
  rx_output_Mcompar_n0017_inst_cy_79_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_79_CYMUXG,
      O => rx_output_Mcompar_n0017_inst_cy_79
    );
  rx_output_Mcompar_n0017_inst_cy_79_1050 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_79_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_78,
      SEL => rx_output_Mcompar_n0017_inst_lut4_1,
      O => rx_output_Mcompar_n0017_inst_cy_79_CYMUXG
    );
  rx_output_Mcompar_n0017_inst_cy_81_LOGIC_ZERO_1051 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0017_inst_cy_81_LOGIC_ZERO
    );
  rx_output_Mcompar_n0017_inst_cy_80_1052 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_81_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_81_CYINIT,
      SEL => rx_output_Mcompar_n0017_inst_lut4_2,
      O => rx_output_Mcompar_n0017_inst_cy_80
    );
  rx_output_Mcompar_n0017_inst_lut4_21 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rxbp(5),
      ADR1 => rxfbbp(5),
      ADR2 => rxbp(4),
      ADR3 => rxfbbp(4),
      O => rx_output_Mcompar_n0017_inst_lut4_2
    );
  rx_output_Mcompar_n0017_inst_lut4_31 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rxbp(6),
      ADR1 => rxbp(7),
      ADR2 => rxfbbp(7),
      ADR3 => rxfbbp(6),
      O => rx_output_Mcompar_n0017_inst_lut4_3
    );
  rx_output_Mcompar_n0017_inst_cy_81_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_81_CYMUXG,
      O => rx_output_Mcompar_n0017_inst_cy_81
    );
  rx_output_Mcompar_n0017_inst_cy_81_1053 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_81_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_80,
      SEL => rx_output_Mcompar_n0017_inst_lut4_3,
      O => rx_output_Mcompar_n0017_inst_cy_81_CYMUXG
    );
  rx_output_Mcompar_n0017_inst_cy_81_CYINIT_1054 : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_79,
      O => rx_output_Mcompar_n0017_inst_cy_81_CYINIT
    );
  rx_input_fifo_control_DATA_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(2),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_2_FFY_RST,
      O => rx_input_data(2)
    );
  rx_input_data_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_2_FFY_RST
    );
  rx_output_Mcompar_n0017_inst_cy_83_LOGIC_ZERO_1055 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0017_inst_cy_83_LOGIC_ZERO
    );
  rx_output_Mcompar_n0017_inst_cy_82_1056 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_83_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_83_CYINIT,
      SEL => rx_output_Mcompar_n0017_inst_lut4_4,
      O => rx_output_Mcompar_n0017_inst_cy_82
    );
  rx_output_Mcompar_n0017_inst_lut4_41 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rxbp(9),
      ADR1 => rxfbbp(8),
      ADR2 => rxfbbp(9),
      ADR3 => rxbp(8),
      O => rx_output_Mcompar_n0017_inst_lut4_4
    );
  rx_output_Mcompar_n0017_inst_lut4_51 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rxbp(11),
      ADR1 => rxfbbp(11),
      ADR2 => rxbp(10),
      ADR3 => rxfbbp(10),
      O => rx_output_Mcompar_n0017_inst_lut4_5
    );
  rx_output_Mcompar_n0017_inst_cy_83_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_83_CYMUXG,
      O => rx_output_Mcompar_n0017_inst_cy_83
    );
  rx_output_Mcompar_n0017_inst_cy_83_1057 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0017_inst_cy_83_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_82,
      SEL => rx_output_Mcompar_n0017_inst_lut4_5,
      O => rx_output_Mcompar_n0017_inst_cy_83_CYMUXG
    );
  rx_output_Mcompar_n0017_inst_cy_83_CYINIT_1058 : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_81,
      O => rx_output_Mcompar_n0017_inst_cy_83_CYINIT
    );
  rx_output_n0017_LOGIC_ZERO_1059 : X_ZERO
    port map (
      O => rx_output_n0017_LOGIC_ZERO
    );
  rx_output_Mcompar_n0017_inst_cy_84_1060 : X_MUX2
    port map (
      IA => rx_output_n0017_LOGIC_ZERO,
      IB => rx_output_n0017_CYINIT,
      SEL => rx_output_Mcompar_n0017_inst_lut4_6,
      O => rx_output_Mcompar_n0017_inst_cy_84
    );
  rx_output_Mcompar_n0017_inst_lut4_61 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rxfbbp(12),
      ADR1 => rxbp(12),
      ADR2 => rxbp(13),
      ADR3 => rxfbbp(13),
      O => rx_output_Mcompar_n0017_inst_lut4_6
    );
  rx_output_Mcompar_n0017_inst_lut4_71 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rxbp(15),
      ADR1 => rxbp(14),
      ADR2 => rxfbbp(14),
      ADR3 => rxfbbp(15),
      O => rx_output_Mcompar_n0017_inst_lut4_7
    );
  rx_output_n0017_COUTUSED : X_BUF
    port map (
      I => rx_output_n0017_CYMUXG,
      O => rx_output_n0017
    );
  rx_output_Mcompar_n0017_inst_cy_85 : X_MUX2
    port map (
      IA => rx_output_n0017_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0017_inst_cy_84,
      SEL => rx_output_Mcompar_n0017_inst_lut4_7,
      O => rx_output_n0017_CYMUXG
    );
  rx_output_n0017_CYINIT_1061 : X_BUF
    port map (
      I => rx_output_Mcompar_n0017_inst_cy_83,
      O => rx_output_n0017_CYINIT
    );
  rx_fifocheck_diff_0_LOGIC_ONE_1062 : X_ONE
    port map (
      O => rx_fifocheck_diff_0_LOGIC_ONE
    );
  rx_fifocheck_Msub_n0001_inst_cy_161_1063 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(0),
      IB => rx_fifocheck_diff_0_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_111,
      O => rx_fifocheck_Msub_n0001_inst_cy_161
    );
  rx_fifocheck_Msub_n0001_inst_sum_143 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_0_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_111,
      O => rx_fifocheck_n0001(0)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1111 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(0),
      ADR1 => rx_fifocheck_bpl(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_111
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1121 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(1),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(1),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_112
    );
  rx_fifocheck_diff_0_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_0_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_162
    );
  rx_fifocheck_Msub_n0001_inst_cy_162_1064 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(1),
      IB => rx_fifocheck_Msub_n0001_inst_cy_161,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_112,
      O => rx_fifocheck_diff_0_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_144 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_161,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_112,
      O => rx_fifocheck_n0001(1)
    );
  rx_fifocheck_diff_0_CYINIT_1065 : X_BUF
    port map (
      I => rx_fifocheck_diff_0_LOGIC_ONE,
      O => rx_fifocheck_diff_0_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_163_1066 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(2),
      IB => rx_fifocheck_diff_2_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_113,
      O => rx_fifocheck_Msub_n0001_inst_cy_163
    );
  rx_fifocheck_Msub_n0001_inst_sum_145 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_2_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_113,
      O => rx_fifocheck_n0001(2)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1131 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_bpl(2),
      O => rx_fifocheck_Msub_n0001_inst_lut2_113
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1141 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_bpl(3),
      O => rx_fifocheck_Msub_n0001_inst_lut2_114
    );
  rx_fifocheck_diff_2_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_2_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_164
    );
  rx_fifocheck_Msub_n0001_inst_cy_164_1067 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(3),
      IB => rx_fifocheck_Msub_n0001_inst_cy_163,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_114,
      O => rx_fifocheck_diff_2_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_146 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_163,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_114,
      O => rx_fifocheck_n0001(3)
    );
  rx_fifocheck_diff_2_CYINIT_1068 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_162,
      O => rx_fifocheck_diff_2_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_165_1069 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(4),
      IB => rx_fifocheck_diff_4_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_115,
      O => rx_fifocheck_Msub_n0001_inst_cy_165
    );
  rx_fifocheck_Msub_n0001_inst_sum_147 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_4_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_115,
      O => rx_fifocheck_n0001(4)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1151 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_bpl(4),
      O => rx_fifocheck_Msub_n0001_inst_lut2_115
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1161 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(5),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(5),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_116
    );
  rx_fifocheck_diff_4_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_4_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_166
    );
  rx_fifocheck_Msub_n0001_inst_cy_166_1070 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(5),
      IB => rx_fifocheck_Msub_n0001_inst_cy_165,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_116,
      O => rx_fifocheck_diff_4_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_148 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_165,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_116,
      O => rx_fifocheck_n0001(5)
    );
  rx_fifocheck_diff_4_CYINIT_1071 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_164,
      O => rx_fifocheck_diff_4_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_167_1072 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(6),
      IB => rx_fifocheck_diff_6_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_117,
      O => rx_fifocheck_Msub_n0001_inst_cy_167
    );
  rx_fifocheck_Msub_n0001_inst_sum_149 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_6_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_117,
      O => rx_fifocheck_n0001(6)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1171 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(6),
      ADR1 => rx_fifocheck_bpl(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_117
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1181 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(7),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(7),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_118
    );
  rx_fifocheck_diff_6_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_6_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_168
    );
  rx_fifocheck_Msub_n0001_inst_cy_168_1073 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(7),
      IB => rx_fifocheck_Msub_n0001_inst_cy_167,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_118,
      O => rx_fifocheck_diff_6_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_150 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_167,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_118,
      O => rx_fifocheck_n0001(7)
    );
  rx_fifocheck_diff_6_CYINIT_1074 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_166,
      O => rx_fifocheck_diff_6_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_169_1075 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(8),
      IB => rx_fifocheck_diff_8_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_119,
      O => rx_fifocheck_Msub_n0001_inst_cy_169
    );
  rx_fifocheck_Msub_n0001_inst_sum_151 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_8_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_119,
      O => rx_fifocheck_n0001(8)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1191 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(8),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(8),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_119
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1201 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_fifocheck_bpl(9),
      O => rx_fifocheck_Msub_n0001_inst_lut2_120
    );
  rx_fifocheck_diff_8_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_8_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_170
    );
  rx_fifocheck_Msub_n0001_inst_cy_170_1076 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(9),
      IB => rx_fifocheck_Msub_n0001_inst_cy_169,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_120,
      O => rx_fifocheck_diff_8_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_152 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_169,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_120,
      O => rx_fifocheck_n0001(9)
    );
  rx_fifocheck_diff_8_CYINIT_1077 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_168,
      O => rx_fifocheck_diff_8_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_171_1078 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(10),
      IB => rx_fifocheck_diff_10_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_121,
      O => rx_fifocheck_Msub_n0001_inst_cy_171
    );
  rx_fifocheck_Msub_n0001_inst_sum_153 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_10_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_121,
      O => rx_fifocheck_n0001(10)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1211 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(10),
      ADR1 => rx_fifocheck_bpl(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_121
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1221 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(11),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(11),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_122
    );
  rx_fifocheck_diff_10_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_10_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_172
    );
  rx_fifocheck_Msub_n0001_inst_cy_172_1079 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(11),
      IB => rx_fifocheck_Msub_n0001_inst_cy_171,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_122,
      O => rx_fifocheck_diff_10_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_154 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_171,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_122,
      O => rx_fifocheck_n0001(11)
    );
  rx_fifocheck_diff_10_CYINIT_1080 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_170,
      O => rx_fifocheck_diff_10_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_173_1081 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(12),
      IB => rx_fifocheck_diff_12_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_123,
      O => rx_fifocheck_Msub_n0001_inst_cy_173
    );
  rx_fifocheck_Msub_n0001_inst_sum_155 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_12_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_123,
      O => rx_fifocheck_n0001(12)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1231 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(12),
      ADR1 => rx_fifocheck_bpl(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_123
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1241 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(13),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(13),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_124
    );
  rx_fifocheck_diff_12_COUTUSED : X_BUF
    port map (
      I => rx_fifocheck_diff_12_CYMUXG,
      O => rx_fifocheck_Msub_n0001_inst_cy_174
    );
  rx_fifocheck_Msub_n0001_inst_cy_174_1082 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(13),
      IB => rx_fifocheck_Msub_n0001_inst_cy_173,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_124,
      O => rx_fifocheck_diff_12_CYMUXG
    );
  rx_fifocheck_Msub_n0001_inst_sum_156 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_173,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_124,
      O => rx_fifocheck_n0001(13)
    );
  rx_fifocheck_diff_12_CYINIT_1083 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_172,
      O => rx_fifocheck_diff_12_CYINIT
    );
  rx_fifocheck_Msub_n0001_inst_cy_175_1084 : X_MUX2
    port map (
      IA => rx_fifocheck_fbbpl(14),
      IB => rx_fifocheck_diff_14_CYINIT,
      SEL => rx_fifocheck_Msub_n0001_inst_lut2_125,
      O => rx_fifocheck_Msub_n0001_inst_cy_175
    );
  rx_fifocheck_Msub_n0001_inst_sum_157 : X_XOR2
    port map (
      I0 => rx_fifocheck_diff_14_CYINIT,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_125,
      O => rx_fifocheck_n0001(14)
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1251 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(14),
      ADR1 => rx_fifocheck_bpl(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_125
    );
  rx_fifocheck_Msub_n0001_inst_lut2_1261 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_fifocheck_fbbpl(15),
      ADR1 => VCC,
      ADR2 => rx_fifocheck_bpl(15),
      ADR3 => VCC,
      O => rx_fifocheck_Msub_n0001_inst_lut2_126
    );
  rx_fifocheck_Msub_n0001_inst_sum_158 : X_XOR2
    port map (
      I0 => rx_fifocheck_Msub_n0001_inst_cy_175,
      I1 => rx_fifocheck_Msub_n0001_inst_lut2_126,
      O => rx_fifocheck_n0001(15)
    );
  rx_fifocheck_diff_14_CYINIT_1085 : X_BUF
    port map (
      I => rx_fifocheck_Msub_n0001_inst_cy_174,
      O => rx_fifocheck_diff_14_CYINIT
    );
  tx_fifocheck_diff_0_LOGIC_ONE_1086 : X_ONE
    port map (
      O => tx_fifocheck_diff_0_LOGIC_ONE
    );
  tx_fifocheck_Msub_n0001_inst_cy_161_1087 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(0),
      IB => tx_fifocheck_diff_0_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_111,
      O => tx_fifocheck_Msub_n0001_inst_cy_161
    );
  tx_fifocheck_Msub_n0001_inst_sum_143 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_0_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_111,
      O => tx_fifocheck_n0001(0)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1111 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(0),
      O => tx_fifocheck_Msub_n0001_inst_lut2_111
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1121 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(1),
      ADR1 => VCC,
      ADR2 => tx_fifocheck_bpl(1),
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_112
    );
  tx_fifocheck_diff_0_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_0_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_162
    );
  tx_fifocheck_Msub_n0001_inst_cy_162_1088 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(1),
      IB => tx_fifocheck_Msub_n0001_inst_cy_161,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_112,
      O => tx_fifocheck_diff_0_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_144 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_161,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_112,
      O => tx_fifocheck_n0001(1)
    );
  tx_fifocheck_diff_0_CYINIT_1089 : X_BUF
    port map (
      I => tx_fifocheck_diff_0_LOGIC_ONE,
      O => tx_fifocheck_diff_0_CYINIT
    );
  tx_fifocheck_diff_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_2_FFY_RST
    );
  tx_fifocheck_diff_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_2_FFY_RST,
      O => tx_fifocheck_diff(3)
    );
  tx_fifocheck_Msub_n0001_inst_cy_163_1090 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(2),
      IB => tx_fifocheck_diff_2_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_113,
      O => tx_fifocheck_Msub_n0001_inst_cy_163
    );
  tx_fifocheck_Msub_n0001_inst_sum_145 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_2_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_113,
      O => tx_fifocheck_n0001(2)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1131 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(2),
      ADR1 => tx_fifocheck_bpl(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_113
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1141 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(3),
      ADR1 => tx_fifocheck_bpl(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_114
    );
  tx_fifocheck_diff_2_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_2_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_164
    );
  tx_fifocheck_Msub_n0001_inst_cy_164_1091 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(3),
      IB => tx_fifocheck_Msub_n0001_inst_cy_163,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_114,
      O => tx_fifocheck_diff_2_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_146 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_163,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_114,
      O => tx_fifocheck_n0001(3)
    );
  tx_fifocheck_diff_2_CYINIT_1092 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_162,
      O => tx_fifocheck_diff_2_CYINIT
    );
  tx_fifocheck_diff_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_4_FFY_RST
    );
  tx_fifocheck_diff_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_4_FFY_RST,
      O => tx_fifocheck_diff(5)
    );
  tx_fifocheck_Msub_n0001_inst_cy_165_1093 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(4),
      IB => tx_fifocheck_diff_4_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_115,
      O => tx_fifocheck_Msub_n0001_inst_cy_165
    );
  tx_fifocheck_Msub_n0001_inst_sum_147 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_4_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_115,
      O => tx_fifocheck_n0001(4)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1151 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(4),
      ADR1 => VCC,
      ADR2 => tx_fifocheck_bpl(4),
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_115
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1161 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(5),
      O => tx_fifocheck_Msub_n0001_inst_lut2_116
    );
  tx_fifocheck_diff_4_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_4_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_166
    );
  tx_fifocheck_Msub_n0001_inst_cy_166_1094 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(5),
      IB => tx_fifocheck_Msub_n0001_inst_cy_165,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_116,
      O => tx_fifocheck_diff_4_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_148 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_165,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_116,
      O => tx_fifocheck_n0001(5)
    );
  tx_fifocheck_diff_4_CYINIT_1095 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_164,
      O => tx_fifocheck_diff_4_CYINIT
    );
  tx_fifocheck_diff_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_6_FFY_RST
    );
  tx_fifocheck_diff_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_6_FFY_RST,
      O => tx_fifocheck_diff(7)
    );
  tx_fifocheck_Msub_n0001_inst_cy_167_1096 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(6),
      IB => tx_fifocheck_diff_6_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_117,
      O => tx_fifocheck_Msub_n0001_inst_cy_167
    );
  tx_fifocheck_Msub_n0001_inst_sum_149 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_6_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_117,
      O => tx_fifocheck_n0001(6)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1171 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(6),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(6),
      O => tx_fifocheck_Msub_n0001_inst_lut2_117
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1181 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(7),
      ADR1 => VCC,
      ADR2 => tx_fifocheck_bpl(7),
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_118
    );
  tx_fifocheck_diff_6_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_6_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_168
    );
  tx_fifocheck_Msub_n0001_inst_cy_168_1097 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(7),
      IB => tx_fifocheck_Msub_n0001_inst_cy_167,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_118,
      O => tx_fifocheck_diff_6_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_150 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_167,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_118,
      O => tx_fifocheck_n0001(7)
    );
  tx_fifocheck_diff_6_CYINIT_1098 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_166,
      O => tx_fifocheck_diff_6_CYINIT
    );
  tx_fifocheck_diff_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_8_FFY_RST
    );
  tx_fifocheck_diff_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_8_FFY_RST,
      O => tx_fifocheck_diff(9)
    );
  tx_fifocheck_Msub_n0001_inst_cy_169_1099 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(8),
      IB => tx_fifocheck_diff_8_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_119,
      O => tx_fifocheck_Msub_n0001_inst_cy_169
    );
  tx_fifocheck_Msub_n0001_inst_sum_151 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_8_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_119,
      O => tx_fifocheck_n0001(8)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1191 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(8),
      ADR1 => tx_fifocheck_bpl(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_119
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1201 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(9),
      ADR1 => tx_fifocheck_bpl(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_120
    );
  tx_fifocheck_diff_8_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_8_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_170
    );
  tx_fifocheck_Msub_n0001_inst_cy_170_1100 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(9),
      IB => tx_fifocheck_Msub_n0001_inst_cy_169,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_120,
      O => tx_fifocheck_diff_8_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_152 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_169,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_120,
      O => tx_fifocheck_n0001(9)
    );
  tx_fifocheck_diff_8_CYINIT_1101 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_168,
      O => tx_fifocheck_diff_8_CYINIT
    );
  rx_input_fifo_control_DATA_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(3),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_3_FFY_RST,
      O => rx_input_data(3)
    );
  rx_input_data_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_3_FFY_RST
    );
  tx_fifocheck_diff_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_10_FFY_RST
    );
  tx_fifocheck_diff_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_10_FFY_RST,
      O => tx_fifocheck_diff(11)
    );
  tx_fifocheck_Msub_n0001_inst_cy_171_1102 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(10),
      IB => tx_fifocheck_diff_10_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_121,
      O => tx_fifocheck_Msub_n0001_inst_cy_171
    );
  tx_fifocheck_Msub_n0001_inst_sum_153 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_10_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_121,
      O => tx_fifocheck_n0001(10)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1211 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(10),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(10),
      O => tx_fifocheck_Msub_n0001_inst_lut2_121
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1221 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(11),
      ADR1 => VCC,
      ADR2 => tx_fifocheck_bpl(11),
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_122
    );
  tx_fifocheck_diff_10_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_10_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_172
    );
  tx_fifocheck_Msub_n0001_inst_cy_172_1103 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(11),
      IB => tx_fifocheck_Msub_n0001_inst_cy_171,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_122,
      O => tx_fifocheck_diff_10_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_154 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_171,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_122,
      O => tx_fifocheck_n0001(11)
    );
  tx_fifocheck_diff_10_CYINIT_1104 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_170,
      O => tx_fifocheck_diff_10_CYINIT
    );
  tx_fifocheck_diff_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_12_FFY_RST
    );
  tx_fifocheck_diff_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_12_FFY_RST,
      O => tx_fifocheck_diff(13)
    );
  tx_fifocheck_Msub_n0001_inst_cy_173_1105 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(12),
      IB => tx_fifocheck_diff_12_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_123,
      O => tx_fifocheck_Msub_n0001_inst_cy_173
    );
  tx_fifocheck_Msub_n0001_inst_sum_155 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_12_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_123,
      O => tx_fifocheck_n0001(12)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1231 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(12),
      ADR1 => tx_fifocheck_bpl(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_123
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1241 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(13),
      ADR1 => tx_fifocheck_bpl(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_124
    );
  tx_fifocheck_diff_12_COUTUSED : X_BUF
    port map (
      I => tx_fifocheck_diff_12_CYMUXG,
      O => tx_fifocheck_Msub_n0001_inst_cy_174
    );
  tx_fifocheck_Msub_n0001_inst_cy_174_1106 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(13),
      IB => tx_fifocheck_Msub_n0001_inst_cy_173,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_124,
      O => tx_fifocheck_diff_12_CYMUXG
    );
  tx_fifocheck_Msub_n0001_inst_sum_156 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_173,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_124,
      O => tx_fifocheck_n0001(13)
    );
  tx_fifocheck_diff_12_CYINIT_1107 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_172,
      O => tx_fifocheck_diff_12_CYINIT
    );
  tx_fifocheck_diff_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_14_FFY_RST
    );
  tx_fifocheck_diff_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_14_FFY_RST,
      O => tx_fifocheck_diff(15)
    );
  tx_fifocheck_Msub_n0001_inst_cy_175_1108 : X_MUX2
    port map (
      IA => tx_fifocheck_fbbpl(14),
      IB => tx_fifocheck_diff_14_CYINIT,
      SEL => tx_fifocheck_Msub_n0001_inst_lut2_125,
      O => tx_fifocheck_Msub_n0001_inst_cy_175
    );
  tx_fifocheck_Msub_n0001_inst_sum_157 : X_XOR2
    port map (
      I0 => tx_fifocheck_diff_14_CYINIT,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_125,
      O => tx_fifocheck_n0001(14)
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1251 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(14),
      ADR1 => VCC,
      ADR2 => tx_fifocheck_bpl(14),
      ADR3 => VCC,
      O => tx_fifocheck_Msub_n0001_inst_lut2_125
    );
  tx_fifocheck_Msub_n0001_inst_lut2_1261 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => tx_fifocheck_fbbpl(15),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_bpl(15),
      O => tx_fifocheck_Msub_n0001_inst_lut2_126
    );
  tx_fifocheck_Msub_n0001_inst_sum_158 : X_XOR2
    port map (
      I0 => tx_fifocheck_Msub_n0001_inst_cy_175,
      I1 => tx_fifocheck_Msub_n0001_inst_lut2_126,
      O => tx_fifocheck_n0001(15)
    );
  tx_fifocheck_diff_14_CYINIT_1109 : X_BUF
    port map (
      I => tx_fifocheck_Msub_n0001_inst_cy_174,
      O => tx_fifocheck_diff_14_CYINIT
    );
  mac_control_ledtx_cnt_142_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_142_FFY_RST
    );
  mac_control_ledtx_cnt_142_1110 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_289,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_142_FFY_RST,
      O => mac_control_ledtx_cnt_142
    );
  mac_control_ledtx_cnt_142_LOGIC_ONE_1111 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_142_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_327_1112 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_18,
      IB => mac_control_ledtx_cnt_142_LOGIC_ONE,
      SEL => mac_control_ledtx_rst_rt,
      O => mac_control_ledtx_cnt_inst_cy_327
    );
  mac_control_ledtx_rst_rt_1113 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_18,
      ADR1 => mac_control_ledtx_rst,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_ledtx_rst_rt
    );
  mac_control_ledtx_cnt_inst_lut3_2241 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_11,
      ADR1 => VCC,
      ADR2 => mac_control_ledtx_rst,
      ADR3 => mac_control_ledtx_cnt_142,
      O => mac_control_ledtx_cnt_inst_lut3_224
    );
  mac_control_ledtx_cnt_142_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_142_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_328
    );
  mac_control_ledtx_cnt_inst_cy_328_1114 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_11,
      IB => mac_control_ledtx_cnt_inst_cy_327,
      SEL => mac_control_ledtx_cnt_inst_lut3_224,
      O => mac_control_ledtx_cnt_142_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_289_1115 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_327,
      I1 => mac_control_ledtx_cnt_inst_lut3_224,
      O => mac_control_ledtx_cnt_inst_sum_289
    );
  mac_control_ledtx_cnt_143_LOGIC_ONE_1116 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_143_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_329_1117 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_143_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_143_CYINIT,
      SEL => mac_control_ledtx_cnt_inst_lut3_225,
      O => mac_control_ledtx_cnt_inst_cy_329
    );
  mac_control_ledtx_cnt_inst_sum_290_1118 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_143_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_225,
      O => mac_control_ledtx_cnt_inst_sum_290
    );
  mac_control_ledtx_cnt_inst_lut3_2251 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledtx_cnt_143,
      ADR2 => mac_control_ledtx_rst,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_225
    );
  mac_control_ledtx_cnt_inst_lut3_2261 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledtx_rst,
      ADR3 => mac_control_ledtx_cnt_144,
      O => mac_control_ledtx_cnt_inst_lut3_226
    );
  mac_control_ledtx_cnt_143_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_143_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_330
    );
  mac_control_ledtx_cnt_inst_cy_330_1119 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_143_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_inst_cy_329,
      SEL => mac_control_ledtx_cnt_inst_lut3_226,
      O => mac_control_ledtx_cnt_143_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_291_1120 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_329,
      I1 => mac_control_ledtx_cnt_inst_lut3_226,
      O => mac_control_ledtx_cnt_inst_sum_291
    );
  mac_control_ledtx_cnt_143_CYINIT_1121 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_328,
      O => mac_control_ledtx_cnt_143_CYINIT
    );
  mac_control_ledtx_cnt_145_LOGIC_ONE_1122 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_145_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_331_1123 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_145_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_145_CYINIT,
      SEL => mac_control_ledtx_cnt_inst_lut3_227,
      O => mac_control_ledtx_cnt_inst_cy_331
    );
  mac_control_ledtx_cnt_inst_sum_292_1124 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_145_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_227,
      O => mac_control_ledtx_cnt_inst_sum_292
    );
  mac_control_ledtx_cnt_inst_lut3_2271 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledtx_rst,
      ADR2 => mac_control_ledtx_cnt_145,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_227
    );
  mac_control_ledtx_cnt_inst_lut3_2281 : X_LUT4
    generic map(
      INIT => X"0303"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_ledtx_rst,
      ADR2 => mac_control_ledtx_cnt_146,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_228
    );
  mac_control_ledtx_cnt_145_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_145_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_332
    );
  mac_control_ledtx_cnt_inst_cy_332_1125 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_145_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_inst_cy_331,
      SEL => mac_control_ledtx_cnt_inst_lut3_228,
      O => mac_control_ledtx_cnt_145_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_293_1126 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_331,
      I1 => mac_control_ledtx_cnt_inst_lut3_228,
      O => mac_control_ledtx_cnt_inst_sum_293
    );
  mac_control_ledtx_cnt_145_CYINIT_1127 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_330,
      O => mac_control_ledtx_cnt_145_CYINIT
    );
  mac_control_ledtx_cnt_147_LOGIC_ONE_1128 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_147_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_333_1129 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_147_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_147_CYINIT,
      SEL => mac_control_ledtx_cnt_inst_lut3_229,
      O => mac_control_ledtx_cnt_inst_cy_333
    );
  mac_control_ledtx_cnt_inst_sum_294_1130 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_147_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_229,
      O => mac_control_ledtx_cnt_inst_sum_294
    );
  mac_control_ledtx_cnt_inst_lut3_2291 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => mac_control_ledtx_rst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_ledtx_cnt_147,
      O => mac_control_ledtx_cnt_inst_lut3_229
    );
  mac_control_ledtx_cnt_inst_lut3_2301 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => mac_control_ledtx_rst,
      ADR1 => VCC,
      ADR2 => mac_control_ledtx_cnt_148,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_230
    );
  mac_control_ledtx_cnt_147_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_147_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_334
    );
  mac_control_ledtx_cnt_inst_cy_334_1131 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_147_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_inst_cy_333,
      SEL => mac_control_ledtx_cnt_inst_lut3_230,
      O => mac_control_ledtx_cnt_147_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_295_1132 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_333,
      I1 => mac_control_ledtx_cnt_inst_lut3_230,
      O => mac_control_ledtx_cnt_inst_sum_295
    );
  mac_control_ledtx_cnt_147_CYINIT_1133 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_332,
      O => mac_control_ledtx_cnt_147_CYINIT
    );
  mac_control_ledtx_cnt_149_LOGIC_ONE_1134 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_149_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_335_1135 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_149_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_149_CYINIT,
      SEL => mac_control_ledtx_cnt_inst_lut3_231,
      O => mac_control_ledtx_cnt_inst_cy_335
    );
  mac_control_ledtx_cnt_inst_sum_296_1136 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_149_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_231,
      O => mac_control_ledtx_cnt_inst_sum_296
    );
  mac_control_ledtx_cnt_inst_lut3_2311 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => mac_control_ledtx_rst,
      ADR1 => VCC,
      ADR2 => mac_control_ledtx_cnt_149,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_231
    );
  mac_control_ledtx_cnt_inst_lut3_2321 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => mac_control_ledtx_rst,
      ADR1 => VCC,
      ADR2 => mac_control_ledtx_cnt_150,
      ADR3 => VCC,
      O => mac_control_ledtx_cnt_inst_lut3_232
    );
  mac_control_ledtx_cnt_149_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_149_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_336
    );
  mac_control_ledtx_cnt_inst_cy_336_1137 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_149_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_inst_cy_335,
      SEL => mac_control_ledtx_cnt_inst_lut3_232,
      O => mac_control_ledtx_cnt_149_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_297_1138 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_335,
      I1 => mac_control_ledtx_cnt_inst_lut3_232,
      O => mac_control_ledtx_cnt_inst_sum_297
    );
  mac_control_ledtx_cnt_149_CYINIT_1139 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_334,
      O => mac_control_ledtx_cnt_149_CYINIT
    );
  mac_control_ledtx_cnt_151_LOGIC_ONE_1140 : X_ONE
    port map (
      O => mac_control_ledtx_cnt_151_LOGIC_ONE
    );
  mac_control_ledtx_cnt_inst_cy_337_1141 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_151_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_151_CYINIT,
      SEL => mac_control_ledtx_cnt_inst_lut3_233,
      O => mac_control_ledtx_cnt_inst_cy_337
    );
  mac_control_ledtx_cnt_inst_sum_298_1142 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_151_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_233,
      O => mac_control_ledtx_cnt_inst_sum_298
    );
  mac_control_ledtx_cnt_inst_lut3_2331 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => mac_control_ledtx_rst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_ledtx_cnt_151,
      O => mac_control_ledtx_cnt_inst_lut3_233
    );
  mac_control_ledtx_cnt_inst_lut3_2341 : X_LUT4
    generic map(
      INIT => X"0055"
    )
    port map (
      ADR0 => mac_control_ledtx_rst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_ledtx_cnt_152,
      O => mac_control_ledtx_cnt_inst_lut3_234
    );
  mac_control_ledtx_cnt_151_COUTUSED : X_BUF
    port map (
      I => mac_control_ledtx_cnt_151_CYMUXG,
      O => mac_control_ledtx_cnt_inst_cy_338
    );
  mac_control_ledtx_cnt_inst_cy_338_1143 : X_MUX2
    port map (
      IA => mac_control_ledtx_cnt_151_LOGIC_ONE,
      IB => mac_control_ledtx_cnt_inst_cy_337,
      SEL => mac_control_ledtx_cnt_inst_lut3_234,
      O => mac_control_ledtx_cnt_151_CYMUXG
    );
  mac_control_ledtx_cnt_inst_sum_299_1144 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_inst_cy_337,
      I1 => mac_control_ledtx_cnt_inst_lut3_234,
      O => mac_control_ledtx_cnt_inst_sum_299
    );
  mac_control_ledtx_cnt_151_CYINIT_1145 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_336,
      O => mac_control_ledtx_cnt_151_CYINIT
    );
  mac_control_ledtx_cnt_inst_sum_300_1146 : X_XOR2
    port map (
      I0 => mac_control_ledtx_cnt_153_CYINIT,
      I1 => mac_control_ledtx_cnt_inst_lut3_235,
      O => mac_control_ledtx_cnt_inst_sum_300
    );
  mac_control_ledtx_cnt_inst_lut3_2351 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_ledtx_rst,
      ADR3 => mac_control_ledtx_cnt_153,
      O => mac_control_ledtx_cnt_inst_lut3_235
    );
  mac_control_ledtx_cnt_153_CYINIT_1147 : X_BUF
    port map (
      I => mac_control_ledtx_cnt_inst_cy_338,
      O => mac_control_ledtx_cnt_153_CYINIT
    );
  tx_output_bcnt_53_1148 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_186,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_53_FFX_RST,
      O => tx_output_bcnt_53
    );
  tx_output_bcnt_53_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_53_FFX_RST
    );
  rx_output_fifo_N17_LOGIC_ZERO_1149 : X_ZERO
    port map (
      O => rx_output_fifo_N17_LOGIC_ZERO
    );
  rx_output_fifo_BU38 : X_MUX2
    port map (
      IA => rx_output_fifo_N17,
      IB => rx_output_fifo_N17_CYINIT,
      SEL => rx_output_fifo_N1912,
      O => rx_output_fifo_N1914
    );
  rx_output_fifo_BU39 : X_XOR2
    port map (
      I0 => rx_output_fifo_N17_CYINIT,
      I1 => rx_output_fifo_N1912,
      O => rx_output_fifo_N1904
    );
  rx_output_fifo_BU37 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_output_fifo_N17,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N1912
    );
  rx_output_fifo_N17_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N16,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N17_GROM
    );
  rx_output_fifo_N17_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N17_CYMUXG,
      O => rx_output_fifo_N1919
    );
  rx_output_fifo_BU44 : X_MUX2
    port map (
      IA => rx_output_fifo_N16,
      IB => rx_output_fifo_N1914,
      SEL => rx_output_fifo_N17_GROM,
      O => rx_output_fifo_N17_CYMUXG
    );
  rx_output_fifo_BU45 : X_XOR2
    port map (
      I0 => rx_output_fifo_N1914,
      I1 => rx_output_fifo_N17_GROM,
      O => rx_output_fifo_N1905
    );
  rx_output_fifo_N17_CYINIT_1150 : X_BUF
    port map (
      I => rx_output_fifo_N17_LOGIC_ZERO,
      O => rx_output_fifo_N17_CYINIT
    );
  rx_output_fifo_BU50 : X_MUX2
    port map (
      IA => rx_output_fifo_N15,
      IB => rx_output_fifo_N15_CYINIT,
      SEL => rx_output_fifo_N15_FROM,
      O => rx_output_fifo_N1924
    );
  rx_output_fifo_BU51 : X_XOR2
    port map (
      I0 => rx_output_fifo_N15_CYINIT,
      I1 => rx_output_fifo_N15_FROM,
      O => rx_output_fifo_N1906
    );
  rx_output_fifo_N15_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N15,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N15_FROM
    );
  rx_output_fifo_N15_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N14,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N15_GROM
    );
  rx_output_fifo_N15_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N15_CYMUXG,
      O => rx_output_fifo_N1929
    );
  rx_output_fifo_BU56 : X_MUX2
    port map (
      IA => rx_output_fifo_N14,
      IB => rx_output_fifo_N1924,
      SEL => rx_output_fifo_N15_GROM,
      O => rx_output_fifo_N15_CYMUXG
    );
  rx_output_fifo_BU57 : X_XOR2
    port map (
      I0 => rx_output_fifo_N1924,
      I1 => rx_output_fifo_N15_GROM,
      O => rx_output_fifo_N1907
    );
  rx_output_fifo_N15_CYINIT_1151 : X_BUF
    port map (
      I => rx_output_fifo_N1919,
      O => rx_output_fifo_N15_CYINIT
    );
  rx_output_fifo_BU62 : X_MUX2
    port map (
      IA => rx_output_fifo_N13,
      IB => rx_output_fifo_N13_CYINIT,
      SEL => rx_output_fifo_N13_FROM,
      O => rx_output_fifo_N1934
    );
  rx_output_fifo_BU63 : X_XOR2
    port map (
      I0 => rx_output_fifo_N13_CYINIT,
      I1 => rx_output_fifo_N13_FROM,
      O => rx_output_fifo_N1908
    );
  rx_output_fifo_N13_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N13,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N13_FROM
    );
  rx_output_fifo_N13_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N12,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N13_GROM
    );
  rx_output_fifo_N13_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N13_CYMUXG,
      O => rx_output_fifo_N1939
    );
  rx_output_fifo_BU68 : X_MUX2
    port map (
      IA => rx_output_fifo_N12,
      IB => rx_output_fifo_N1934,
      SEL => rx_output_fifo_N13_GROM,
      O => rx_output_fifo_N13_CYMUXG
    );
  rx_output_fifo_BU69 : X_XOR2
    port map (
      I0 => rx_output_fifo_N1934,
      I1 => rx_output_fifo_N13_GROM,
      O => rx_output_fifo_N1909
    );
  rx_output_fifo_N13_CYINIT_1152 : X_BUF
    port map (
      I => rx_output_fifo_N1929,
      O => rx_output_fifo_N13_CYINIT
    );
  rx_output_fifo_BU74 : X_MUX2
    port map (
      IA => rx_output_fifo_N11,
      IB => rx_output_fifo_N11_CYINIT,
      SEL => rx_output_fifo_N11_FROM,
      O => rx_output_fifo_N1944
    );
  rx_output_fifo_BU75 : X_XOR2
    port map (
      I0 => rx_output_fifo_N11_CYINIT,
      I1 => rx_output_fifo_N11_FROM,
      O => rx_output_fifo_N1910
    );
  rx_output_fifo_N11_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N11,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N11_FROM
    );
  rx_output_fifo_N10_rt_1153 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N10,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N10_rt
    );
  rx_output_fifo_BU80 : X_XOR2
    port map (
      I0 => rx_output_fifo_N1944,
      I1 => rx_output_fifo_N10_rt,
      O => rx_output_fifo_N1911
    );
  rx_output_fifo_N11_CYINIT_1154 : X_BUF
    port map (
      I => rx_output_fifo_N1939,
      O => rx_output_fifo_N11_CYINIT
    );
  tx_input_n0074_0_LOGIC_ONE_1155 : X_ONE
    port map (
      O => tx_input_n0074_0_LOGIC_ONE
    );
  tx_input_Msub_n0034_inst_cy_118_1156 : X_MUX2
    port map (
      IA => tx_input_CNT(0),
      IB => tx_input_n0074_0_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_95,
      O => tx_input_Msub_n0034_inst_cy_118
    );
  tx_input_Msub_n0034_inst_sum_111 : X_XOR2
    port map (
      I0 => tx_input_n0074_0_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_95,
      O => tx_input_n0074_0_XORF
    );
  tx_input_Msub_n0034_inst_lut2_951 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_95
    );
  tx_input_n0074_0_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_20,
      ADR1 => VCC,
      ADR2 => tx_input_CNT(1),
      ADR3 => VCC,
      O => tx_input_n0074_0_GROM
    );
  tx_input_n0074_0_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_0_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_119
    );
  tx_input_n0074_0_XUSED : X_BUF
    port map (
      I => tx_input_n0074_0_XORF,
      O => tx_input_n0074(0)
    );
  tx_input_n0074_0_YUSED : X_BUF
    port map (
      I => tx_input_n0074_0_XORG,
      O => tx_input_n0074(1)
    );
  tx_input_Msub_n0034_inst_cy_119_1157 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_20,
      IB => tx_input_Msub_n0034_inst_cy_118,
      SEL => tx_input_n0074_0_GROM,
      O => tx_input_n0074_0_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_112 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_118,
      I1 => tx_input_n0074_0_GROM,
      O => tx_input_n0074_0_XORG
    );
  tx_input_n0074_0_CYINIT_1158 : X_BUF
    port map (
      I => tx_input_n0074_0_LOGIC_ONE,
      O => tx_input_n0074_0_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_120_1159 : X_MUX2
    port map (
      IA => tx_input_CNT(2),
      IB => tx_input_n0074_2_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_97,
      O => tx_input_Msub_n0034_inst_cy_120
    );
  tx_input_Msub_n0034_inst_sum_113 : X_XOR2
    port map (
      I0 => tx_input_n0074_2_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_97,
      O => tx_input_n0074_2_XORF
    );
  tx_input_Msub_n0034_inst_lut2_971 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_97
    );
  tx_input_Msub_n0034_inst_lut2_981 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_98
    );
  tx_input_n0074_2_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_2_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_121
    );
  tx_input_n0074_2_XUSED : X_BUF
    port map (
      I => tx_input_n0074_2_XORF,
      O => tx_input_n0074(2)
    );
  tx_input_n0074_2_YUSED : X_BUF
    port map (
      I => tx_input_n0074_2_XORG,
      O => tx_input_n0074(3)
    );
  tx_input_Msub_n0034_inst_cy_121_1160 : X_MUX2
    port map (
      IA => tx_input_CNT(3),
      IB => tx_input_Msub_n0034_inst_cy_120,
      SEL => tx_input_Msub_n0034_inst_lut2_98,
      O => tx_input_n0074_2_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_114 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_120,
      I1 => tx_input_Msub_n0034_inst_lut2_98,
      O => tx_input_n0074_2_XORG
    );
  tx_input_n0074_2_CYINIT_1161 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_119,
      O => tx_input_n0074_2_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_122_1162 : X_MUX2
    port map (
      IA => tx_input_CNT(4),
      IB => tx_input_n0074_4_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_99,
      O => tx_input_Msub_n0034_inst_cy_122
    );
  tx_input_Msub_n0034_inst_sum_115 : X_XOR2
    port map (
      I0 => tx_input_n0074_4_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_99,
      O => tx_input_n0074_4_XORF
    );
  tx_input_Msub_n0034_inst_lut2_991 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_99
    );
  tx_input_Msub_n0034_inst_lut2_1001 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_100
    );
  tx_input_n0074_4_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_4_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_123
    );
  tx_input_n0074_4_XUSED : X_BUF
    port map (
      I => tx_input_n0074_4_XORF,
      O => tx_input_n0074(4)
    );
  tx_input_n0074_4_YUSED : X_BUF
    port map (
      I => tx_input_n0074_4_XORG,
      O => tx_input_n0074(5)
    );
  tx_input_Msub_n0034_inst_cy_123_1163 : X_MUX2
    port map (
      IA => tx_input_CNT(5),
      IB => tx_input_Msub_n0034_inst_cy_122,
      SEL => tx_input_Msub_n0034_inst_lut2_100,
      O => tx_input_n0074_4_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_116 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_122,
      I1 => tx_input_Msub_n0034_inst_lut2_100,
      O => tx_input_n0074_4_XORG
    );
  tx_input_n0074_4_CYINIT_1164 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_121,
      O => tx_input_n0074_4_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_124_1165 : X_MUX2
    port map (
      IA => tx_input_CNT(6),
      IB => tx_input_n0074_6_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_101,
      O => tx_input_Msub_n0034_inst_cy_124
    );
  tx_input_Msub_n0034_inst_sum_117 : X_XOR2
    port map (
      I0 => tx_input_n0074_6_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_101,
      O => tx_input_n0074_6_XORF
    );
  tx_input_Msub_n0034_inst_lut2_1011 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(6),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_101
    );
  tx_input_Msub_n0034_inst_lut2_1021 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(7),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_102
    );
  tx_input_n0074_6_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_6_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_125
    );
  tx_input_n0074_6_XUSED : X_BUF
    port map (
      I => tx_input_n0074_6_XORF,
      O => tx_input_n0074(6)
    );
  tx_input_n0074_6_YUSED : X_BUF
    port map (
      I => tx_input_n0074_6_XORG,
      O => tx_input_n0074(7)
    );
  tx_input_Msub_n0034_inst_cy_125_1166 : X_MUX2
    port map (
      IA => tx_input_CNT(7),
      IB => tx_input_Msub_n0034_inst_cy_124,
      SEL => tx_input_Msub_n0034_inst_lut2_102,
      O => tx_input_n0074_6_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_118 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_124,
      I1 => tx_input_Msub_n0034_inst_lut2_102,
      O => tx_input_n0074_6_XORG
    );
  tx_input_n0074_6_CYINIT_1167 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_123,
      O => tx_input_n0074_6_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_126_1168 : X_MUX2
    port map (
      IA => tx_input_CNT(8),
      IB => tx_input_n0074_8_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_103,
      O => tx_input_Msub_n0034_inst_cy_126
    );
  tx_input_Msub_n0034_inst_sum_119 : X_XOR2
    port map (
      I0 => tx_input_n0074_8_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_103,
      O => tx_input_n0074_8_XORF
    );
  tx_input_Msub_n0034_inst_lut2_1031 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_103
    );
  tx_input_Msub_n0034_inst_lut2_1041 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_104
    );
  tx_input_n0074_8_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_8_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_127
    );
  tx_input_n0074_8_XUSED : X_BUF
    port map (
      I => tx_input_n0074_8_XORF,
      O => tx_input_n0074(8)
    );
  tx_input_n0074_8_YUSED : X_BUF
    port map (
      I => tx_input_n0074_8_XORG,
      O => tx_input_n0074(9)
    );
  tx_input_Msub_n0034_inst_cy_127_1169 : X_MUX2
    port map (
      IA => tx_input_CNT(9),
      IB => tx_input_Msub_n0034_inst_cy_126,
      SEL => tx_input_Msub_n0034_inst_lut2_104,
      O => tx_input_n0074_8_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_120 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_126,
      I1 => tx_input_Msub_n0034_inst_lut2_104,
      O => tx_input_n0074_8_XORG
    );
  tx_input_n0074_8_CYINIT_1170 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_125,
      O => tx_input_n0074_8_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_128_1171 : X_MUX2
    port map (
      IA => tx_input_CNT(10),
      IB => tx_input_n0074_10_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_105,
      O => tx_input_Msub_n0034_inst_cy_128
    );
  tx_input_Msub_n0034_inst_sum_121 : X_XOR2
    port map (
      I0 => tx_input_n0074_10_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_105,
      O => tx_input_n0074_10_XORF
    );
  tx_input_Msub_n0034_inst_lut2_1051 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(10),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_105
    );
  tx_input_Msub_n0034_inst_lut2_1061 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(11),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_106
    );
  tx_input_n0074_10_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_10_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_129
    );
  tx_input_n0074_10_XUSED : X_BUF
    port map (
      I => tx_input_n0074_10_XORF,
      O => tx_input_n0074(10)
    );
  tx_input_n0074_10_YUSED : X_BUF
    port map (
      I => tx_input_n0074_10_XORG,
      O => tx_input_n0074(11)
    );
  tx_input_Msub_n0034_inst_cy_129_1172 : X_MUX2
    port map (
      IA => tx_input_CNT(11),
      IB => tx_input_Msub_n0034_inst_cy_128,
      SEL => tx_input_Msub_n0034_inst_lut2_106,
      O => tx_input_n0074_10_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_122 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_128,
      I1 => tx_input_Msub_n0034_inst_lut2_106,
      O => tx_input_n0074_10_XORG
    );
  tx_input_n0074_10_CYINIT_1173 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_127,
      O => tx_input_n0074_10_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_130_1174 : X_MUX2
    port map (
      IA => tx_input_CNT(12),
      IB => tx_input_n0074_12_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_107,
      O => tx_input_Msub_n0034_inst_cy_130
    );
  tx_input_Msub_n0034_inst_sum_123 : X_XOR2
    port map (
      I0 => tx_input_n0074_12_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_107,
      O => tx_input_n0074_12_XORF
    );
  tx_input_Msub_n0034_inst_lut2_1071 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(12),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_107
    );
  tx_input_Msub_n0034_inst_lut2_1081 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_108
    );
  tx_input_n0074_12_COUTUSED : X_BUF
    port map (
      I => tx_input_n0074_12_CYMUXG,
      O => tx_input_Msub_n0034_inst_cy_131
    );
  tx_input_n0074_12_XUSED : X_BUF
    port map (
      I => tx_input_n0074_12_XORF,
      O => tx_input_n0074(12)
    );
  tx_input_n0074_12_YUSED : X_BUF
    port map (
      I => tx_input_n0074_12_XORG,
      O => tx_input_n0074(13)
    );
  tx_input_Msub_n0034_inst_cy_131_1175 : X_MUX2
    port map (
      IA => tx_input_CNT(13),
      IB => tx_input_Msub_n0034_inst_cy_130,
      SEL => tx_input_Msub_n0034_inst_lut2_108,
      O => tx_input_n0074_12_CYMUXG
    );
  tx_input_Msub_n0034_inst_sum_124 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_130,
      I1 => tx_input_Msub_n0034_inst_lut2_108,
      O => tx_input_n0074_12_XORG
    );
  tx_input_n0074_12_CYINIT_1176 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_129,
      O => tx_input_n0074_12_CYINIT
    );
  tx_input_Msub_n0034_inst_cy_132_1177 : X_MUX2
    port map (
      IA => tx_input_CNT(14),
      IB => tx_input_n0074_14_CYINIT,
      SEL => tx_input_Msub_n0034_inst_lut2_109,
      O => tx_input_Msub_n0034_inst_cy_132
    );
  tx_input_Msub_n0034_inst_sum_125 : X_XOR2
    port map (
      I0 => tx_input_n0074_14_CYINIT,
      I1 => tx_input_Msub_n0034_inst_lut2_109,
      O => tx_input_n0074_14_XORF
    );
  tx_input_Msub_n0034_inst_lut2_1091 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(14),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_109
    );
  tx_input_Msub_n0034_inst_lut2_1101 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => tx_input_CNT(15),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_input_Msub_n0034_inst_lut2_110
    );
  tx_input_n0074_14_XUSED : X_BUF
    port map (
      I => tx_input_n0074_14_XORF,
      O => tx_input_n0074(14)
    );
  tx_input_n0074_14_YUSED : X_BUF
    port map (
      I => tx_input_n0074_14_XORG,
      O => tx_input_n0074(15)
    );
  tx_input_Msub_n0034_inst_sum_126 : X_XOR2
    port map (
      I0 => tx_input_Msub_n0034_inst_cy_132,
      I1 => tx_input_Msub_n0034_inst_lut2_110,
      O => tx_input_n0074_14_XORG
    );
  tx_input_n0074_14_CYINIT_1178 : X_BUF
    port map (
      I => tx_input_Msub_n0034_inst_cy_131,
      O => tx_input_n0074_14_CYINIT
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ONE_1179 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ZERO_1180 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_177_1181 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(32),
      ADR1 => rx_input_memio_addrchk_macaddrl(33),
      ADR2 => rx_input_memio_addrchk_datal(33),
      ADR3 => rx_input_memio_addrchk_macaddrl(32),
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(34),
      ADR1 => rx_input_memio_addrchk_macaddrl(34),
      ADR2 => rx_input_memio_addrchk_macaddrl(35),
      ADR3 => rx_input_memio_addrchk_datal(35),
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_1182 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_1_LOGIC_ZERO_1183 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_1_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_179_1184 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_1_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_1_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(36),
      ADR1 => rx_input_memio_addrchk_macaddrl(37),
      ADR2 => rx_input_memio_addrchk_datal(37),
      ADR3 => rx_input_memio_addrchk_datal(36),
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(38),
      ADR1 => rx_input_memio_addrchk_macaddrl(38),
      ADR2 => rx_input_memio_addrchk_datal(39),
      ADR3 => rx_input_memio_addrchk_macaddrl(39),
      O => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_1_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_1_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(1)
    );
  rx_input_memio_addrchk_Mcompar_n0045_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_1_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0045_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_1_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_1_CYINIT_1185 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0045_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_1_CYINIT
    );
  mac_control_PHY_status_MII_Interface_mdccnt_32_LOGIC_ZERO_1186 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_mdccnt_32_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_187_1187 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_32,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_32_LOGIC_ZERO,
      SEL => mac_control_PHY_status_MII_Interface_cs_FFd5_rt,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_187
    );
  mac_control_PHY_status_MII_Interface_cs_FFd5_rt_1188 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_32,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_cs_FFd5_rt
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_341 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_49,
      ADR1 => mac_control_PHY_status_MII_Interface_mdccnt_32,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_34
    );
  mac_control_PHY_status_MII_Interface_mdccnt_32_COUTUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_32_CYMUXG,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_188
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_188_1189 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_49,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_187,
      SEL => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_34,
      O => mac_control_PHY_status_MII_Interface_mdccnt_32_CYMUXG
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_165_1190 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_187,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_34,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_165
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_LOGIC_ZERO_1191 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_mdccnt_33_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_189_1192 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_mdccnt_33_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_33_CYINIT,
      SEL => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_35,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_189
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_166_1193 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_33_CYINIT,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_35,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_166
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_351 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => mac_control_PHY_status_MII_Interface_mdccnt_33,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_35
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_361 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_mdccnt_34,
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_36
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_COUTUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_33_CYMUXG,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_190
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_190_1194 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_mdccnt_33_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_189,
      SEL => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_36,
      O => mac_control_PHY_status_MII_Interface_mdccnt_33_CYMUXG
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_167_1195 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_189,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_36,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_167
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_CYINIT_1196 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_188,
      O => mac_control_PHY_status_MII_Interface_mdccnt_33_CYINIT
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_LOGIC_ZERO_1197 : X_ZERO
    port map (
      O => mac_control_PHY_status_MII_Interface_mdccnt_35_LOGIC_ZERO
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_191_1198 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_mdccnt_35_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_35_CYINIT,
      SEL => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_37,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_191
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_168_1199 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_35_CYINIT,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_37,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_168
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_371 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_MII_Interface_mdccnt_35,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => VCC,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_37
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_381 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_mdccnt_36,
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_38
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_COUTUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_35_CYMUXG,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_192
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_192_1200 : X_MUX2
    port map (
      IA => mac_control_PHY_status_MII_Interface_mdccnt_35_LOGIC_ZERO,
      IB => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_191,
      SEL => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_38,
      O => mac_control_PHY_status_MII_Interface_mdccnt_35_CYMUXG
    );
  mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_169_1201 : X_XOR2
    port map (
      I0 => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_191,
      I1 => mac_control_PHY_status_MII_Interface_mdccnt_inst_lut3_38,
      O => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_169
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_CYINIT_1202 : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_cy_190,
      O => mac_control_PHY_status_MII_Interface_mdccnt_35_CYINIT
    );
  rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ONE_1203 : X_ONE
    port map (
      O => rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ONE
    );
  rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ZERO_1204 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ZERO
    );
  rx_output_Mcompar_n0018_inst_cy_78_1205 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ONE,
      SEL => rx_output_Mcompar_n0018_inst_lut4_0,
      O => rx_output_Mcompar_n0018_inst_cy_78
    );
  rx_output_Mcompar_n0018_inst_lut4_01 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rxfbbp(0),
      ADR1 => addr3ext(0),
      ADR2 => addr3ext(1),
      ADR3 => rxfbbp(1),
      O => rx_output_Mcompar_n0018_inst_lut4_0
    );
  rx_output_Mcompar_n0018_inst_lut4_11 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rxfbbp(3),
      ADR1 => rxfbbp(2),
      ADR2 => addr3ext(3),
      ADR3 => addr3ext(2),
      O => rx_output_Mcompar_n0018_inst_lut4_1
    );
  rx_output_Mcompar_n0018_inst_cy_79_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_79_CYMUXG,
      O => rx_output_Mcompar_n0018_inst_cy_79
    );
  rx_output_Mcompar_n0018_inst_cy_79_1206 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_79_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_78,
      SEL => rx_output_Mcompar_n0018_inst_lut4_1,
      O => rx_output_Mcompar_n0018_inst_cy_79_CYMUXG
    );
  rx_output_Mcompar_n0018_inst_cy_81_LOGIC_ZERO_1207 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0018_inst_cy_81_LOGIC_ZERO
    );
  rx_output_Mcompar_n0018_inst_cy_80_1208 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_81_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_81_CYINIT,
      SEL => rx_output_Mcompar_n0018_inst_lut4_2,
      O => rx_output_Mcompar_n0018_inst_cy_80
    );
  rx_output_Mcompar_n0018_inst_lut4_21 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => addr3ext(4),
      ADR1 => addr3ext(5),
      ADR2 => rxfbbp(4),
      ADR3 => rxfbbp(5),
      O => rx_output_Mcompar_n0018_inst_lut4_2
    );
  rx_output_Mcompar_n0018_inst_lut4_31 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => addr3ext(6),
      ADR1 => rxfbbp(6),
      ADR2 => addr3ext(7),
      ADR3 => rxfbbp(7),
      O => rx_output_Mcompar_n0018_inst_lut4_3
    );
  rx_output_Mcompar_n0018_inst_cy_81_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_81_CYMUXG,
      O => rx_output_Mcompar_n0018_inst_cy_81
    );
  rx_output_Mcompar_n0018_inst_cy_81_1209 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_81_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_80,
      SEL => rx_output_Mcompar_n0018_inst_lut4_3,
      O => rx_output_Mcompar_n0018_inst_cy_81_CYMUXG
    );
  rx_output_Mcompar_n0018_inst_cy_81_CYINIT_1210 : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_79,
      O => rx_output_Mcompar_n0018_inst_cy_81_CYINIT
    );
  rx_output_Mcompar_n0018_inst_cy_83_LOGIC_ZERO_1211 : X_ZERO
    port map (
      O => rx_output_Mcompar_n0018_inst_cy_83_LOGIC_ZERO
    );
  rx_output_Mcompar_n0018_inst_cy_82_1212 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_83_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_83_CYINIT,
      SEL => rx_output_Mcompar_n0018_inst_lut4_4,
      O => rx_output_Mcompar_n0018_inst_cy_82
    );
  rx_output_Mcompar_n0018_inst_lut4_41 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rxfbbp(9),
      ADR1 => addr3ext(8),
      ADR2 => addr3ext(9),
      ADR3 => rxfbbp(8),
      O => rx_output_Mcompar_n0018_inst_lut4_4
    );
  rx_output_Mcompar_n0018_inst_lut4_51 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => addr3ext(10),
      ADR1 => rxfbbp(10),
      ADR2 => addr3ext(11),
      ADR3 => rxfbbp(11),
      O => rx_output_Mcompar_n0018_inst_lut4_5
    );
  rx_output_Mcompar_n0018_inst_cy_83_COUTUSED : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_83_CYMUXG,
      O => rx_output_Mcompar_n0018_inst_cy_83
    );
  rx_output_Mcompar_n0018_inst_cy_83_1213 : X_MUX2
    port map (
      IA => rx_output_Mcompar_n0018_inst_cy_83_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_82,
      SEL => rx_output_Mcompar_n0018_inst_lut4_5,
      O => rx_output_Mcompar_n0018_inst_cy_83_CYMUXG
    );
  rx_output_Mcompar_n0018_inst_cy_83_CYINIT_1214 : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_81,
      O => rx_output_Mcompar_n0018_inst_cy_83_CYINIT
    );
  rx_output_n0018_LOGIC_ZERO_1215 : X_ZERO
    port map (
      O => rx_output_n0018_LOGIC_ZERO
    );
  rx_output_Mcompar_n0018_inst_cy_84_1216 : X_MUX2
    port map (
      IA => rx_output_n0018_LOGIC_ZERO,
      IB => rx_output_n0018_CYINIT,
      SEL => rx_output_Mcompar_n0018_inst_lut4_6,
      O => rx_output_Mcompar_n0018_inst_cy_84
    );
  rx_output_Mcompar_n0018_inst_lut4_61 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rxfbbp(12),
      ADR1 => rxfbbp(13),
      ADR2 => addr3ext(12),
      ADR3 => addr3ext(13),
      O => rx_output_Mcompar_n0018_inst_lut4_6
    );
  rx_output_Mcompar_n0018_inst_lut4_71 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rxfbbp(14),
      ADR1 => rxfbbp(15),
      ADR2 => addr3ext(14),
      ADR3 => addr3ext(15),
      O => rx_output_Mcompar_n0018_inst_lut4_7
    );
  rx_output_n0018_COUTUSED : X_BUF
    port map (
      I => rx_output_n0018_CYMUXG,
      O => rx_output_n0018
    );
  rx_output_Mcompar_n0018_inst_cy_85 : X_MUX2
    port map (
      IA => rx_output_n0018_LOGIC_ZERO,
      IB => rx_output_Mcompar_n0018_inst_cy_84,
      SEL => rx_output_Mcompar_n0018_inst_lut4_7,
      O => rx_output_n0018_CYMUXG
    );
  rx_output_n0018_CYINIT_1217 : X_BUF
    port map (
      I => rx_output_Mcompar_n0018_inst_cy_83,
      O => rx_output_n0018_CYINIT
    );
  mac_control_txf_cnt_0_LOGIC_ZERO_1218 : X_ZERO
    port map (
      O => mac_control_txf_cnt_0_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_16_1219 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_16,
      IB => mac_control_txf_cnt_0_LOGIC_ZERO,
      SEL => mac_control_txf_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_txf_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_16,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(0),
      O => mac_control_txf_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_txf_cnt_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_23,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(1),
      O => mac_control_txf_cnt_0_GROM
    );
  mac_control_txf_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_0_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_17_1220 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_23,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_txf_cnt_0_GROM,
      O => mac_control_txf_cnt_0_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_txf_cnt_0_GROM,
      O => mac_control_txf_cnt_n0000(1)
    );
  mac_control_txf_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(3),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(3)
    );
  mac_control_txf_cnt_2_LOGIC_ZERO_1221 : X_ZERO
    port map (
      O => mac_control_txf_cnt_2_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_18_1222 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_2_LOGIC_ZERO,
      IB => mac_control_txf_cnt_2_CYINIT,
      SEL => mac_control_txf_cnt_2_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_2_CYINIT,
      I1 => mac_control_txf_cnt_2_FROM,
      O => mac_control_txf_cnt_n0000(2)
    );
  mac_control_txf_cnt_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(2),
      O => mac_control_txf_cnt_2_FROM
    );
  mac_control_txf_cnt_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(3),
      O => mac_control_txf_cnt_2_GROM
    );
  mac_control_txf_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_2_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_19_1223 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_2_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_txf_cnt_2_GROM,
      O => mac_control_txf_cnt_2_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_txf_cnt_2_GROM,
      O => mac_control_txf_cnt_n0000(3)
    );
  mac_control_txf_cnt_2_CYINIT_1224 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_txf_cnt_2_CYINIT
    );
  mac_control_txf_cnt_4_LOGIC_ZERO_1225 : X_ZERO
    port map (
      O => mac_control_txf_cnt_4_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_20_1226 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_4_LOGIC_ZERO,
      IB => mac_control_txf_cnt_4_CYINIT,
      SEL => mac_control_txf_cnt_4_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_4_CYINIT,
      I1 => mac_control_txf_cnt_4_FROM,
      O => mac_control_txf_cnt_n0000(4)
    );
  mac_control_txf_cnt_4_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(4),
      O => mac_control_txf_cnt_4_FROM
    );
  mac_control_txf_cnt_4_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(5),
      O => mac_control_txf_cnt_4_GROM
    );
  mac_control_txf_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_4_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_21_1227 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_4_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_txf_cnt_4_GROM,
      O => mac_control_txf_cnt_4_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_txf_cnt_4_GROM,
      O => mac_control_txf_cnt_n0000(5)
    );
  mac_control_txf_cnt_4_CYINIT_1228 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_txf_cnt_4_CYINIT
    );
  mac_control_txf_cnt_6_LOGIC_ZERO_1229 : X_ZERO
    port map (
      O => mac_control_txf_cnt_6_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_22_1230 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_6_LOGIC_ZERO,
      IB => mac_control_txf_cnt_6_CYINIT,
      SEL => mac_control_txf_cnt_6_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_6_CYINIT,
      I1 => mac_control_txf_cnt_6_FROM,
      O => mac_control_txf_cnt_n0000(6)
    );
  mac_control_txf_cnt_6_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(6),
      O => mac_control_txf_cnt_6_FROM
    );
  mac_control_txf_cnt_6_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(7),
      O => mac_control_txf_cnt_6_GROM
    );
  mac_control_txf_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_6_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_23_1231 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_6_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_txf_cnt_6_GROM,
      O => mac_control_txf_cnt_6_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_txf_cnt_6_GROM,
      O => mac_control_txf_cnt_n0000(7)
    );
  mac_control_txf_cnt_6_CYINIT_1232 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_txf_cnt_6_CYINIT
    );
  mac_control_txf_cnt_8_LOGIC_ZERO_1233 : X_ZERO
    port map (
      O => mac_control_txf_cnt_8_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_24_1234 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_8_LOGIC_ZERO,
      IB => mac_control_txf_cnt_8_CYINIT,
      SEL => mac_control_txf_cnt_8_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_8_CYINIT,
      I1 => mac_control_txf_cnt_8_FROM,
      O => mac_control_txf_cnt_n0000(8)
    );
  mac_control_txf_cnt_8_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(8),
      O => mac_control_txf_cnt_8_FROM
    );
  mac_control_txf_cnt_8_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(9),
      O => mac_control_txf_cnt_8_GROM
    );
  mac_control_txf_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_8_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_25_1235 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_8_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_txf_cnt_8_GROM,
      O => mac_control_txf_cnt_8_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_txf_cnt_8_GROM,
      O => mac_control_txf_cnt_n0000(9)
    );
  mac_control_txf_cnt_8_CYINIT_1236 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_txf_cnt_8_CYINIT
    );
  mac_control_txf_cnt_10_LOGIC_ZERO_1237 : X_ZERO
    port map (
      O => mac_control_txf_cnt_10_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_26_1238 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_10_LOGIC_ZERO,
      IB => mac_control_txf_cnt_10_CYINIT,
      SEL => mac_control_txf_cnt_10_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_10_CYINIT,
      I1 => mac_control_txf_cnt_10_FROM,
      O => mac_control_txf_cnt_n0000(10)
    );
  mac_control_txf_cnt_10_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(10),
      O => mac_control_txf_cnt_10_FROM
    );
  mac_control_txf_cnt_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(11),
      O => mac_control_txf_cnt_10_GROM
    );
  mac_control_txf_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_10_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_27_1239 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_10_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_txf_cnt_10_GROM,
      O => mac_control_txf_cnt_10_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_txf_cnt_10_GROM,
      O => mac_control_txf_cnt_n0000(11)
    );
  mac_control_txf_cnt_10_CYINIT_1240 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_txf_cnt_10_CYINIT
    );
  mac_control_txf_cnt_12_LOGIC_ZERO_1241 : X_ZERO
    port map (
      O => mac_control_txf_cnt_12_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_28_1242 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_12_LOGIC_ZERO,
      IB => mac_control_txf_cnt_12_CYINIT,
      SEL => mac_control_txf_cnt_12_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_12_CYINIT,
      I1 => mac_control_txf_cnt_12_FROM,
      O => mac_control_txf_cnt_n0000(12)
    );
  mac_control_txf_cnt_12_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(12),
      O => mac_control_txf_cnt_12_FROM
    );
  mac_control_txf_cnt_12_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(13),
      O => mac_control_txf_cnt_12_GROM
    );
  mac_control_txf_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_12_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_29_1243 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_12_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_txf_cnt_12_GROM,
      O => mac_control_txf_cnt_12_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_txf_cnt_12_GROM,
      O => mac_control_txf_cnt_n0000(13)
    );
  mac_control_txf_cnt_12_CYINIT_1244 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_txf_cnt_12_CYINIT
    );
  tx_output_cs_FFd4_1_1245 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd4_GROM,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd4_FFY_RST,
      O => tx_output_cs_FFd4_1
    );
  tx_output_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd4_FFY_RST
    );
  mac_control_txf_cnt_14_LOGIC_ZERO_1246 : X_ZERO
    port map (
      O => mac_control_txf_cnt_14_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_30_1247 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_14_LOGIC_ZERO,
      IB => mac_control_txf_cnt_14_CYINIT,
      SEL => mac_control_txf_cnt_14_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_14_CYINIT,
      I1 => mac_control_txf_cnt_14_FROM,
      O => mac_control_txf_cnt_n0000(14)
    );
  mac_control_txf_cnt_14_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(14),
      O => mac_control_txf_cnt_14_FROM
    );
  mac_control_txf_cnt_14_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(15),
      O => mac_control_txf_cnt_14_GROM
    );
  mac_control_txf_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_14_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_31_1248 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_14_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_txf_cnt_14_GROM,
      O => mac_control_txf_cnt_14_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_txf_cnt_14_GROM,
      O => mac_control_txf_cnt_n0000(15)
    );
  mac_control_txf_cnt_14_CYINIT_1249 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_txf_cnt_14_CYINIT
    );
  mac_control_txf_cnt_16_LOGIC_ZERO_1250 : X_ZERO
    port map (
      O => mac_control_txf_cnt_16_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_32_1251 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_16_LOGIC_ZERO,
      IB => mac_control_txf_cnt_16_CYINIT,
      SEL => mac_control_txf_cnt_16_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_16_CYINIT,
      I1 => mac_control_txf_cnt_16_FROM,
      O => mac_control_txf_cnt_n0000(16)
    );
  mac_control_txf_cnt_16_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(16),
      O => mac_control_txf_cnt_16_FROM
    );
  mac_control_txf_cnt_16_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(17),
      O => mac_control_txf_cnt_16_GROM
    );
  mac_control_txf_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_16_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_33_1252 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_16_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_txf_cnt_16_GROM,
      O => mac_control_txf_cnt_16_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_txf_cnt_16_GROM,
      O => mac_control_txf_cnt_n0000(17)
    );
  mac_control_txf_cnt_16_CYINIT_1253 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_txf_cnt_16_CYINIT
    );
  mac_control_txf_cnt_18_LOGIC_ZERO_1254 : X_ZERO
    port map (
      O => mac_control_txf_cnt_18_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_34_1255 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_18_LOGIC_ZERO,
      IB => mac_control_txf_cnt_18_CYINIT,
      SEL => mac_control_txf_cnt_18_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_18_CYINIT,
      I1 => mac_control_txf_cnt_18_FROM,
      O => mac_control_txf_cnt_n0000(18)
    );
  mac_control_txf_cnt_18_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(18),
      O => mac_control_txf_cnt_18_FROM
    );
  mac_control_txf_cnt_18_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(19),
      O => mac_control_txf_cnt_18_GROM
    );
  mac_control_txf_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_18_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_35_1256 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_18_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_txf_cnt_18_GROM,
      O => mac_control_txf_cnt_18_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_txf_cnt_18_GROM,
      O => mac_control_txf_cnt_n0000(19)
    );
  mac_control_txf_cnt_18_CYINIT_1257 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_txf_cnt_18_CYINIT
    );
  mac_control_txf_cnt_20_LOGIC_ZERO_1258 : X_ZERO
    port map (
      O => mac_control_txf_cnt_20_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_36_1259 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_20_LOGIC_ZERO,
      IB => mac_control_txf_cnt_20_CYINIT,
      SEL => mac_control_txf_cnt_20_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_20_CYINIT,
      I1 => mac_control_txf_cnt_20_FROM,
      O => mac_control_txf_cnt_n0000(20)
    );
  mac_control_txf_cnt_20_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(20),
      O => mac_control_txf_cnt_20_FROM
    );
  mac_control_txf_cnt_20_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(21),
      O => mac_control_txf_cnt_20_GROM
    );
  mac_control_txf_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_20_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_37_1260 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_20_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_txf_cnt_20_GROM,
      O => mac_control_txf_cnt_20_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_txf_cnt_20_GROM,
      O => mac_control_txf_cnt_n0000(21)
    );
  mac_control_txf_cnt_20_CYINIT_1261 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_txf_cnt_20_CYINIT
    );
  mac_control_txf_cnt_22_LOGIC_ZERO_1262 : X_ZERO
    port map (
      O => mac_control_txf_cnt_22_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_38_1263 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_22_LOGIC_ZERO,
      IB => mac_control_txf_cnt_22_CYINIT,
      SEL => mac_control_txf_cnt_22_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_22_CYINIT,
      I1 => mac_control_txf_cnt_22_FROM,
      O => mac_control_txf_cnt_n0000(22)
    );
  mac_control_txf_cnt_22_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_txf_cnt(22),
      ADR3 => VCC,
      O => mac_control_txf_cnt_22_FROM
    );
  mac_control_txf_cnt_22_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(23),
      O => mac_control_txf_cnt_22_GROM
    );
  mac_control_txf_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_22_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_39_1264 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_22_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_txf_cnt_22_GROM,
      O => mac_control_txf_cnt_22_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_txf_cnt_22_GROM,
      O => mac_control_txf_cnt_n0000(23)
    );
  mac_control_txf_cnt_22_CYINIT_1265 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_txf_cnt_22_CYINIT
    );
  mac_control_txf_cnt_24_LOGIC_ZERO_1266 : X_ZERO
    port map (
      O => mac_control_txf_cnt_24_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_40_1267 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_24_LOGIC_ZERO,
      IB => mac_control_txf_cnt_24_CYINIT,
      SEL => mac_control_txf_cnt_24_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_24_CYINIT,
      I1 => mac_control_txf_cnt_24_FROM,
      O => mac_control_txf_cnt_n0000(24)
    );
  mac_control_txf_cnt_24_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(24),
      O => mac_control_txf_cnt_24_FROM
    );
  mac_control_txf_cnt_24_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(25),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_24_GROM
    );
  mac_control_txf_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_24_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_41_1268 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_24_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_txf_cnt_24_GROM,
      O => mac_control_txf_cnt_24_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_txf_cnt_24_GROM,
      O => mac_control_txf_cnt_n0000(25)
    );
  mac_control_txf_cnt_24_CYINIT_1269 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_txf_cnt_24_CYINIT
    );
  mac_control_txf_cnt_26_LOGIC_ZERO_1270 : X_ZERO
    port map (
      O => mac_control_txf_cnt_26_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_42_1271 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_26_LOGIC_ZERO,
      IB => mac_control_txf_cnt_26_CYINIT,
      SEL => mac_control_txf_cnt_26_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_26_CYINIT,
      I1 => mac_control_txf_cnt_26_FROM,
      O => mac_control_txf_cnt_n0000(26)
    );
  mac_control_txf_cnt_26_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(26),
      O => mac_control_txf_cnt_26_FROM
    );
  mac_control_txf_cnt_26_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(27),
      O => mac_control_txf_cnt_26_GROM
    );
  mac_control_txf_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_26_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_43_1272 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_26_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_txf_cnt_26_GROM,
      O => mac_control_txf_cnt_26_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_txf_cnt_26_GROM,
      O => mac_control_txf_cnt_n0000(27)
    );
  mac_control_txf_cnt_26_CYINIT_1273 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_txf_cnt_26_CYINIT
    );
  mac_control_txf_cnt_28_LOGIC_ZERO_1274 : X_ZERO
    port map (
      O => mac_control_txf_cnt_28_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_44_1275 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_28_LOGIC_ZERO,
      IB => mac_control_txf_cnt_28_CYINIT,
      SEL => mac_control_txf_cnt_28_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_28_CYINIT,
      I1 => mac_control_txf_cnt_28_FROM,
      O => mac_control_txf_cnt_n0000(28)
    );
  mac_control_txf_cnt_28_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(28),
      O => mac_control_txf_cnt_28_FROM
    );
  mac_control_txf_cnt_28_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_txf_cnt(29),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_txf_cnt_28_GROM
    );
  mac_control_txf_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_txf_cnt_28_CYMUXG,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_45_1276 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_28_LOGIC_ZERO,
      IB => mac_control_txf_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_txf_cnt_28_GROM,
      O => mac_control_txf_cnt_28_CYMUXG
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_txf_cnt_28_GROM,
      O => mac_control_txf_cnt_n0000(29)
    );
  mac_control_txf_cnt_28_CYINIT_1277 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_txf_cnt_28_CYINIT
    );
  mac_control_txf_cnt_30_LOGIC_ZERO_1278 : X_ZERO
    port map (
      O => mac_control_txf_cnt_30_LOGIC_ZERO
    );
  mac_control_txf_cnt_Madd_n0000_inst_cy_46_1279 : X_MUX2
    port map (
      IA => mac_control_txf_cnt_30_LOGIC_ZERO,
      IB => mac_control_txf_cnt_30_CYINIT,
      SEL => mac_control_txf_cnt_30_FROM,
      O => mac_control_txf_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_30_CYINIT,
      I1 => mac_control_txf_cnt_30_FROM,
      O => mac_control_txf_cnt_n0000(30)
    );
  mac_control_txf_cnt_30_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(30),
      O => mac_control_txf_cnt_30_FROM
    );
  mac_control_txf_cnt_31_rt_1280 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_txf_cnt(31),
      O => mac_control_txf_cnt_31_rt
    );
  mac_control_txf_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_txf_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_txf_cnt_31_rt,
      O => mac_control_txf_cnt_n0000(31)
    );
  mac_control_txf_cnt_30_CYINIT_1281 : X_BUF
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_txf_cnt_30_CYINIT
    );
  addr3ext_0_LOGIC_ZERO_1282 : X_ZERO
    port map (
      O => addr3ext_0_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_101_1283 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_7,
      IB => addr3ext_0_LOGIC_ZERO,
      SEL => rx_output_cs_FFd19_rt,
      O => rx_output_macnt_inst_cy_101
    );
  rx_output_cs_FFd19_rt_1284 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_7,
      ADR1 => VCC,
      ADR2 => rx_output_cs_FFd19,
      ADR3 => VCC,
      O => rx_output_cs_FFd19_rt
    );
  rx_output_macnt_inst_lut3_01 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_14,
      ADR1 => rx_output_bp(0),
      ADR2 => rx_output_cs_FFd19,
      ADR3 => addr3ext(0),
      O => rx_output_macnt_inst_lut3_0
    );
  addr3ext_0_COUTUSED : X_BUF
    port map (
      I => addr3ext_0_CYMUXG,
      O => rx_output_macnt_inst_cy_102
    );
  rx_output_macnt_inst_cy_102_1285 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_14,
      IB => rx_output_macnt_inst_cy_101,
      SEL => rx_output_macnt_inst_lut3_0,
      O => addr3ext_0_CYMUXG
    );
  rx_output_macnt_inst_sum_95_1286 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_101,
      I1 => rx_output_macnt_inst_lut3_0,
      O => rx_output_macnt_inst_sum_95
    );
  addr3ext_1_LOGIC_ZERO_1287 : X_ZERO
    port map (
      O => addr3ext_1_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_103_1288 : X_MUX2
    port map (
      IA => addr3ext_1_LOGIC_ZERO,
      IB => addr3ext_1_CYINIT,
      SEL => rx_output_macnt_inst_lut3_1,
      O => rx_output_macnt_inst_cy_103
    );
  rx_output_macnt_inst_sum_96_1289 : X_XOR2
    port map (
      I0 => addr3ext_1_CYINIT,
      I1 => rx_output_macnt_inst_lut3_1,
      O => rx_output_macnt_inst_sum_96
    );
  rx_output_macnt_inst_lut3_16 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => VCC,
      ADR2 => rx_output_bp(1),
      ADR3 => addr3ext(1),
      O => rx_output_macnt_inst_lut3_1
    );
  rx_output_macnt_inst_lut3_21 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => addr3ext(2),
      ADR2 => rx_output_bp(2),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_2
    );
  addr3ext_1_COUTUSED : X_BUF
    port map (
      I => addr3ext_1_CYMUXG,
      O => rx_output_macnt_inst_cy_104
    );
  rx_output_macnt_inst_cy_104_1290 : X_MUX2
    port map (
      IA => addr3ext_1_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_103,
      SEL => rx_output_macnt_inst_lut3_2,
      O => addr3ext_1_CYMUXG
    );
  rx_output_macnt_inst_sum_97_1291 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_103,
      I1 => rx_output_macnt_inst_lut3_2,
      O => rx_output_macnt_inst_sum_97
    );
  addr3ext_1_CYINIT_1292 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_102,
      O => addr3ext_1_CYINIT
    );
  rx_input_fifo_control_DATA_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(4),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_4_FFY_RST,
      O => rx_input_data(4)
    );
  rx_input_data_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_4_FFY_RST
    );
  addr3ext_3_LOGIC_ZERO_1293 : X_ZERO
    port map (
      O => addr3ext_3_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_105_1294 : X_MUX2
    port map (
      IA => addr3ext_3_LOGIC_ZERO,
      IB => addr3ext_3_CYINIT,
      SEL => rx_output_macnt_inst_lut3_3,
      O => rx_output_macnt_inst_cy_105
    );
  rx_output_macnt_inst_sum_98_1295 : X_XOR2
    port map (
      I0 => addr3ext_3_CYINIT,
      I1 => rx_output_macnt_inst_lut3_3,
      O => rx_output_macnt_inst_sum_98
    );
  rx_output_macnt_inst_lut3_31 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_output_cs_FFd19,
      ADR1 => VCC,
      ADR2 => rx_output_bp(3),
      ADR3 => addr3ext(3),
      O => rx_output_macnt_inst_lut3_3
    );
  rx_output_macnt_inst_lut3_41 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => addr3ext(4),
      ADR1 => VCC,
      ADR2 => rx_output_bp(4),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_4
    );
  addr3ext_3_COUTUSED : X_BUF
    port map (
      I => addr3ext_3_CYMUXG,
      O => rx_output_macnt_inst_cy_106
    );
  rx_output_macnt_inst_cy_106_1296 : X_MUX2
    port map (
      IA => addr3ext_3_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_105,
      SEL => rx_output_macnt_inst_lut3_4,
      O => addr3ext_3_CYMUXG
    );
  rx_output_macnt_inst_sum_99_1297 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_105,
      I1 => rx_output_macnt_inst_lut3_4,
      O => rx_output_macnt_inst_sum_99
    );
  addr3ext_3_CYINIT_1298 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_104,
      O => addr3ext_3_CYINIT
    );
  addr3ext_5_LOGIC_ZERO_1299 : X_ZERO
    port map (
      O => addr3ext_5_LOGIC_ZERO
    );
  rx_output_macnt_inst_cy_107_1300 : X_MUX2
    port map (
      IA => addr3ext_5_LOGIC_ZERO,
      IB => addr3ext_5_CYINIT,
      SEL => rx_output_macnt_inst_lut3_5,
      O => rx_output_macnt_inst_cy_107
    );
  rx_output_macnt_inst_sum_100_1301 : X_XOR2
    port map (
      I0 => addr3ext_5_CYINIT,
      I1 => rx_output_macnt_inst_lut3_5,
      O => rx_output_macnt_inst_sum_100
    );
  rx_output_macnt_inst_lut3_51 : X_LUT4
    generic map(
      INIT => X"F3C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_cs_FFd19,
      ADR2 => rx_output_bp(5),
      ADR3 => addr3ext(5),
      O => rx_output_macnt_inst_lut3_5
    );
  rx_output_macnt_inst_lut3_61 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_bp(6),
      ADR2 => addr3ext(6),
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_macnt_inst_lut3_6
    );
  addr3ext_5_COUTUSED : X_BUF
    port map (
      I => addr3ext_5_CYMUXG,
      O => rx_output_macnt_inst_cy_108
    );
  rx_output_macnt_inst_cy_108_1302 : X_MUX2
    port map (
      IA => addr3ext_5_LOGIC_ZERO,
      IB => rx_output_macnt_inst_cy_107,
      SEL => rx_output_macnt_inst_lut3_6,
      O => addr3ext_5_CYMUXG
    );
  rx_output_macnt_inst_sum_101_1303 : X_XOR2
    port map (
      I0 => rx_output_macnt_inst_cy_107,
      I1 => rx_output_macnt_inst_lut3_6,
      O => rx_output_macnt_inst_sum_101
    );
  addr3ext_5_CYINIT_1304 : X_BUF
    port map (
      I => rx_output_macnt_inst_cy_106,
      O => addr3ext_5_CYINIT
    );
  tx_output_data_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(0),
      CE => tx_output_data_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_0_FFY_RST,
      O => tx_output_data(0)
    );
  tx_output_data_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_0_FFY_RST
    );
  rx_input_memio_macnt_75_LOGIC_ZERO_1305 : X_ZERO
    port map (
      O => rx_input_memio_macnt_75_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_259_1306 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_75_LOGIC_ZERO,
      IB => rx_input_memio_macnt_75_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_61,
      O => rx_input_memio_macnt_inst_cy_259
    );
  rx_input_memio_macnt_inst_sum_224_1307 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_75_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_61,
      O => rx_input_memio_macnt_inst_sum_224
    );
  rx_input_memio_macnt_inst_lut3_611 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => rx_input_memio_bp(5),
      ADR1 => rx_input_memio_macnt_75,
      ADR2 => rx_input_memio_cs_FFd16_2,
      ADR3 => VCC,
      O => rx_input_memio_macnt_inst_lut3_61
    );
  rx_input_memio_macnt_inst_lut3_621 : X_LUT4
    generic map(
      INIT => X"B8B8"
    )
    port map (
      ADR0 => rx_input_memio_bp(6),
      ADR1 => rx_input_memio_cs_FFd16_2,
      ADR2 => rx_input_memio_macnt_76,
      ADR3 => VCC,
      O => rx_input_memio_macnt_inst_lut3_62
    );
  rx_input_memio_macnt_75_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_75_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_260
    );
  rx_input_memio_macnt_inst_cy_260_1308 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_75_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_259,
      SEL => rx_input_memio_macnt_inst_lut3_62,
      O => rx_input_memio_macnt_75_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_225_1309 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_259,
      I1 => rx_input_memio_macnt_inst_lut3_62,
      O => rx_input_memio_macnt_inst_sum_225
    );
  rx_input_memio_macnt_75_CYINIT_1310 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_258,
      O => rx_input_memio_macnt_75_CYINIT
    );
  rx_input_memio_macnt_77_LOGIC_ZERO_1311 : X_ZERO
    port map (
      O => rx_input_memio_macnt_77_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_261_1312 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_77_LOGIC_ZERO,
      IB => rx_input_memio_macnt_77_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_63,
      O => rx_input_memio_macnt_inst_cy_261
    );
  rx_input_memio_macnt_inst_sum_226_1313 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_77_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_63,
      O => rx_input_memio_macnt_inst_sum_226
    );
  rx_input_memio_macnt_inst_lut3_631 : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_macnt_77,
      ADR2 => rx_input_memio_cs_FFd16_2,
      ADR3 => rx_input_memio_bp(7),
      O => rx_input_memio_macnt_inst_lut3_63
    );
  rx_input_memio_macnt_inst_lut3_641 : X_LUT4
    generic map(
      INIT => X"B8B8"
    )
    port map (
      ADR0 => rx_input_memio_bp(8),
      ADR1 => rx_input_memio_cs_FFd16_2,
      ADR2 => rx_input_memio_macnt_78,
      ADR3 => VCC,
      O => rx_input_memio_macnt_inst_lut3_64
    );
  rx_input_memio_macnt_77_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_77_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_262
    );
  rx_input_memio_macnt_inst_cy_262_1314 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_77_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_261,
      SEL => rx_input_memio_macnt_inst_lut3_64,
      O => rx_input_memio_macnt_77_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_227_1315 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_261,
      I1 => rx_input_memio_macnt_inst_lut3_64,
      O => rx_input_memio_macnt_inst_sum_227
    );
  rx_input_memio_macnt_77_CYINIT_1316 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_260,
      O => rx_input_memio_macnt_77_CYINIT
    );
  rx_input_memio_macnt_79_LOGIC_ZERO_1317 : X_ZERO
    port map (
      O => rx_input_memio_macnt_79_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_263_1318 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_79_LOGIC_ZERO,
      IB => rx_input_memio_macnt_79_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_65,
      O => rx_input_memio_macnt_inst_cy_263
    );
  rx_input_memio_macnt_inst_sum_228_1319 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_79_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_65,
      O => rx_input_memio_macnt_inst_sum_228
    );
  rx_input_memio_macnt_inst_lut3_651 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => rx_input_memio_macnt_79,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bp(9),
      ADR3 => rx_input_memio_cs_FFd16_2,
      O => rx_input_memio_macnt_inst_lut3_65
    );
  rx_input_memio_macnt_inst_lut3_661 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bp(10),
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_80,
      ADR3 => rx_input_memio_cs_FFd16_2,
      O => rx_input_memio_macnt_inst_lut3_66
    );
  rx_input_memio_macnt_79_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_79_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_264
    );
  rx_input_memio_macnt_inst_cy_264_1320 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_79_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_263,
      SEL => rx_input_memio_macnt_inst_lut3_66,
      O => rx_input_memio_macnt_79_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_229_1321 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_263,
      I1 => rx_input_memio_macnt_inst_lut3_66,
      O => rx_input_memio_macnt_inst_sum_229
    );
  rx_input_memio_macnt_79_CYINIT_1322 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_262,
      O => rx_input_memio_macnt_79_CYINIT
    );
  rx_input_memio_macnt_81_LOGIC_ZERO_1323 : X_ZERO
    port map (
      O => rx_input_memio_macnt_81_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_265_1324 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_81_LOGIC_ZERO,
      IB => rx_input_memio_macnt_81_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_67,
      O => rx_input_memio_macnt_inst_cy_265
    );
  rx_input_memio_macnt_inst_sum_230_1325 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_81_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_67,
      O => rx_input_memio_macnt_inst_sum_230
    );
  rx_input_memio_macnt_inst_lut3_671 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16_2,
      ADR1 => rx_input_memio_macnt_81,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bp(11),
      O => rx_input_memio_macnt_inst_lut3_67
    );
  rx_input_memio_macnt_inst_lut3_681 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bp(12),
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_82,
      ADR3 => rx_input_memio_cs_FFd16_2,
      O => rx_input_memio_macnt_inst_lut3_68
    );
  rx_input_memio_macnt_81_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_81_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_266
    );
  rx_input_memio_macnt_inst_cy_266_1326 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_81_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_265,
      SEL => rx_input_memio_macnt_inst_lut3_68,
      O => rx_input_memio_macnt_81_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_231_1327 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_265,
      I1 => rx_input_memio_macnt_inst_lut3_68,
      O => rx_input_memio_macnt_inst_sum_231
    );
  rx_input_memio_macnt_81_CYINIT_1328 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_264,
      O => rx_input_memio_macnt_81_CYINIT
    );
  rx_input_memio_macnt_83_LOGIC_ZERO_1329 : X_ZERO
    port map (
      O => rx_input_memio_macnt_83_LOGIC_ZERO
    );
  rx_input_memio_macnt_inst_cy_267_1330 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_83_LOGIC_ZERO,
      IB => rx_input_memio_macnt_83_CYINIT,
      SEL => rx_input_memio_macnt_inst_lut3_69,
      O => rx_input_memio_macnt_inst_cy_267
    );
  rx_input_memio_macnt_inst_sum_232_1331 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_83_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_69,
      O => rx_input_memio_macnt_inst_sum_232
    );
  rx_input_memio_macnt_inst_lut3_691 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => rx_input_memio_bp(13),
      ADR1 => rx_input_memio_macnt_83,
      ADR2 => rx_input_memio_cs_FFd16_2,
      ADR3 => VCC,
      O => rx_input_memio_macnt_inst_lut3_69
    );
  rx_input_memio_macnt_inst_lut3_701 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_cs_FFd16_2,
      ADR2 => rx_input_memio_macnt_84,
      ADR3 => rx_input_memio_bp(14),
      O => rx_input_memio_macnt_inst_lut3_70
    );
  rx_input_memio_macnt_83_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_macnt_83_CYMUXG,
      O => rx_input_memio_macnt_inst_cy_268
    );
  rx_input_memio_macnt_inst_cy_268_1332 : X_MUX2
    port map (
      IA => rx_input_memio_macnt_83_LOGIC_ZERO,
      IB => rx_input_memio_macnt_inst_cy_267,
      SEL => rx_input_memio_macnt_inst_lut3_70,
      O => rx_input_memio_macnt_83_CYMUXG
    );
  rx_input_memio_macnt_inst_sum_233_1333 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_inst_cy_267,
      I1 => rx_input_memio_macnt_inst_lut3_70,
      O => rx_input_memio_macnt_inst_sum_233
    );
  rx_input_memio_macnt_83_CYINIT_1334 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_266,
      O => rx_input_memio_macnt_83_CYINIT
    );
  rx_input_memio_macnt_inst_sum_234_1335 : X_XOR2
    port map (
      I0 => rx_input_memio_macnt_85_CYINIT,
      I1 => rx_input_memio_macnt_inst_lut3_71,
      O => rx_input_memio_macnt_inst_sum_234
    );
  rx_input_memio_macnt_inst_lut3_711 : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_macnt_85,
      ADR2 => rx_input_memio_cs_FFd16_2,
      ADR3 => rx_input_memio_bp(15),
      O => rx_input_memio_macnt_inst_lut3_71
    );
  rx_input_memio_macnt_85_CYINIT_1336 : X_BUF
    port map (
      I => rx_input_memio_macnt_inst_cy_268,
      O => rx_input_memio_macnt_85_CYINIT
    );
  rx_output_n0070_2_LOGIC_ZERO_1337 : X_ZERO
    port map (
      O => rx_output_n0070_2_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_63_1338 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_19,
      IB => rx_output_n0070_2_LOGIC_ZERO,
      SEL => rx_output_Madd_n0047_inst_lut2_641_O,
      O => rx_output_Madd_n0047_inst_cy_63
    );
  rx_output_Madd_n0047_inst_lut2_641 : X_LUT4
    generic map(
      INIT => X"0F0F"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_19,
      ADR1 => VCC,
      ADR2 => rx_output_len(1),
      ADR3 => VCC,
      O => rx_output_Madd_n0047_inst_lut2_641_O
    );
  rx_output_n0070_2_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_28,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(2),
      O => rx_output_n0070_2_GROM
    );
  rx_output_n0070_2_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_2_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_64
    );
  rx_output_n0070_2_YUSED : X_BUF
    port map (
      I => rx_output_n0070_2_XORG,
      O => rx_output_n0070(2)
    );
  rx_output_Madd_n0047_inst_cy_64_1339 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_28,
      IB => rx_output_Madd_n0047_inst_cy_63,
      SEL => rx_output_n0070_2_GROM,
      O => rx_output_n0070_2_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_65 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_63,
      I1 => rx_output_n0070_2_GROM,
      O => rx_output_n0070_2_XORG
    );
  rx_output_n0070_3_LOGIC_ZERO_1340 : X_ZERO
    port map (
      O => rx_output_n0070_3_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_65_1341 : X_MUX2
    port map (
      IA => rx_output_n0070_3_LOGIC_ZERO,
      IB => rx_output_n0070_3_CYINIT,
      SEL => rx_output_n0070_3_FROM,
      O => rx_output_Madd_n0047_inst_cy_65
    );
  rx_output_Madd_n0047_inst_sum_66 : X_XOR2
    port map (
      I0 => rx_output_n0070_3_CYINIT,
      I1 => rx_output_n0070_3_FROM,
      O => rx_output_n0070_3_XORF
    );
  rx_output_n0070_3_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_len(3),
      O => rx_output_n0070_3_FROM
    );
  rx_output_n0070_3_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(4),
      ADR3 => VCC,
      O => rx_output_n0070_3_GROM
    );
  rx_output_n0070_3_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_3_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_66
    );
  rx_output_n0070_3_XUSED : X_BUF
    port map (
      I => rx_output_n0070_3_XORF,
      O => rx_output_n0070(3)
    );
  rx_output_n0070_3_YUSED : X_BUF
    port map (
      I => rx_output_n0070_3_XORG,
      O => rx_output_n0070(4)
    );
  rx_output_Madd_n0047_inst_cy_66_1342 : X_MUX2
    port map (
      IA => rx_output_n0070_3_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_65,
      SEL => rx_output_n0070_3_GROM,
      O => rx_output_n0070_3_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_67 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_65,
      I1 => rx_output_n0070_3_GROM,
      O => rx_output_n0070_3_XORG
    );
  rx_output_n0070_3_CYINIT_1343 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_64,
      O => rx_output_n0070_3_CYINIT
    );
  rx_output_n0070_5_LOGIC_ZERO_1344 : X_ZERO
    port map (
      O => rx_output_n0070_5_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_67_1345 : X_MUX2
    port map (
      IA => rx_output_n0070_5_LOGIC_ZERO,
      IB => rx_output_n0070_5_CYINIT,
      SEL => rx_output_n0070_5_FROM,
      O => rx_output_Madd_n0047_inst_cy_67
    );
  rx_output_Madd_n0047_inst_sum_68 : X_XOR2
    port map (
      I0 => rx_output_n0070_5_CYINIT,
      I1 => rx_output_n0070_5_FROM,
      O => rx_output_n0070_5_XORF
    );
  rx_output_n0070_5_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_5_FROM
    );
  rx_output_n0070_5_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(6),
      ADR3 => VCC,
      O => rx_output_n0070_5_GROM
    );
  rx_output_n0070_5_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_5_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_68
    );
  rx_output_n0070_5_XUSED : X_BUF
    port map (
      I => rx_output_n0070_5_XORF,
      O => rx_output_n0070(5)
    );
  rx_output_n0070_5_YUSED : X_BUF
    port map (
      I => rx_output_n0070_5_XORG,
      O => rx_output_n0070(6)
    );
  rx_output_Madd_n0047_inst_cy_68_1346 : X_MUX2
    port map (
      IA => rx_output_n0070_5_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_67,
      SEL => rx_output_n0070_5_GROM,
      O => rx_output_n0070_5_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_69 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_67,
      I1 => rx_output_n0070_5_GROM,
      O => rx_output_n0070_5_XORG
    );
  rx_output_n0070_5_CYINIT_1347 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_66,
      O => rx_output_n0070_5_CYINIT
    );
  rx_output_n0070_7_LOGIC_ZERO_1348 : X_ZERO
    port map (
      O => rx_output_n0070_7_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_69_1349 : X_MUX2
    port map (
      IA => rx_output_n0070_7_LOGIC_ZERO,
      IB => rx_output_n0070_7_CYINIT,
      SEL => rx_output_n0070_7_FROM,
      O => rx_output_Madd_n0047_inst_cy_69
    );
  rx_output_Madd_n0047_inst_sum_70 : X_XOR2
    port map (
      I0 => rx_output_n0070_7_CYINIT,
      I1 => rx_output_n0070_7_FROM,
      O => rx_output_n0070_7_XORF
    );
  rx_output_n0070_7_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_7_FROM
    );
  rx_output_n0070_7_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(8),
      ADR3 => VCC,
      O => rx_output_n0070_7_GROM
    );
  rx_output_n0070_7_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_7_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_70
    );
  rx_output_n0070_7_XUSED : X_BUF
    port map (
      I => rx_output_n0070_7_XORF,
      O => rx_output_n0070(7)
    );
  rx_output_n0070_7_YUSED : X_BUF
    port map (
      I => rx_output_n0070_7_XORG,
      O => rx_output_n0070(8)
    );
  rx_output_Madd_n0047_inst_cy_70_1350 : X_MUX2
    port map (
      IA => rx_output_n0070_7_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_69,
      SEL => rx_output_n0070_7_GROM,
      O => rx_output_n0070_7_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_71 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_69,
      I1 => rx_output_n0070_7_GROM,
      O => rx_output_n0070_7_XORG
    );
  rx_output_n0070_7_CYINIT_1351 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_68,
      O => rx_output_n0070_7_CYINIT
    );
  rx_output_n0070_9_LOGIC_ZERO_1352 : X_ZERO
    port map (
      O => rx_output_n0070_9_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_71_1353 : X_MUX2
    port map (
      IA => rx_output_n0070_9_LOGIC_ZERO,
      IB => rx_output_n0070_9_CYINIT,
      SEL => rx_output_n0070_9_FROM,
      O => rx_output_Madd_n0047_inst_cy_71
    );
  rx_output_Madd_n0047_inst_sum_72 : X_XOR2
    port map (
      I0 => rx_output_n0070_9_CYINIT,
      I1 => rx_output_n0070_9_FROM,
      O => rx_output_n0070_9_XORF
    );
  rx_output_n0070_9_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_9_FROM
    );
  rx_output_n0070_9_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(10),
      ADR3 => VCC,
      O => rx_output_n0070_9_GROM
    );
  rx_output_n0070_9_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_9_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_72
    );
  rx_output_n0070_9_XUSED : X_BUF
    port map (
      I => rx_output_n0070_9_XORF,
      O => rx_output_n0070(9)
    );
  rx_output_n0070_9_YUSED : X_BUF
    port map (
      I => rx_output_n0070_9_XORG,
      O => rx_output_n0070(10)
    );
  rx_output_Madd_n0047_inst_cy_72_1354 : X_MUX2
    port map (
      IA => rx_output_n0070_9_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_71,
      SEL => rx_output_n0070_9_GROM,
      O => rx_output_n0070_9_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_73 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_71,
      I1 => rx_output_n0070_9_GROM,
      O => rx_output_n0070_9_XORG
    );
  rx_output_n0070_9_CYINIT_1355 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_70,
      O => rx_output_n0070_9_CYINIT
    );
  rx_output_n0070_11_LOGIC_ZERO_1356 : X_ZERO
    port map (
      O => rx_output_n0070_11_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_73_1357 : X_MUX2
    port map (
      IA => rx_output_n0070_11_LOGIC_ZERO,
      IB => rx_output_n0070_11_CYINIT,
      SEL => rx_output_n0070_11_FROM,
      O => rx_output_Madd_n0047_inst_cy_73
    );
  rx_output_Madd_n0047_inst_sum_74 : X_XOR2
    port map (
      I0 => rx_output_n0070_11_CYINIT,
      I1 => rx_output_n0070_11_FROM,
      O => rx_output_n0070_11_XORF
    );
  rx_output_n0070_11_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(11),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_11_FROM
    );
  rx_output_n0070_11_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(12),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_11_GROM
    );
  rx_output_n0070_11_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_11_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_74
    );
  rx_output_n0070_11_XUSED : X_BUF
    port map (
      I => rx_output_n0070_11_XORF,
      O => rx_output_n0070(11)
    );
  rx_output_n0070_11_YUSED : X_BUF
    port map (
      I => rx_output_n0070_11_XORG,
      O => rx_output_n0070(12)
    );
  rx_output_Madd_n0047_inst_cy_74_1358 : X_MUX2
    port map (
      IA => rx_output_n0070_11_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_73,
      SEL => rx_output_n0070_11_GROM,
      O => rx_output_n0070_11_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_75 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_73,
      I1 => rx_output_n0070_11_GROM,
      O => rx_output_n0070_11_XORG
    );
  rx_output_n0070_11_CYINIT_1359 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_72,
      O => rx_output_n0070_11_CYINIT
    );
  rx_output_n0070_13_LOGIC_ZERO_1360 : X_ZERO
    port map (
      O => rx_output_n0070_13_LOGIC_ZERO
    );
  rx_output_Madd_n0047_inst_cy_75_1361 : X_MUX2
    port map (
      IA => rx_output_n0070_13_LOGIC_ZERO,
      IB => rx_output_n0070_13_CYINIT,
      SEL => rx_output_n0070_13_FROM,
      O => rx_output_Madd_n0047_inst_cy_75
    );
  rx_output_Madd_n0047_inst_sum_76 : X_XOR2
    port map (
      I0 => rx_output_n0070_13_CYINIT,
      I1 => rx_output_n0070_13_FROM,
      O => rx_output_n0070_13_XORF
    );
  rx_output_n0070_13_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_len(13),
      ADR3 => VCC,
      O => rx_output_n0070_13_FROM
    );
  rx_output_n0070_13_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_len(14),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_n0070_13_GROM
    );
  rx_output_n0070_13_COUTUSED : X_BUF
    port map (
      I => rx_output_n0070_13_CYMUXG,
      O => rx_output_Madd_n0047_inst_cy_76
    );
  rx_output_n0070_13_XUSED : X_BUF
    port map (
      I => rx_output_n0070_13_XORF,
      O => rx_output_n0070(13)
    );
  rx_output_n0070_13_YUSED : X_BUF
    port map (
      I => rx_output_n0070_13_XORG,
      O => rx_output_n0070(14)
    );
  rx_output_Madd_n0047_inst_cy_76_1362 : X_MUX2
    port map (
      IA => rx_output_n0070_13_LOGIC_ZERO,
      IB => rx_output_Madd_n0047_inst_cy_75,
      SEL => rx_output_n0070_13_GROM,
      O => rx_output_n0070_13_CYMUXG
    );
  rx_output_Madd_n0047_inst_sum_77 : X_XOR2
    port map (
      I0 => rx_output_Madd_n0047_inst_cy_75,
      I1 => rx_output_n0070_13_GROM,
      O => rx_output_n0070_13_XORG
    );
  rx_output_n0070_13_CYINIT_1363 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_74,
      O => rx_output_n0070_13_CYINIT
    );
  rx_output_Madd_n0047_inst_sum_78 : X_XOR2
    port map (
      I0 => rx_output_n0070_15_CYINIT,
      I1 => rx_output_SIG_38,
      O => rx_output_n0070_15_XORF
    );
  rx_output_BEL_19 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(15),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_SIG_38
    );
  rx_output_n0070_15_XUSED : X_BUF
    port map (
      I => rx_output_n0070_15_XORF,
      O => rx_output_n0070(15)
    );
  rx_output_n0070_15_CYINIT_1364 : X_BUF
    port map (
      I => rx_output_Madd_n0047_inst_cy_76,
      O => rx_output_n0070_15_CYINIT
    );
  rx_input_fifo_control_DATA_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(7),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_data_7_FFY_RST,
      O => rx_input_data(7)
    );
  rx_input_data_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_data_7_FFY_RST
    );
  tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ONE_1365 : X_ONE
    port map (
      O => tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ONE
    );
  tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ZERO_1366 : X_ZERO
    port map (
      O => tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ZERO
    );
  tx_output_Mcompar_n0006_inst_cy_78_1367 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ONE,
      SEL => tx_output_Mcompar_n0006_inst_lut4_0,
      O => tx_output_Mcompar_n0006_inst_cy_78
    );
  tx_output_Mcompar_n0006_inst_lut4_01 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => txfbbp(0),
      ADR1 => txfbbp(1),
      ADR2 => tx_output_bpl(0),
      ADR3 => tx_output_bpl(1),
      O => tx_output_Mcompar_n0006_inst_lut4_0
    );
  tx_output_Mcompar_n0006_inst_lut4_11 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => txfbbp(3),
      ADR1 => txfbbp(2),
      ADR2 => tx_output_bpl(2),
      ADR3 => tx_output_bpl(3),
      O => tx_output_Mcompar_n0006_inst_lut4_1
    );
  tx_output_Mcompar_n0006_inst_cy_79_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_79_CYMUXG,
      O => tx_output_Mcompar_n0006_inst_cy_79
    );
  tx_output_Mcompar_n0006_inst_cy_79_1368 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_79_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_78,
      SEL => tx_output_Mcompar_n0006_inst_lut4_1,
      O => tx_output_Mcompar_n0006_inst_cy_79_CYMUXG
    );
  tx_output_Mcompar_n0006_inst_cy_81_LOGIC_ZERO_1369 : X_ZERO
    port map (
      O => tx_output_Mcompar_n0006_inst_cy_81_LOGIC_ZERO
    );
  tx_output_Mcompar_n0006_inst_cy_80_1370 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_81_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_81_CYINIT,
      SEL => tx_output_Mcompar_n0006_inst_lut4_2,
      O => tx_output_Mcompar_n0006_inst_cy_80
    );
  tx_output_Mcompar_n0006_inst_lut4_21 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => txfbbp(5),
      ADR1 => tx_output_bpl(4),
      ADR2 => tx_output_bpl(5),
      ADR3 => txfbbp(4),
      O => tx_output_Mcompar_n0006_inst_lut4_2
    );
  tx_output_Mcompar_n0006_inst_lut4_31 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => txfbbp(6),
      ADR1 => txfbbp(7),
      ADR2 => tx_output_bpl(7),
      ADR3 => tx_output_bpl(6),
      O => tx_output_Mcompar_n0006_inst_lut4_3
    );
  tx_output_Mcompar_n0006_inst_cy_81_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_81_CYMUXG,
      O => tx_output_Mcompar_n0006_inst_cy_81
    );
  tx_output_Mcompar_n0006_inst_cy_81_1371 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_81_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_80,
      SEL => tx_output_Mcompar_n0006_inst_lut4_3,
      O => tx_output_Mcompar_n0006_inst_cy_81_CYMUXG
    );
  tx_output_Mcompar_n0006_inst_cy_81_CYINIT_1372 : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_79,
      O => tx_output_Mcompar_n0006_inst_cy_81_CYINIT
    );
  tx_output_Mcompar_n0006_inst_cy_83_LOGIC_ZERO_1373 : X_ZERO
    port map (
      O => tx_output_Mcompar_n0006_inst_cy_83_LOGIC_ZERO
    );
  tx_output_Mcompar_n0006_inst_cy_82_1374 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_83_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_83_CYINIT,
      SEL => tx_output_Mcompar_n0006_inst_lut4_4,
      O => tx_output_Mcompar_n0006_inst_cy_82
    );
  tx_output_Mcompar_n0006_inst_lut4_41 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => txfbbp(9),
      ADR1 => tx_output_bpl(8),
      ADR2 => txfbbp(8),
      ADR3 => tx_output_bpl(9),
      O => tx_output_Mcompar_n0006_inst_lut4_4
    );
  tx_output_Mcompar_n0006_inst_lut4_51 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => txfbbp(10),
      ADR1 => txfbbp(11),
      ADR2 => tx_output_bpl(11),
      ADR3 => tx_output_bpl(10),
      O => tx_output_Mcompar_n0006_inst_lut4_5
    );
  tx_output_Mcompar_n0006_inst_cy_83_COUTUSED : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_83_CYMUXG,
      O => tx_output_Mcompar_n0006_inst_cy_83
    );
  tx_output_Mcompar_n0006_inst_cy_83_1375 : X_MUX2
    port map (
      IA => tx_output_Mcompar_n0006_inst_cy_83_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_82,
      SEL => tx_output_Mcompar_n0006_inst_lut4_5,
      O => tx_output_Mcompar_n0006_inst_cy_83_CYMUXG
    );
  tx_output_Mcompar_n0006_inst_cy_83_CYINIT_1376 : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_81,
      O => tx_output_Mcompar_n0006_inst_cy_83_CYINIT
    );
  tx_output_n0006_LOGIC_ZERO_1377 : X_ZERO
    port map (
      O => tx_output_n0006_LOGIC_ZERO
    );
  tx_output_Mcompar_n0006_inst_cy_84_1378 : X_MUX2
    port map (
      IA => tx_output_n0006_LOGIC_ZERO,
      IB => tx_output_n0006_CYINIT,
      SEL => tx_output_Mcompar_n0006_inst_lut4_6,
      O => tx_output_Mcompar_n0006_inst_cy_84
    );
  tx_output_Mcompar_n0006_inst_lut4_61 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => txfbbp(13),
      ADR1 => tx_output_bpl(13),
      ADR2 => txfbbp(12),
      ADR3 => tx_output_bpl(12),
      O => tx_output_Mcompar_n0006_inst_lut4_6
    );
  tx_output_Mcompar_n0006_inst_lut4_71 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => tx_output_bpl(14),
      ADR1 => tx_output_bpl(15),
      ADR2 => txfbbp(15),
      ADR3 => txfbbp(14),
      O => tx_output_Mcompar_n0006_inst_lut4_7
    );
  tx_output_n0006_COUTUSED : X_BUF
    port map (
      I => tx_output_n0006_CYMUXG,
      O => tx_output_n0006
    );
  tx_output_Mcompar_n0006_inst_cy_85 : X_MUX2
    port map (
      IA => tx_output_n0006_LOGIC_ZERO,
      IB => tx_output_Mcompar_n0006_inst_cy_84,
      SEL => tx_output_Mcompar_n0006_inst_lut4_7,
      O => tx_output_n0006_CYMUXG
    );
  tx_output_n0006_CYINIT_1379 : X_BUF
    port map (
      I => tx_output_Mcompar_n0006_inst_cy_83,
      O => tx_output_n0006_CYINIT
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ONE_1380 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ZERO_1381 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_177_1382 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(40),
      ADR1 => rx_input_memio_addrchk_datal(41),
      ADR2 => rx_input_memio_addrchk_macaddrl(41),
      ADR3 => rx_input_memio_addrchk_macaddrl(40),
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(43),
      ADR1 => rx_input_memio_addrchk_macaddrl(42),
      ADR2 => rx_input_memio_addrchk_datal(42),
      ADR3 => rx_input_memio_addrchk_datal(43),
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_1383 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_0_LOGIC_ZERO_1384 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_0_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_179_1385 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_0_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_0_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(44),
      ADR1 => rx_input_memio_addrchk_macaddrl(45),
      ADR2 => rx_input_memio_addrchk_datal(45),
      ADR3 => rx_input_memio_addrchk_macaddrl(44),
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(47),
      ADR1 => rx_input_memio_addrchk_datal(47),
      ADR2 => rx_input_memio_addrchk_macaddrl(46),
      ADR3 => rx_input_memio_addrchk_datal(46),
      O => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_0_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_0_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(0)
    );
  rx_input_memio_addrchk_Mcompar_n0048_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_0_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0048_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_0_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_0_CYINIT_1386 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0048_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_0_CYINIT
    );
  rx_input_memio_bcntl_0_LOGIC_ONE_1387 : X_ONE
    port map (
      O => rx_input_memio_bcntl_0_LOGIC_ONE
    );
  rx_input_memio_Msub_n0042_inst_cy_237_1388 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_86,
      IB => rx_input_memio_bcntl_0_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_149,
      O => rx_input_memio_Msub_n0042_inst_cy_237
    );
  rx_input_memio_Msub_n0042_inst_sum_203 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_0_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_149,
      O => rx_input_memio_n0042(0)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1491 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_86,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_149
    );
  rx_input_memio_Msub_n0042_inst_lut2_1501 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_87,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_150
    );
  rx_input_memio_bcntl_0_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_0_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_238
    );
  rx_input_memio_Msub_n0042_inst_cy_238_1389 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_87,
      IB => rx_input_memio_Msub_n0042_inst_cy_237,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_150,
      O => rx_input_memio_bcntl_0_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_204 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_237,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_150,
      O => rx_input_memio_n0042(1)
    );
  rx_input_memio_bcntl_0_CYINIT_1390 : X_BUF
    port map (
      I => rx_input_memio_bcntl_0_LOGIC_ONE,
      O => rx_input_memio_bcntl_0_CYINIT
    );
  rx_input_memio_bcntl_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_2_FFY_RST
    );
  rx_input_memio_bcntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(3),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_2_FFY_RST,
      O => rx_input_memio_bcntl(3)
    );
  rx_input_memio_Msub_n0042_inst_cy_239_1391 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_7,
      IB => rx_input_memio_bcntl_2_CYINIT,
      SEL => rx_input_memio_bcntl_2_FROM,
      O => rx_input_memio_Msub_n0042_inst_cy_239
    );
  rx_input_memio_Msub_n0042_inst_sum_205 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_2_CYINIT,
      I1 => rx_input_memio_bcntl_2_FROM,
      O => rx_input_memio_n0042(2)
    );
  rx_input_memio_bcntl_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_7,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bcnt_88,
      O => rx_input_memio_bcntl_2_FROM
    );
  rx_input_memio_Msub_n0042_inst_lut2_1521 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_89,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_152
    );
  rx_input_memio_bcntl_2_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_2_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_240
    );
  rx_input_memio_Msub_n0042_inst_cy_240_1392 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_89,
      IB => rx_input_memio_Msub_n0042_inst_cy_239,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_152,
      O => rx_input_memio_bcntl_2_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_206 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_239,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_152,
      O => rx_input_memio_n0042(3)
    );
  rx_input_memio_bcntl_2_CYINIT_1393 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_238,
      O => rx_input_memio_bcntl_2_CYINIT
    );
  rx_input_memio_bcntl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_4_FFY_RST
    );
  rx_input_memio_bcntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(5),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_4_FFY_RST,
      O => rx_input_memio_bcntl(5)
    );
  rx_input_memio_Msub_n0042_inst_cy_241_1394 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_90,
      IB => rx_input_memio_bcntl_4_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_153,
      O => rx_input_memio_Msub_n0042_inst_cy_241
    );
  rx_input_memio_Msub_n0042_inst_sum_207 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_4_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_153,
      O => rx_input_memio_n0042(4)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1531 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_90,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_153
    );
  rx_input_memio_Msub_n0042_inst_lut2_1541 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_91,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_154
    );
  rx_input_memio_bcntl_4_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_4_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_242
    );
  rx_input_memio_Msub_n0042_inst_cy_242_1395 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_91,
      IB => rx_input_memio_Msub_n0042_inst_cy_241,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_154,
      O => rx_input_memio_bcntl_4_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_208 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_241,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_154,
      O => rx_input_memio_n0042(5)
    );
  rx_input_memio_bcntl_4_CYINIT_1396 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_240,
      O => rx_input_memio_bcntl_4_CYINIT
    );
  rx_input_memio_bcntl_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_6_FFY_RST
    );
  rx_input_memio_bcntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(7),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_6_FFY_RST,
      O => rx_input_memio_bcntl(7)
    );
  rx_input_memio_Msub_n0042_inst_cy_243_1397 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_92,
      IB => rx_input_memio_bcntl_6_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_155,
      O => rx_input_memio_Msub_n0042_inst_cy_243
    );
  rx_input_memio_Msub_n0042_inst_sum_209 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_6_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_155,
      O => rx_input_memio_n0042(6)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1551 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_92,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_155
    );
  rx_input_memio_Msub_n0042_inst_lut2_1561 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_93,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_156
    );
  rx_input_memio_bcntl_6_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_6_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_244
    );
  rx_input_memio_Msub_n0042_inst_cy_244_1398 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_93,
      IB => rx_input_memio_Msub_n0042_inst_cy_243,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_156,
      O => rx_input_memio_bcntl_6_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_210 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_243,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_156,
      O => rx_input_memio_n0042(7)
    );
  rx_input_memio_bcntl_6_CYINIT_1399 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_242,
      O => rx_input_memio_bcntl_6_CYINIT
    );
  rx_input_memio_bcntl_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_8_FFY_RST
    );
  rx_input_memio_bcntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(9),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_8_FFY_RST,
      O => rx_input_memio_bcntl(9)
    );
  rx_input_memio_Msub_n0042_inst_cy_245_1400 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_94,
      IB => rx_input_memio_bcntl_8_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_157,
      O => rx_input_memio_Msub_n0042_inst_cy_245
    );
  rx_input_memio_Msub_n0042_inst_sum_211 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_8_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_157,
      O => rx_input_memio_n0042(8)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1571 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_94,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_157
    );
  rx_input_memio_Msub_n0042_inst_lut2_1581 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_95,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_158
    );
  rx_input_memio_bcntl_8_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_8_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_246
    );
  rx_input_memio_Msub_n0042_inst_cy_246_1401 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_95,
      IB => rx_input_memio_Msub_n0042_inst_cy_245,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_158,
      O => rx_input_memio_bcntl_8_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_212 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_245,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_158,
      O => rx_input_memio_n0042(9)
    );
  rx_input_memio_bcntl_8_CYINIT_1402 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_244,
      O => rx_input_memio_bcntl_8_CYINIT
    );
  rx_input_fifo_control_cs_FFd3_1403 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_cs_FFd3_FFX_RST,
      O => rx_input_fifo_control_cs_FFd3
    );
  rx_input_fifo_control_cs_FFd3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_cs_FFd3_FFX_RST
    );
  rx_input_memio_bcntl_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_10_FFY_RST
    );
  rx_input_memio_bcntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(11),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_10_FFY_RST,
      O => rx_input_memio_bcntl(11)
    );
  rx_input_memio_Msub_n0042_inst_cy_247_1404 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_96,
      IB => rx_input_memio_bcntl_10_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_159,
      O => rx_input_memio_Msub_n0042_inst_cy_247
    );
  rx_input_memio_Msub_n0042_inst_sum_213 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_10_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_159,
      O => rx_input_memio_n0042(10)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1591 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_96,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_159
    );
  rx_input_memio_Msub_n0042_inst_lut2_1601 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_97,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_160
    );
  rx_input_memio_bcntl_10_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_10_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_248
    );
  rx_input_memio_Msub_n0042_inst_cy_248_1405 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_97,
      IB => rx_input_memio_Msub_n0042_inst_cy_247,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_160,
      O => rx_input_memio_bcntl_10_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_214 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_247,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_160,
      O => rx_input_memio_n0042(11)
    );
  rx_input_memio_bcntl_10_CYINIT_1406 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_246,
      O => rx_input_memio_bcntl_10_CYINIT
    );
  rx_input_memio_bcntl_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_12_FFY_RST
    );
  rx_input_memio_bcntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(13),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_12_FFY_RST,
      O => rx_input_memio_bcntl(13)
    );
  rx_input_memio_Msub_n0042_inst_cy_249_1407 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_98,
      IB => rx_input_memio_bcntl_12_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_161,
      O => rx_input_memio_Msub_n0042_inst_cy_249
    );
  rx_input_memio_Msub_n0042_inst_sum_215 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_12_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_161,
      O => rx_input_memio_n0042(12)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1611 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_98,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_161
    );
  rx_input_memio_Msub_n0042_inst_lut2_1621 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_99,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_162
    );
  rx_input_memio_bcntl_12_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_bcntl_12_CYMUXG,
      O => rx_input_memio_Msub_n0042_inst_cy_250
    );
  rx_input_memio_Msub_n0042_inst_cy_250_1408 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_99,
      IB => rx_input_memio_Msub_n0042_inst_cy_249,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_162,
      O => rx_input_memio_bcntl_12_CYMUXG
    );
  rx_input_memio_Msub_n0042_inst_sum_216 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_249,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_162,
      O => rx_input_memio_n0042(13)
    );
  rx_input_memio_bcntl_12_CYINIT_1409 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_248,
      O => rx_input_memio_bcntl_12_CYINIT
    );
  rx_input_memio_bcntl_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_14_FFY_RST
    );
  rx_input_memio_bcntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(15),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_14_FFY_RST,
      O => rx_input_memio_bcntl(15)
    );
  rx_input_memio_Msub_n0042_inst_cy_251_1410 : X_MUX2
    port map (
      IA => rx_input_memio_bcnt_100,
      IB => rx_input_memio_bcntl_14_CYINIT,
      SEL => rx_input_memio_Msub_n0042_inst_lut2_163,
      O => rx_input_memio_Msub_n0042_inst_cy_251
    );
  rx_input_memio_Msub_n0042_inst_sum_217 : X_XOR2
    port map (
      I0 => rx_input_memio_bcntl_14_CYINIT,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_163,
      O => rx_input_memio_n0042(14)
    );
  rx_input_memio_Msub_n0042_inst_lut2_1631 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_100,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_163
    );
  rx_input_memio_Msub_n0042_inst_lut2_1641 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_input_memio_bcnt_101,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_Msub_n0042_inst_lut2_164
    );
  rx_input_memio_Msub_n0042_inst_sum_218 : X_XOR2
    port map (
      I0 => rx_input_memio_Msub_n0042_inst_cy_251,
      I1 => rx_input_memio_Msub_n0042_inst_lut2_164,
      O => rx_input_memio_n0042(15)
    );
  rx_input_memio_bcntl_14_CYINIT_1411 : X_BUF
    port map (
      I => rx_input_memio_Msub_n0042_inst_cy_250,
      O => rx_input_memio_bcntl_14_CYINIT
    );
  tx_input_addr_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_16_FFY_RST
    );
  tx_input_addr_16_1412 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_127,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_16_FFY_RST,
      O => tx_input_addr_16
    );
  tx_input_addr_16_LOGIC_ZERO_1413 : X_ZERO
    port map (
      O => tx_input_addr_16_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_134_1414 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_12,
      IB => tx_input_addr_16_LOGIC_ZERO,
      SEL => tx_input_cs_FFd12_rt,
      O => tx_input_addr_inst_cy_134
    );
  tx_input_cs_FFd12_rt_1415 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_12,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_cs_FFd12_rt
    );
  tx_input_addr_inst_lut3_161 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_19,
      ADR1 => txbp(0),
      ADR2 => tx_input_addr_16,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_addr_inst_lut3_16
    );
  tx_input_addr_16_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_16_CYMUXG,
      O => tx_input_addr_inst_cy_135
    );
  tx_input_addr_inst_cy_135_1416 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_19,
      IB => tx_input_addr_inst_cy_134,
      SEL => tx_input_addr_inst_lut3_16,
      O => tx_input_addr_16_CYMUXG
    );
  tx_input_addr_inst_sum_127_1417 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_134,
      I1 => tx_input_addr_inst_lut3_16,
      O => tx_input_addr_inst_sum_127
    );
  tx_input_addr_17_LOGIC_ZERO_1418 : X_ZERO
    port map (
      O => tx_input_addr_17_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_136_1419 : X_MUX2
    port map (
      IA => tx_input_addr_17_LOGIC_ZERO,
      IB => tx_input_addr_17_CYINIT,
      SEL => tx_input_addr_inst_lut3_17,
      O => tx_input_addr_inst_cy_136
    );
  tx_input_addr_inst_sum_128_1420 : X_XOR2
    port map (
      I0 => tx_input_addr_17_CYINIT,
      I1 => tx_input_addr_inst_lut3_17,
      O => tx_input_addr_inst_sum_128
    );
  tx_input_addr_inst_lut3_171 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => tx_input_addr_17,
      ADR1 => txbp(1),
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_addr_inst_lut3_17
    );
  tx_input_addr_inst_lut3_181 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => VCC,
      ADR2 => tx_input_addr_18,
      ADR3 => txbp(2),
      O => tx_input_addr_inst_lut3_18
    );
  tx_input_addr_17_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_17_CYMUXG,
      O => tx_input_addr_inst_cy_137
    );
  tx_input_addr_inst_cy_137_1421 : X_MUX2
    port map (
      IA => tx_input_addr_17_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_136,
      SEL => tx_input_addr_inst_lut3_18,
      O => tx_input_addr_17_CYMUXG
    );
  tx_input_addr_inst_sum_129_1422 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_136,
      I1 => tx_input_addr_inst_lut3_18,
      O => tx_input_addr_inst_sum_129
    );
  tx_input_addr_17_CYINIT_1423 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_135,
      O => tx_input_addr_17_CYINIT
    );
  tx_input_addr_19_LOGIC_ZERO_1424 : X_ZERO
    port map (
      O => tx_input_addr_19_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_138_1425 : X_MUX2
    port map (
      IA => tx_input_addr_19_LOGIC_ZERO,
      IB => tx_input_addr_19_CYINIT,
      SEL => tx_input_addr_inst_lut3_19,
      O => tx_input_addr_inst_cy_138
    );
  tx_input_addr_inst_sum_130_1426 : X_XOR2
    port map (
      I0 => tx_input_addr_19_CYINIT,
      I1 => tx_input_addr_inst_lut3_19,
      O => tx_input_addr_inst_sum_130
    );
  tx_input_addr_inst_lut3_191 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => tx_input_addr_19,
      ADR3 => txbp(3),
      O => tx_input_addr_inst_lut3_19
    );
  tx_input_addr_inst_lut3_201 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => txbp(4),
      ADR1 => VCC,
      ADR2 => tx_input_addr_20,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_addr_inst_lut3_20
    );
  tx_input_addr_19_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_19_CYMUXG,
      O => tx_input_addr_inst_cy_139
    );
  tx_input_addr_inst_cy_139_1427 : X_MUX2
    port map (
      IA => tx_input_addr_19_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_138,
      SEL => tx_input_addr_inst_lut3_20,
      O => tx_input_addr_19_CYMUXG
    );
  tx_input_addr_inst_sum_131_1428 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_138,
      I1 => tx_input_addr_inst_lut3_20,
      O => tx_input_addr_inst_sum_131
    );
  tx_input_addr_19_CYINIT_1429 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_137,
      O => tx_input_addr_19_CYINIT
    );
  tx_input_addr_21_LOGIC_ZERO_1430 : X_ZERO
    port map (
      O => tx_input_addr_21_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_140_1431 : X_MUX2
    port map (
      IA => tx_input_addr_21_LOGIC_ZERO,
      IB => tx_input_addr_21_CYINIT,
      SEL => tx_input_addr_inst_lut3_21,
      O => tx_input_addr_inst_cy_140
    );
  tx_input_addr_inst_sum_132_1432 : X_XOR2
    port map (
      I0 => tx_input_addr_21_CYINIT,
      I1 => tx_input_addr_inst_lut3_21,
      O => tx_input_addr_inst_sum_132
    );
  tx_input_addr_inst_lut3_211 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => tx_input_addr_21,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => VCC,
      ADR3 => txbp(5),
      O => tx_input_addr_inst_lut3_21
    );
  tx_input_addr_inst_lut3_221 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => txbp(6),
      ADR1 => tx_input_addr_22,
      ADR2 => tx_input_cs_FFd12,
      ADR3 => VCC,
      O => tx_input_addr_inst_lut3_22
    );
  tx_input_addr_21_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_21_CYMUXG,
      O => tx_input_addr_inst_cy_141
    );
  tx_input_addr_inst_cy_141_1433 : X_MUX2
    port map (
      IA => tx_input_addr_21_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_140,
      SEL => tx_input_addr_inst_lut3_22,
      O => tx_input_addr_21_CYMUXG
    );
  tx_input_addr_inst_sum_133_1434 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_140,
      I1 => tx_input_addr_inst_lut3_22,
      O => tx_input_addr_inst_sum_133
    );
  tx_input_addr_21_CYINIT_1435 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_139,
      O => tx_input_addr_21_CYINIT
    );
  tx_input_addr_23_LOGIC_ZERO_1436 : X_ZERO
    port map (
      O => tx_input_addr_23_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_142_1437 : X_MUX2
    port map (
      IA => tx_input_addr_23_LOGIC_ZERO,
      IB => tx_input_addr_23_CYINIT,
      SEL => tx_input_addr_inst_lut3_23,
      O => tx_input_addr_inst_cy_142
    );
  tx_input_addr_inst_sum_134_1438 : X_XOR2
    port map (
      I0 => tx_input_addr_23_CYINIT,
      I1 => tx_input_addr_inst_lut3_23,
      O => tx_input_addr_inst_sum_134
    );
  tx_input_addr_inst_lut3_231 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => tx_input_addr_23,
      ADR2 => VCC,
      ADR3 => txbp(7),
      O => tx_input_addr_inst_lut3_23
    );
  tx_input_addr_inst_lut3_241 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => VCC,
      ADR2 => txbp(8),
      ADR3 => tx_input_addr_24,
      O => tx_input_addr_inst_lut3_24
    );
  tx_input_addr_23_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_23_CYMUXG,
      O => tx_input_addr_inst_cy_143
    );
  tx_input_addr_inst_cy_143_1439 : X_MUX2
    port map (
      IA => tx_input_addr_23_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_142,
      SEL => tx_input_addr_inst_lut3_24,
      O => tx_input_addr_23_CYMUXG
    );
  tx_input_addr_inst_sum_135_1440 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_142,
      I1 => tx_input_addr_inst_lut3_24,
      O => tx_input_addr_inst_sum_135
    );
  tx_input_addr_23_CYINIT_1441 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_141,
      O => tx_input_addr_23_CYINIT
    );
  tx_input_addr_25_LOGIC_ZERO_1442 : X_ZERO
    port map (
      O => tx_input_addr_25_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_144_1443 : X_MUX2
    port map (
      IA => tx_input_addr_25_LOGIC_ZERO,
      IB => tx_input_addr_25_CYINIT,
      SEL => tx_input_addr_inst_lut3_25,
      O => tx_input_addr_inst_cy_144
    );
  tx_input_addr_inst_sum_136_1444 : X_XOR2
    port map (
      I0 => tx_input_addr_25_CYINIT,
      I1 => tx_input_addr_inst_lut3_25,
      O => tx_input_addr_inst_sum_136
    );
  tx_input_addr_inst_lut3_251 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => VCC,
      ADR2 => tx_input_addr_25,
      ADR3 => txbp(9),
      O => tx_input_addr_inst_lut3_25
    );
  tx_input_addr_inst_lut3_261 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => VCC,
      ADR2 => txbp(10),
      ADR3 => tx_input_addr_26,
      O => tx_input_addr_inst_lut3_26
    );
  tx_input_addr_25_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_25_CYMUXG,
      O => tx_input_addr_inst_cy_145
    );
  tx_input_addr_inst_cy_145_1445 : X_MUX2
    port map (
      IA => tx_input_addr_25_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_144,
      SEL => tx_input_addr_inst_lut3_26,
      O => tx_input_addr_25_CYMUXG
    );
  tx_input_addr_inst_sum_137_1446 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_144,
      I1 => tx_input_addr_inst_lut3_26,
      O => tx_input_addr_inst_sum_137
    );
  tx_input_addr_25_CYINIT_1447 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_143,
      O => tx_input_addr_25_CYINIT
    );
  tx_input_addr_27_LOGIC_ZERO_1448 : X_ZERO
    port map (
      O => tx_input_addr_27_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_146_1449 : X_MUX2
    port map (
      IA => tx_input_addr_27_LOGIC_ZERO,
      IB => tx_input_addr_27_CYINIT,
      SEL => tx_input_addr_inst_lut3_27,
      O => tx_input_addr_inst_cy_146
    );
  tx_input_addr_inst_sum_138_1450 : X_XOR2
    port map (
      I0 => tx_input_addr_27_CYINIT,
      I1 => tx_input_addr_inst_lut3_27,
      O => tx_input_addr_inst_sum_138
    );
  tx_input_addr_inst_lut3_271 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => tx_input_addr_27,
      ADR2 => VCC,
      ADR3 => txbp(11),
      O => tx_input_addr_inst_lut3_27
    );
  tx_input_addr_inst_lut3_281 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => VCC,
      ADR2 => tx_input_addr_28,
      ADR3 => txbp(12),
      O => tx_input_addr_inst_lut3_28
    );
  tx_input_addr_27_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_27_CYMUXG,
      O => tx_input_addr_inst_cy_147
    );
  tx_input_addr_inst_cy_147_1451 : X_MUX2
    port map (
      IA => tx_input_addr_27_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_146,
      SEL => tx_input_addr_inst_lut3_28,
      O => tx_input_addr_27_CYMUXG
    );
  tx_input_addr_inst_sum_139_1452 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_146,
      I1 => tx_input_addr_inst_lut3_28,
      O => tx_input_addr_inst_sum_139
    );
  tx_input_addr_27_CYINIT_1453 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_145,
      O => tx_input_addr_27_CYINIT
    );
  tx_input_addr_29_LOGIC_ZERO_1454 : X_ZERO
    port map (
      O => tx_input_addr_29_LOGIC_ZERO
    );
  tx_input_addr_inst_cy_148_1455 : X_MUX2
    port map (
      IA => tx_input_addr_29_LOGIC_ZERO,
      IB => tx_input_addr_29_CYINIT,
      SEL => tx_input_addr_inst_lut3_29,
      O => tx_input_addr_inst_cy_148
    );
  tx_input_addr_inst_sum_140_1456 : X_XOR2
    port map (
      I0 => tx_input_addr_29_CYINIT,
      I1 => tx_input_addr_inst_lut3_29,
      O => tx_input_addr_inst_sum_140
    );
  tx_input_addr_inst_lut3_291 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => tx_input_addr_29,
      ADR2 => txbp(13),
      ADR3 => VCC,
      O => tx_input_addr_inst_lut3_29
    );
  tx_input_addr_inst_lut3_301 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => VCC,
      ADR2 => tx_input_addr_30,
      ADR3 => txbp(14),
      O => tx_input_addr_inst_lut3_30
    );
  tx_input_addr_29_COUTUSED : X_BUF
    port map (
      I => tx_input_addr_29_CYMUXG,
      O => tx_input_addr_inst_cy_149
    );
  tx_input_addr_inst_cy_149_1457 : X_MUX2
    port map (
      IA => tx_input_addr_29_LOGIC_ZERO,
      IB => tx_input_addr_inst_cy_148,
      SEL => tx_input_addr_inst_lut3_30,
      O => tx_input_addr_29_CYMUXG
    );
  tx_input_addr_inst_sum_141_1458 : X_XOR2
    port map (
      I0 => tx_input_addr_inst_cy_148,
      I1 => tx_input_addr_inst_lut3_30,
      O => tx_input_addr_inst_sum_141
    );
  tx_input_addr_29_CYINIT_1459 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_147,
      O => tx_input_addr_29_CYINIT
    );
  tx_input_addr_inst_sum_142_1460 : X_XOR2
    port map (
      I0 => tx_input_addr_31_CYINIT,
      I1 => tx_input_addr_inst_lut3_31,
      O => tx_input_addr_inst_sum_142
    );
  tx_input_addr_inst_lut3_311 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => txbp(15),
      ADR1 => tx_input_addr_31,
      ADR2 => tx_input_cs_FFd12,
      ADR3 => VCC,
      O => tx_input_addr_inst_lut3_31
    );
  tx_input_addr_31_CYINIT_1461 : X_BUF
    port map (
      I => tx_input_addr_inst_cy_149,
      O => tx_input_addr_31_CYINIT
    );
  mac_control_rxf_cnt_0_LOGIC_ZERO_1462 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_0_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_16_1463 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_26,
      IB => mac_control_rxf_cnt_0_LOGIC_ZERO,
      SEL => mac_control_rxf_cnt_Madd_n0000_inst_lut2_16,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_16
    );
  mac_control_rxf_cnt_Madd_n0000_inst_lut2_161 : X_LUT4
    generic map(
      INIT => X"00FF"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_26,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(0),
      O => mac_control_rxf_cnt_Madd_n0000_inst_lut2_16
    );
  mac_control_rxf_cnt_0_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_41,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(1),
      O => mac_control_rxf_cnt_0_GROM
    );
  mac_control_rxf_cnt_0_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_0_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_17
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_17_1464 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_41,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_16,
      SEL => mac_control_rxf_cnt_0_GROM,
      O => mac_control_rxf_cnt_0_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_17 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_16,
      I1 => mac_control_rxf_cnt_0_GROM,
      O => mac_control_rxf_cnt_n0000(1)
    );
  mac_control_rxf_cnt_2_LOGIC_ZERO_1465 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_2_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_18_1466 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_2_CYINIT,
      SEL => mac_control_rxf_cnt_2_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_18
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_18 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_2_CYINIT,
      I1 => mac_control_rxf_cnt_2_FROM,
      O => mac_control_rxf_cnt_n0000(2)
    );
  mac_control_rxf_cnt_2_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(2),
      O => mac_control_rxf_cnt_2_FROM
    );
  mac_control_rxf_cnt_2_G : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxf_cnt(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxf_cnt_2_GROM
    );
  mac_control_rxf_cnt_2_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_2_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_19
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_19_1467 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_2_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_18,
      SEL => mac_control_rxf_cnt_2_GROM,
      O => mac_control_rxf_cnt_2_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_19 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_18,
      I1 => mac_control_rxf_cnt_2_GROM,
      O => mac_control_rxf_cnt_n0000(3)
    );
  mac_control_rxf_cnt_2_CYINIT_1468 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_17,
      O => mac_control_rxf_cnt_2_CYINIT
    );
  mac_control_rxf_cnt_4_LOGIC_ZERO_1469 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_4_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_20_1470 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_4_CYINIT,
      SEL => mac_control_rxf_cnt_4_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_20
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_20 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_4_CYINIT,
      I1 => mac_control_rxf_cnt_4_FROM,
      O => mac_control_rxf_cnt_n0000(4)
    );
  mac_control_rxf_cnt_4_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(4),
      O => mac_control_rxf_cnt_4_FROM
    );
  mac_control_rxf_cnt_4_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(5),
      O => mac_control_rxf_cnt_4_GROM
    );
  mac_control_rxf_cnt_4_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_4_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_21
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_21_1471 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_4_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_20,
      SEL => mac_control_rxf_cnt_4_GROM,
      O => mac_control_rxf_cnt_4_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_21 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_20,
      I1 => mac_control_rxf_cnt_4_GROM,
      O => mac_control_rxf_cnt_n0000(5)
    );
  mac_control_rxf_cnt_4_CYINIT_1472 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_19,
      O => mac_control_rxf_cnt_4_CYINIT
    );
  mac_control_rxf_cnt_6_LOGIC_ZERO_1473 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_6_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_22_1474 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_6_CYINIT,
      SEL => mac_control_rxf_cnt_6_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_22
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_22 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_6_CYINIT,
      I1 => mac_control_rxf_cnt_6_FROM,
      O => mac_control_rxf_cnt_n0000(6)
    );
  mac_control_rxf_cnt_6_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(6),
      O => mac_control_rxf_cnt_6_FROM
    );
  mac_control_rxf_cnt_6_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(7),
      O => mac_control_rxf_cnt_6_GROM
    );
  mac_control_rxf_cnt_6_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_6_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_23
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_23_1475 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_6_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_22,
      SEL => mac_control_rxf_cnt_6_GROM,
      O => mac_control_rxf_cnt_6_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_23 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_22,
      I1 => mac_control_rxf_cnt_6_GROM,
      O => mac_control_rxf_cnt_n0000(7)
    );
  mac_control_rxf_cnt_6_CYINIT_1476 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_21,
      O => mac_control_rxf_cnt_6_CYINIT
    );
  mac_control_rxf_cnt_8_LOGIC_ZERO_1477 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_8_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_24_1478 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_8_CYINIT,
      SEL => mac_control_rxf_cnt_8_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_24
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_24 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_8_CYINIT,
      I1 => mac_control_rxf_cnt_8_FROM,
      O => mac_control_rxf_cnt_n0000(8)
    );
  mac_control_rxf_cnt_8_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(8),
      O => mac_control_rxf_cnt_8_FROM
    );
  mac_control_rxf_cnt_8_G : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(9),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_8_GROM
    );
  mac_control_rxf_cnt_8_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_8_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_25
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_25_1479 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_8_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_24,
      SEL => mac_control_rxf_cnt_8_GROM,
      O => mac_control_rxf_cnt_8_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_25 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_24,
      I1 => mac_control_rxf_cnt_8_GROM,
      O => mac_control_rxf_cnt_n0000(9)
    );
  mac_control_rxf_cnt_8_CYINIT_1480 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_23,
      O => mac_control_rxf_cnt_8_CYINIT
    );
  mac_control_rxf_cnt_10_LOGIC_ZERO_1481 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_10_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_26_1482 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_10_CYINIT,
      SEL => mac_control_rxf_cnt_10_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_26
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_26 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_10_CYINIT,
      I1 => mac_control_rxf_cnt_10_FROM,
      O => mac_control_rxf_cnt_n0000(10)
    );
  mac_control_rxf_cnt_10_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(10),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_10_FROM
    );
  mac_control_rxf_cnt_10_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(11),
      O => mac_control_rxf_cnt_10_GROM
    );
  mac_control_rxf_cnt_10_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_10_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_27
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_27_1483 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_10_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_26,
      SEL => mac_control_rxf_cnt_10_GROM,
      O => mac_control_rxf_cnt_10_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_27 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_26,
      I1 => mac_control_rxf_cnt_10_GROM,
      O => mac_control_rxf_cnt_n0000(11)
    );
  mac_control_rxf_cnt_10_CYINIT_1484 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_25,
      O => mac_control_rxf_cnt_10_CYINIT
    );
  rx_output_cs_FFd9_1485 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd9_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd9_FFY_RST,
      O => rx_output_cs_FFd9
    );
  rx_output_cs_FFd9_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd9_FFY_RST
    );
  mac_control_rxf_cnt_12_LOGIC_ZERO_1486 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_12_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_28_1487 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_12_CYINIT,
      SEL => mac_control_rxf_cnt_12_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_28
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_28 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_12_CYINIT,
      I1 => mac_control_rxf_cnt_12_FROM,
      O => mac_control_rxf_cnt_n0000(12)
    );
  mac_control_rxf_cnt_12_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(12),
      O => mac_control_rxf_cnt_12_FROM
    );
  mac_control_rxf_cnt_12_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(13),
      O => mac_control_rxf_cnt_12_GROM
    );
  mac_control_rxf_cnt_12_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_12_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_29
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_29_1488 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_12_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_28,
      SEL => mac_control_rxf_cnt_12_GROM,
      O => mac_control_rxf_cnt_12_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_29 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_28,
      I1 => mac_control_rxf_cnt_12_GROM,
      O => mac_control_rxf_cnt_n0000(13)
    );
  mac_control_rxf_cnt_12_CYINIT_1489 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_27,
      O => mac_control_rxf_cnt_12_CYINIT
    );
  mac_control_rxf_cnt_14_LOGIC_ZERO_1490 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_14_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_30_1491 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_14_CYINIT,
      SEL => mac_control_rxf_cnt_14_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_30
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_30 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_14_CYINIT,
      I1 => mac_control_rxf_cnt_14_FROM,
      O => mac_control_rxf_cnt_n0000(14)
    );
  mac_control_rxf_cnt_14_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(14),
      O => mac_control_rxf_cnt_14_FROM
    );
  mac_control_rxf_cnt_14_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(15),
      O => mac_control_rxf_cnt_14_GROM
    );
  mac_control_rxf_cnt_14_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_14_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_31
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_31_1492 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_14_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_30,
      SEL => mac_control_rxf_cnt_14_GROM,
      O => mac_control_rxf_cnt_14_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_31 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_30,
      I1 => mac_control_rxf_cnt_14_GROM,
      O => mac_control_rxf_cnt_n0000(15)
    );
  mac_control_rxf_cnt_14_CYINIT_1493 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_29,
      O => mac_control_rxf_cnt_14_CYINIT
    );
  mac_control_rxf_cnt_16_LOGIC_ZERO_1494 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_16_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_32_1495 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_16_CYINIT,
      SEL => mac_control_rxf_cnt_16_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_32
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_32 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_16_CYINIT,
      I1 => mac_control_rxf_cnt_16_FROM,
      O => mac_control_rxf_cnt_n0000(16)
    );
  mac_control_rxf_cnt_16_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(16),
      O => mac_control_rxf_cnt_16_FROM
    );
  mac_control_rxf_cnt_16_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(17),
      O => mac_control_rxf_cnt_16_GROM
    );
  mac_control_rxf_cnt_16_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_16_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_33
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_33_1496 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_16_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_32,
      SEL => mac_control_rxf_cnt_16_GROM,
      O => mac_control_rxf_cnt_16_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_33 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_32,
      I1 => mac_control_rxf_cnt_16_GROM,
      O => mac_control_rxf_cnt_n0000(17)
    );
  mac_control_rxf_cnt_16_CYINIT_1497 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_31,
      O => mac_control_rxf_cnt_16_CYINIT
    );
  mac_control_rxf_cnt_18_LOGIC_ZERO_1498 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_18_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_34_1499 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_18_CYINIT,
      SEL => mac_control_rxf_cnt_18_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_34
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_34 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_18_CYINIT,
      I1 => mac_control_rxf_cnt_18_FROM,
      O => mac_control_rxf_cnt_n0000(18)
    );
  mac_control_rxf_cnt_18_F : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_rxf_cnt(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_rxf_cnt_18_FROM
    );
  mac_control_rxf_cnt_18_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(19),
      O => mac_control_rxf_cnt_18_GROM
    );
  mac_control_rxf_cnt_18_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_18_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_35
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_35_1500 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_18_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_34,
      SEL => mac_control_rxf_cnt_18_GROM,
      O => mac_control_rxf_cnt_18_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_35 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_34,
      I1 => mac_control_rxf_cnt_18_GROM,
      O => mac_control_rxf_cnt_n0000(19)
    );
  mac_control_rxf_cnt_18_CYINIT_1501 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_33,
      O => mac_control_rxf_cnt_18_CYINIT
    );
  mac_control_rxf_cnt_20_LOGIC_ZERO_1502 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_20_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_36_1503 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_20_CYINIT,
      SEL => mac_control_rxf_cnt_20_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_36
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_36 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_20_CYINIT,
      I1 => mac_control_rxf_cnt_20_FROM,
      O => mac_control_rxf_cnt_n0000(20)
    );
  mac_control_rxf_cnt_20_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(20),
      O => mac_control_rxf_cnt_20_FROM
    );
  mac_control_rxf_cnt_20_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(21),
      O => mac_control_rxf_cnt_20_GROM
    );
  mac_control_rxf_cnt_20_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_20_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_37
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_37_1504 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_20_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_36,
      SEL => mac_control_rxf_cnt_20_GROM,
      O => mac_control_rxf_cnt_20_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_37 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_36,
      I1 => mac_control_rxf_cnt_20_GROM,
      O => mac_control_rxf_cnt_n0000(21)
    );
  mac_control_rxf_cnt_20_CYINIT_1505 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_35,
      O => mac_control_rxf_cnt_20_CYINIT
    );
  mac_control_rxf_cnt_22_LOGIC_ZERO_1506 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_22_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_38_1507 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_22_CYINIT,
      SEL => mac_control_rxf_cnt_22_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_38
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_38 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_22_CYINIT,
      I1 => mac_control_rxf_cnt_22_FROM,
      O => mac_control_rxf_cnt_n0000(22)
    );
  mac_control_rxf_cnt_22_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(22),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_22_FROM
    );
  mac_control_rxf_cnt_22_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(23),
      O => mac_control_rxf_cnt_22_GROM
    );
  mac_control_rxf_cnt_22_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_22_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_39
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_39_1508 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_22_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_38,
      SEL => mac_control_rxf_cnt_22_GROM,
      O => mac_control_rxf_cnt_22_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_39 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_38,
      I1 => mac_control_rxf_cnt_22_GROM,
      O => mac_control_rxf_cnt_n0000(23)
    );
  mac_control_rxf_cnt_22_CYINIT_1509 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_37,
      O => mac_control_rxf_cnt_22_CYINIT
    );
  mac_control_rxf_cnt_24_LOGIC_ZERO_1510 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_24_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_40_1511 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_24_CYINIT,
      SEL => mac_control_rxf_cnt_24_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_40
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_40 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_24_CYINIT,
      I1 => mac_control_rxf_cnt_24_FROM,
      O => mac_control_rxf_cnt_n0000(24)
    );
  mac_control_rxf_cnt_24_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(24),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_24_FROM
    );
  mac_control_rxf_cnt_24_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(25),
      O => mac_control_rxf_cnt_24_GROM
    );
  mac_control_rxf_cnt_24_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_24_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_41
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_41_1512 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_24_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_40,
      SEL => mac_control_rxf_cnt_24_GROM,
      O => mac_control_rxf_cnt_24_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_41 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_40,
      I1 => mac_control_rxf_cnt_24_GROM,
      O => mac_control_rxf_cnt_n0000(25)
    );
  mac_control_rxf_cnt_24_CYINIT_1513 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_39,
      O => mac_control_rxf_cnt_24_CYINIT
    );
  mac_control_rxf_cnt_26_LOGIC_ZERO_1514 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_26_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_42_1515 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_26_CYINIT,
      SEL => mac_control_rxf_cnt_26_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_42
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_42 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_26_CYINIT,
      I1 => mac_control_rxf_cnt_26_FROM,
      O => mac_control_rxf_cnt_n0000(26)
    );
  mac_control_rxf_cnt_26_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(26),
      O => mac_control_rxf_cnt_26_FROM
    );
  mac_control_rxf_cnt_26_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(27),
      O => mac_control_rxf_cnt_26_GROM
    );
  mac_control_rxf_cnt_26_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_26_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_43
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_43_1516 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_26_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_42,
      SEL => mac_control_rxf_cnt_26_GROM,
      O => mac_control_rxf_cnt_26_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_43 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_42,
      I1 => mac_control_rxf_cnt_26_GROM,
      O => mac_control_rxf_cnt_n0000(27)
    );
  mac_control_rxf_cnt_26_CYINIT_1517 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_41,
      O => mac_control_rxf_cnt_26_CYINIT
    );
  mac_control_rxf_cnt_28_LOGIC_ZERO_1518 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_28_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_44_1519 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_28_CYINIT,
      SEL => mac_control_rxf_cnt_28_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_44
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_44 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_28_CYINIT,
      I1 => mac_control_rxf_cnt_28_FROM,
      O => mac_control_rxf_cnt_n0000(28)
    );
  mac_control_rxf_cnt_28_F : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(28),
      O => mac_control_rxf_cnt_28_FROM
    );
  mac_control_rxf_cnt_28_G : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(29),
      O => mac_control_rxf_cnt_28_GROM
    );
  mac_control_rxf_cnt_28_COUTUSED : X_BUF
    port map (
      I => mac_control_rxf_cnt_28_CYMUXG,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_45
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_45_1520 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_28_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_Madd_n0000_inst_cy_44,
      SEL => mac_control_rxf_cnt_28_GROM,
      O => mac_control_rxf_cnt_28_CYMUXG
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_45 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_44,
      I1 => mac_control_rxf_cnt_28_GROM,
      O => mac_control_rxf_cnt_n0000(29)
    );
  mac_control_rxf_cnt_28_CYINIT_1521 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_43,
      O => mac_control_rxf_cnt_28_CYINIT
    );
  mac_control_rxf_cnt_30_LOGIC_ZERO_1522 : X_ZERO
    port map (
      O => mac_control_rxf_cnt_30_LOGIC_ZERO
    );
  mac_control_rxf_cnt_Madd_n0000_inst_cy_46_1523 : X_MUX2
    port map (
      IA => mac_control_rxf_cnt_30_LOGIC_ZERO,
      IB => mac_control_rxf_cnt_30_CYINIT,
      SEL => mac_control_rxf_cnt_30_FROM,
      O => mac_control_rxf_cnt_Madd_n0000_inst_cy_46
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_46 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_30_CYINIT,
      I1 => mac_control_rxf_cnt_30_FROM,
      O => mac_control_rxf_cnt_n0000(30)
    );
  mac_control_rxf_cnt_30_F : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_rxf_cnt(30),
      ADR3 => VCC,
      O => mac_control_rxf_cnt_30_FROM
    );
  mac_control_rxf_cnt_31_rt_1524 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_rxf_cnt(31),
      O => mac_control_rxf_cnt_31_rt
    );
  mac_control_rxf_cnt_Madd_n0000_inst_sum_47 : X_XOR2
    port map (
      I0 => mac_control_rxf_cnt_Madd_n0000_inst_cy_46,
      I1 => mac_control_rxf_cnt_31_rt,
      O => mac_control_rxf_cnt_n0000(31)
    );
  mac_control_rxf_cnt_30_CYINIT_1525 : X_BUF
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_cy_45,
      O => mac_control_rxf_cnt_30_CYINIT
    );
  mac_control_PHY_status_MII_Interface_dreg_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(2),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_4_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(3)
    );
  mac_control_PHY_status_MII_Interface_dreg_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_4_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(1),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_2_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(2)
    );
  mac_control_PHY_status_MII_Interface_dreg_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_2_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(3),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_4_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(4)
    );
  mac_control_PHY_status_MII_Interface_dreg_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_4_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(5),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_6_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(6)
    );
  mac_control_PHY_status_MII_Interface_dreg_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_6_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(6),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_8_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(7)
    );
  mac_control_PHY_status_MII_Interface_dreg_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_8_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(7),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_8_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(8)
    );
  mac_control_PHY_status_MII_Interface_dreg_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_8_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(9),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_10_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(10)
    );
  mac_control_PHY_status_MII_Interface_dreg_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_10_FFX_RST
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ONE_1526 : X_ONE
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ONE
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ZERO_1527 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_177_1528 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ONE,
      SEL => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_12,
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_177
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_121 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(1),
      ADR1 => rx_input_memio_addrchk_datal(0),
      ADR2 => rx_input_memio_addrchk_datal(1),
      ADR3 => rx_input_memio_addrchk_macaddrl(0),
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_12
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_131 : X_LUT4
    generic map(
      INIT => X"9009"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_datal(2),
      ADR1 => rx_input_memio_addrchk_macaddrl(2),
      ADR2 => rx_input_memio_addrchk_datal(3),
      ADR3 => rx_input_memio_addrchk_macaddrl(3),
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_13
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_CYMUXG,
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_1529 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_177,
      SEL => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_13,
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_5_LOGIC_ZERO_1530 : X_ZERO
    port map (
      O => rx_input_memio_addrchk_lmaceq_5_LOGIC_ZERO
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_179_1531 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_5_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_lmaceq_5_CYINIT,
      SEL => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_14,
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_179
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_141 : X_LUT4
    generic map(
      INIT => X"8421"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(5),
      ADR1 => rx_input_memio_addrchk_datal(4),
      ADR2 => rx_input_memio_addrchk_datal(5),
      ADR3 => rx_input_memio_addrchk_macaddrl(4),
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_14
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_151 : X_LUT4
    generic map(
      INIT => X"8241"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_macaddrl(7),
      ADR1 => rx_input_memio_addrchk_datal(6),
      ADR2 => rx_input_memio_addrchk_macaddrl(6),
      ADR3 => rx_input_memio_addrchk_datal(7),
      O => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_15
    );
  rx_input_memio_addrchk_lmaceq_5_COUTUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq_5_CYMUXG,
      O => rx_input_memio_addrchk_lmaceq(5)
    );
  rx_input_memio_addrchk_Mcompar_n0033_inst_cy_180 : X_MUX2
    port map (
      IA => rx_input_memio_addrchk_lmaceq_5_LOGIC_ZERO,
      IB => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_179,
      SEL => rx_input_memio_addrchk_Mcompar_n0033_inst_lut4_15,
      O => rx_input_memio_addrchk_lmaceq_5_CYMUXG
    );
  rx_input_memio_addrchk_lmaceq_5_CYINIT_1532 : X_BUF
    port map (
      I => rx_input_memio_addrchk_Mcompar_n0033_inst_cy_178,
      O => rx_input_memio_addrchk_lmaceq_5_CYINIT
    );
  rx_output_fifo_N9_LOGIC_ZERO_1533 : X_ZERO
    port map (
      O => rx_output_fifo_N9_LOGIC_ZERO
    );
  rx_output_fifo_BU199 : X_MUX2
    port map (
      IA => rx_output_fifo_N9,
      IB => rx_output_fifo_N9_CYINIT,
      SEL => rx_output_fifo_N2840,
      O => rx_output_fifo_N2842
    );
  rx_output_fifo_BU200 : X_XOR2
    port map (
      I0 => rx_output_fifo_N9_CYINIT,
      I1 => rx_output_fifo_N2840,
      O => rx_output_fifo_N2832
    );
  rx_output_fifo_BU198 : X_LUT4
    generic map(
      INIT => X"5555"
    )
    port map (
      ADR0 => rx_output_fifo_N9,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N2840
    );
  rx_output_fifo_N9_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N8,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N9_GROM
    );
  rx_output_fifo_N9_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N9_CYMUXG,
      O => rx_output_fifo_N2847
    );
  rx_output_fifo_BU205 : X_MUX2
    port map (
      IA => rx_output_fifo_N8,
      IB => rx_output_fifo_N2842,
      SEL => rx_output_fifo_N9_GROM,
      O => rx_output_fifo_N9_CYMUXG
    );
  rx_output_fifo_BU206 : X_XOR2
    port map (
      I0 => rx_output_fifo_N2842,
      I1 => rx_output_fifo_N9_GROM,
      O => rx_output_fifo_N2833
    );
  rx_output_fifo_N9_CYINIT_1534 : X_BUF
    port map (
      I => rx_output_fifo_N9_LOGIC_ZERO,
      O => rx_output_fifo_N9_CYINIT
    );
  rx_output_fifo_BU211 : X_MUX2
    port map (
      IA => rx_output_fifo_N7,
      IB => rx_output_fifo_N7_CYINIT,
      SEL => rx_output_fifo_N7_FROM,
      O => rx_output_fifo_N2852
    );
  rx_output_fifo_BU212 : X_XOR2
    port map (
      I0 => rx_output_fifo_N7_CYINIT,
      I1 => rx_output_fifo_N7_FROM,
      O => rx_output_fifo_N2834
    );
  rx_output_fifo_N7_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N7,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N7_FROM
    );
  rx_output_fifo_N7_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N6,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N7_GROM
    );
  rx_output_fifo_N7_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N7_CYMUXG,
      O => rx_output_fifo_N2857
    );
  rx_output_fifo_BU217 : X_MUX2
    port map (
      IA => rx_output_fifo_N6,
      IB => rx_output_fifo_N2852,
      SEL => rx_output_fifo_N7_GROM,
      O => rx_output_fifo_N7_CYMUXG
    );
  rx_output_fifo_BU218 : X_XOR2
    port map (
      I0 => rx_output_fifo_N2852,
      I1 => rx_output_fifo_N7_GROM,
      O => rx_output_fifo_N2835
    );
  rx_output_fifo_N7_CYINIT_1535 : X_BUF
    port map (
      I => rx_output_fifo_N2847,
      O => rx_output_fifo_N7_CYINIT
    );
  rx_output_fifo_BU223 : X_MUX2
    port map (
      IA => rx_output_fifo_N5,
      IB => rx_output_fifo_N5_CYINIT,
      SEL => rx_output_fifo_N5_FROM,
      O => rx_output_fifo_N2862
    );
  rx_output_fifo_BU224 : X_XOR2
    port map (
      I0 => rx_output_fifo_N5_CYINIT,
      I1 => rx_output_fifo_N5_FROM,
      O => rx_output_fifo_N2836
    );
  rx_output_fifo_N5_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N5,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N5_FROM
    );
  rx_output_fifo_N5_G : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N4,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N5_GROM
    );
  rx_output_fifo_N5_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N5_CYMUXG,
      O => rx_output_fifo_N2867
    );
  rx_output_fifo_BU229 : X_MUX2
    port map (
      IA => rx_output_fifo_N4,
      IB => rx_output_fifo_N2862,
      SEL => rx_output_fifo_N5_GROM,
      O => rx_output_fifo_N5_CYMUXG
    );
  rx_output_fifo_BU230 : X_XOR2
    port map (
      I0 => rx_output_fifo_N2862,
      I1 => rx_output_fifo_N5_GROM,
      O => rx_output_fifo_N2837
    );
  rx_output_fifo_N5_CYINIT_1536 : X_BUF
    port map (
      I => rx_output_fifo_N2857,
      O => rx_output_fifo_N5_CYINIT
    );
  rx_output_fifo_BU235 : X_MUX2
    port map (
      IA => rx_output_fifo_N3,
      IB => rx_output_fifo_N3_CYINIT,
      SEL => rx_output_fifo_N3_FROM,
      O => rx_output_fifo_N2872
    );
  rx_output_fifo_BU236 : X_XOR2
    port map (
      I0 => rx_output_fifo_N3_CYINIT,
      I1 => rx_output_fifo_N3_FROM,
      O => rx_output_fifo_N2838
    );
  rx_output_fifo_N3_F : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N3_FROM
    );
  rx_output_fifo_N2_rt_1537 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => rx_output_fifo_N2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N2_rt
    );
  rx_output_fifo_BU241 : X_XOR2
    port map (
      I0 => rx_output_fifo_N2872,
      I1 => rx_output_fifo_N2_rt,
      O => rx_output_fifo_N2839
    );
  rx_output_fifo_N3_CYINIT_1538 : X_BUF
    port map (
      I => rx_output_fifo_N2867,
      O => rx_output_fifo_N3_CYINIT
    );
  rx_output_fifo_N2576_LOGIC_ONE_1539 : X_ONE
    port map (
      O => rx_output_fifo_N2576_LOGIC_ONE
    );
  rx_output_fifo_N2576_LOGIC_ZERO_1540 : X_ZERO
    port map (
      O => rx_output_fifo_N2576_LOGIC_ZERO
    );
  rx_output_fifo_BU151 : X_MUX2
    port map (
      IA => rx_output_fifo_N2576_LOGIC_ZERO,
      IB => rx_output_fifo_N2576_LOGIC_ONE,
      SEL => rx_output_fifo_N2569,
      O => rx_output_fifo_N2577
    );
  rx_output_fifo_BU150 : X_LUT4
    generic map(
      INIT => X"99C3"
    )
    port map (
      ADR0 => rx_output_fifo_N1617,
      ADR1 => rx_output_fifo_N1553,
      ADR2 => rx_output_fifo_N1633,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N2569
    );
  rx_output_fifo_BU153 : X_LUT4
    generic map(
      INIT => X"9A95"
    )
    port map (
      ADR0 => rx_output_fifo_N1552,
      ADR1 => rx_output_fifo_N1616,
      ADR2 => rx_output_fifo_empty,
      ADR3 => rx_output_fifo_N1632,
      O => rx_output_fifo_N2568
    );
  rx_output_fifo_N2576_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N2576_CYMUXG,
      O => rx_output_fifo_N2576
    );
  rx_output_fifo_BU154 : X_MUX2
    port map (
      IA => rx_output_fifo_N2576_LOGIC_ZERO,
      IB => rx_output_fifo_N2577,
      SEL => rx_output_fifo_N2568,
      O => rx_output_fifo_N2576_CYMUXG
    );
  rx_output_fifo_N2574_LOGIC_ZERO_1541 : X_ZERO
    port map (
      O => rx_output_fifo_N2574_LOGIC_ZERO
    );
  rx_output_fifo_BU157 : X_MUX2
    port map (
      IA => rx_output_fifo_N2574_LOGIC_ZERO,
      IB => rx_output_fifo_N2574_CYINIT,
      SEL => rx_output_fifo_N2567,
      O => rx_output_fifo_N2575
    );
  rx_output_fifo_BU156 : X_LUT4
    generic map(
      INIT => X"C939"
    )
    port map (
      ADR0 => rx_output_fifo_N1631,
      ADR1 => rx_output_fifo_N1551,
      ADR2 => rx_output_fifo_empty,
      ADR3 => rx_output_fifo_N1615,
      O => rx_output_fifo_N2567
    );
  rx_output_fifo_BU159 : X_LUT4
    generic map(
      INIT => X"A959"
    )
    port map (
      ADR0 => rx_output_fifo_N1550,
      ADR1 => rx_output_fifo_N1630,
      ADR2 => rx_output_fifo_empty,
      ADR3 => rx_output_fifo_N1614,
      O => rx_output_fifo_N2566
    );
  rx_output_fifo_N2574_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N2574_CYMUXG,
      O => rx_output_fifo_N2574
    );
  rx_output_fifo_BU160 : X_MUX2
    port map (
      IA => rx_output_fifo_N2574_LOGIC_ZERO,
      IB => rx_output_fifo_N2575,
      SEL => rx_output_fifo_N2566,
      O => rx_output_fifo_N2574_CYMUXG
    );
  rx_output_fifo_N2574_CYINIT_1542 : X_BUF
    port map (
      I => rx_output_fifo_N2576,
      O => rx_output_fifo_N2574_CYINIT
    );
  rx_output_fifo_N2572_LOGIC_ZERO_1543 : X_ZERO
    port map (
      O => rx_output_fifo_N2572_LOGIC_ZERO
    );
  rx_output_fifo_BU163 : X_MUX2
    port map (
      IA => rx_output_fifo_N2572_LOGIC_ZERO,
      IB => rx_output_fifo_N2572_CYINIT,
      SEL => rx_output_fifo_N2565,
      O => rx_output_fifo_N2573
    );
  rx_output_fifo_BU162 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => rx_output_fifo_N1629,
      ADR1 => rx_output_fifo_N1549,
      ADR2 => rx_output_fifo_N1613,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N2565
    );
  rx_output_fifo_BU165 : X_LUT4
    generic map(
      INIT => X"99A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1548,
      ADR1 => rx_output_fifo_N1612,
      ADR2 => rx_output_fifo_N1628,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N2564
    );
  rx_output_fifo_N2572_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N2572_CYMUXG,
      O => rx_output_fifo_N2572
    );
  rx_output_fifo_BU166 : X_MUX2
    port map (
      IA => rx_output_fifo_N2572_LOGIC_ZERO,
      IB => rx_output_fifo_N2573,
      SEL => rx_output_fifo_N2564,
      O => rx_output_fifo_N2572_CYMUXG
    );
  rx_output_fifo_N2572_CYINIT_1544 : X_BUF
    port map (
      I => rx_output_fifo_N2574,
      O => rx_output_fifo_N2572_CYINIT
    );
  tx_output_crcl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_6_1_O,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_6_FFY_RST,
      O => tx_output_crcl(6)
    );
  tx_output_crcl_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_6_FFY_RST
    );
  rx_output_fifo_BU172_O_LOGIC_ZERO_1545 : X_ZERO
    port map (
      O => rx_output_fifo_BU172_O_LOGIC_ZERO
    );
  rx_output_fifo_BU169 : X_MUX2
    port map (
      IA => rx_output_fifo_BU172_O_LOGIC_ZERO,
      IB => rx_output_fifo_BU172_O_CYINIT,
      SEL => rx_output_fifo_N2563,
      O => rx_output_fifo_N2571
    );
  rx_output_fifo_BU168 : X_LUT4
    generic map(
      INIT => X"99C3"
    )
    port map (
      ADR0 => rx_output_fifo_N1611,
      ADR1 => rx_output_fifo_N1547,
      ADR2 => rx_output_fifo_N1627,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N2563
    );
  rx_output_fifo_BU171 : X_LUT4
    generic map(
      INIT => X"99C3"
    )
    port map (
      ADR0 => rx_output_fifo_N1610,
      ADR1 => rx_output_fifo_N1546,
      ADR2 => rx_output_fifo_N1626,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_fifo_N2562
    );
  rx_output_fifo_BU172_O_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_BU172_O_CYMUXG,
      O => rx_output_fifo_BU172_O
    );
  rx_output_fifo_BU172 : X_MUX2
    port map (
      IA => rx_output_fifo_BU172_O_LOGIC_ZERO,
      IB => rx_output_fifo_N2571,
      SEL => rx_output_fifo_N2562,
      O => rx_output_fifo_BU172_O_CYMUXG
    );
  rx_output_fifo_BU172_O_CYINIT_1546 : X_BUF
    port map (
      I => rx_output_fifo_N2572,
      O => rx_output_fifo_BU172_O_CYINIT
    );
  rx_output_fifo_BU175 : X_XOR2
    port map (
      I0 => rx_output_fifo_empty_CYINIT,
      I1 => rx_output_fifo_empty_FROM,
      O => rx_output_fifo_N2580
    );
  rx_output_fifo_empty_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_empty_FROM
    );
  rx_output_fifo_empty_CYINIT_1547 : X_BUF
    port map (
      I => rx_output_fifo_BU172_O,
      O => rx_output_fifo_empty_CYINIT
    );
  rx_output_fifo_N3614_LOGIC_ONE_1548 : X_ONE
    port map (
      O => rx_output_fifo_N3614_LOGIC_ONE
    );
  rx_output_fifo_N3614_LOGIC_ZERO_1549 : X_ZERO
    port map (
      O => rx_output_fifo_N3614_LOGIC_ZERO
    );
  rx_output_fifo_BU330 : X_MUX2
    port map (
      IA => rx_output_fifo_N3614_LOGIC_ZERO,
      IB => rx_output_fifo_N3614_LOGIC_ONE,
      SEL => rx_output_fifo_N3607,
      O => rx_output_fifo_N3615
    );
  rx_output_fifo_BU329 : X_LUT4
    generic map(
      INIT => X"CA35"
    )
    port map (
      ADR0 => rx_output_fifo_N1577,
      ADR1 => rx_output_fifo_N1569,
      ADR2 => rx_output_fifo_full_0,
      ADR3 => rx_output_fifo_N1617,
      O => rx_output_fifo_N3607
    );
  rx_output_fifo_BU332 : X_LUT4
    generic map(
      INIT => X"9C93"
    )
    port map (
      ADR0 => rx_output_fifo_N1568,
      ADR1 => rx_output_fifo_N1616,
      ADR2 => rx_output_fifo_full_0,
      ADR3 => rx_output_fifo_N1576,
      O => rx_output_fifo_N3606
    );
  rx_output_fifo_N3614_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N3614_CYMUXG,
      O => rx_output_fifo_N3614
    );
  rx_output_fifo_BU333 : X_MUX2
    port map (
      IA => rx_output_fifo_N3614_LOGIC_ZERO,
      IB => rx_output_fifo_N3615,
      SEL => rx_output_fifo_N3606,
      O => rx_output_fifo_N3614_CYMUXG
    );
  rx_output_fifo_N3612_LOGIC_ZERO_1550 : X_ZERO
    port map (
      O => rx_output_fifo_N3612_LOGIC_ZERO
    );
  rx_output_fifo_BU336 : X_MUX2
    port map (
      IA => rx_output_fifo_N3612_LOGIC_ZERO,
      IB => rx_output_fifo_N3612_CYINIT,
      SEL => rx_output_fifo_N3605,
      O => rx_output_fifo_N3613
    );
  rx_output_fifo_BU335 : X_LUT4
    generic map(
      INIT => X"D287"
    )
    port map (
      ADR0 => rx_output_fifo_full_0,
      ADR1 => rx_output_fifo_N1567,
      ADR2 => rx_output_fifo_N1615,
      ADR3 => rx_output_fifo_N1575,
      O => rx_output_fifo_N3605
    );
  rx_output_fifo_BU338 : X_LUT4
    generic map(
      INIT => X"C3A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1574,
      ADR1 => rx_output_fifo_N1566,
      ADR2 => rx_output_fifo_N1614,
      ADR3 => rx_output_fifo_full_0,
      O => rx_output_fifo_N3604
    );
  rx_output_fifo_N3612_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N3612_CYMUXG,
      O => rx_output_fifo_N3612
    );
  rx_output_fifo_BU339 : X_MUX2
    port map (
      IA => rx_output_fifo_N3612_LOGIC_ZERO,
      IB => rx_output_fifo_N3613,
      SEL => rx_output_fifo_N3604,
      O => rx_output_fifo_N3612_CYMUXG
    );
  rx_output_fifo_N3612_CYINIT_1551 : X_BUF
    port map (
      I => rx_output_fifo_N3614,
      O => rx_output_fifo_N3612_CYINIT
    );
  rx_output_fifo_N3610_LOGIC_ZERO_1552 : X_ZERO
    port map (
      O => rx_output_fifo_N3610_LOGIC_ZERO
    );
  rx_output_fifo_BU342 : X_MUX2
    port map (
      IA => rx_output_fifo_N3610_LOGIC_ZERO,
      IB => rx_output_fifo_N3610_CYINIT,
      SEL => rx_output_fifo_N3603,
      O => rx_output_fifo_N3611
    );
  rx_output_fifo_BU341 : X_LUT4
    generic map(
      INIT => X"D287"
    )
    port map (
      ADR0 => rx_output_fifo_full_0,
      ADR1 => rx_output_fifo_N1565,
      ADR2 => rx_output_fifo_N1613,
      ADR3 => rx_output_fifo_N1573,
      O => rx_output_fifo_N3603
    );
  rx_output_fifo_BU344 : X_LUT4
    generic map(
      INIT => X"A695"
    )
    port map (
      ADR0 => rx_output_fifo_N1612,
      ADR1 => rx_output_fifo_full_0,
      ADR2 => rx_output_fifo_N1564,
      ADR3 => rx_output_fifo_N1572,
      O => rx_output_fifo_N3602
    );
  rx_output_fifo_N3610_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N3610_CYMUXG,
      O => rx_output_fifo_N3610
    );
  rx_output_fifo_BU345 : X_MUX2
    port map (
      IA => rx_output_fifo_N3610_LOGIC_ZERO,
      IB => rx_output_fifo_N3611,
      SEL => rx_output_fifo_N3602,
      O => rx_output_fifo_N3610_CYMUXG
    );
  rx_output_fifo_N3610_CYINIT_1553 : X_BUF
    port map (
      I => rx_output_fifo_N3612,
      O => rx_output_fifo_N3610_CYINIT
    );
  rx_output_fifo_BU351_O_LOGIC_ZERO_1554 : X_ZERO
    port map (
      O => rx_output_fifo_BU351_O_LOGIC_ZERO
    );
  rx_output_fifo_BU348 : X_MUX2
    port map (
      IA => rx_output_fifo_BU351_O_LOGIC_ZERO,
      IB => rx_output_fifo_BU351_O_CYINIT,
      SEL => rx_output_fifo_N3601,
      O => rx_output_fifo_N3609
    );
  rx_output_fifo_BU347 : X_LUT4
    generic map(
      INIT => X"CA35"
    )
    port map (
      ADR0 => rx_output_fifo_N1571,
      ADR1 => rx_output_fifo_N1563,
      ADR2 => rx_output_fifo_full_0,
      ADR3 => rx_output_fifo_N1611,
      O => rx_output_fifo_N3601
    );
  rx_output_fifo_BU350 : X_LUT4
    generic map(
      INIT => X"C693"
    )
    port map (
      ADR0 => rx_output_fifo_full_0,
      ADR1 => rx_output_fifo_N1610,
      ADR2 => rx_output_fifo_N1562,
      ADR3 => rx_output_fifo_N1570,
      O => rx_output_fifo_N3600
    );
  rx_output_fifo_BU351_O_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_BU351_O_CYMUXG,
      O => rx_output_fifo_BU351_O
    );
  rx_output_fifo_BU351 : X_MUX2
    port map (
      IA => rx_output_fifo_BU351_O_LOGIC_ZERO,
      IB => rx_output_fifo_N3609,
      SEL => rx_output_fifo_N3600,
      O => rx_output_fifo_BU351_O_CYMUXG
    );
  rx_output_fifo_BU351_O_CYINIT_1555 : X_BUF
    port map (
      I => rx_output_fifo_N3610,
      O => rx_output_fifo_BU351_O_CYINIT
    );
  rx_output_fifo_BU354 : X_XOR2
    port map (
      I0 => rx_output_fifo_full_CYINIT,
      I1 => rx_output_fifo_full_FROM,
      O => rx_output_fifo_N3618
    );
  rx_output_fifo_full_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_full_FROM
    );
  rx_output_fifo_full_CYINIT_1556 : X_BUF
    port map (
      I => rx_output_fifo_BU351_O,
      O => rx_output_fifo_full_CYINIT
    );
  rx_output_fifo_N4763_LOGIC_ONE_1557 : X_ONE
    port map (
      O => rx_output_fifo_N4763_LOGIC_ONE
    );
  rx_output_fifo_BU477 : X_MUX2
    port map (
      IA => rx_output_fifo_N1609,
      IB => rx_output_fifo_N4763_LOGIC_ONE,
      SEL => rx_output_fifo_N4756,
      O => rx_output_fifo_N4759
    );
  rx_output_fifo_BU476 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1609,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N1593,
      ADR3 => VCC,
      O => rx_output_fifo_N4756
    );
  rx_output_fifo_BU479 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => rx_output_fifo_N1608,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N1592,
      O => rx_output_fifo_N4760
    );
  rx_output_fifo_N4763_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N4763_CYMUXG,
      O => rx_output_fifo_N4763
    );
  rx_output_fifo_BU480 : X_MUX2
    port map (
      IA => rx_output_fifo_N1608,
      IB => rx_output_fifo_N4759,
      SEL => rx_output_fifo_N4760,
      O => rx_output_fifo_N4763_CYMUXG
    );
  rx_output_fifo_BU483 : X_MUX2
    port map (
      IA => rx_output_fifo_N1607,
      IB => rx_output_fifo_N4771_CYINIT,
      SEL => rx_output_fifo_N4764,
      O => rx_output_fifo_N4767
    );
  rx_output_fifo_BU482 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_output_fifo_N1607,
      ADR1 => rx_output_fifo_N1591,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N4764
    );
  rx_output_fifo_BU485 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1606,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N1590,
      ADR3 => VCC,
      O => rx_output_fifo_N4768
    );
  rx_output_fifo_N4771_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N4771_CYMUXG,
      O => rx_output_fifo_N4771
    );
  rx_output_fifo_BU486 : X_MUX2
    port map (
      IA => rx_output_fifo_N1606,
      IB => rx_output_fifo_N4767,
      SEL => rx_output_fifo_N4768,
      O => rx_output_fifo_N4771_CYMUXG
    );
  rx_output_fifo_N4771_CYINIT_1558 : X_BUF
    port map (
      I => rx_output_fifo_N4763,
      O => rx_output_fifo_N4771_CYINIT
    );
  rx_output_fifo_BU489 : X_MUX2
    port map (
      IA => rx_output_fifo_N1605,
      IB => rx_output_fifo_N4779_CYINIT,
      SEL => rx_output_fifo_N4772,
      O => rx_output_fifo_N4775
    );
  rx_output_fifo_BU488 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1605,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N1589,
      ADR3 => VCC,
      O => rx_output_fifo_N4772
    );
  rx_output_fifo_BU491 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1604,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N1588,
      ADR3 => VCC,
      O => rx_output_fifo_N4776
    );
  rx_output_fifo_N4779_COUTUSED : X_BUF
    port map (
      I => rx_output_fifo_N4779_CYMUXG,
      O => rx_output_fifo_N4779
    );
  rx_output_fifo_BU492 : X_MUX2
    port map (
      IA => rx_output_fifo_N1604,
      IB => rx_output_fifo_N4775,
      SEL => rx_output_fifo_N4776,
      O => rx_output_fifo_N4779_CYMUXG
    );
  rx_output_fifo_N4779_CYINIT_1559 : X_BUF
    port map (
      I => rx_output_fifo_N4771,
      O => rx_output_fifo_N4779_CYINIT
    );
  rx_output_fifo_BU495 : X_MUX2
    port map (
      IA => rx_output_fifo_N1603,
      IB => rx_output_fifo_wrcount_0_CYINIT,
      SEL => rx_output_fifo_N4780,
      O => rx_output_fifo_N4783
    );
  rx_output_fifo_BU496 : X_XOR2
    port map (
      I0 => rx_output_fifo_wrcount_0_CYINIT,
      I1 => rx_output_fifo_N4780,
      O => rx_output_fifo_N4754
    );
  rx_output_fifo_BU494 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => rx_output_fifo_N1603,
      ADR1 => rx_output_fifo_N1587,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N4780
    );
  rx_output_fifo_BU500 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => rx_output_fifo_N1602,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N1586,
      ADR3 => VCC,
      O => rx_output_fifo_N4786
    );
  rx_output_fifo_BU502 : X_XOR2
    port map (
      I0 => rx_output_fifo_N4783,
      I1 => rx_output_fifo_N4786,
      O => rx_output_fifo_N4755
    );
  rx_output_fifo_wrcount_0_CYINIT_1560 : X_BUF
    port map (
      I => rx_output_fifo_N4779,
      O => rx_output_fifo_wrcount_0_CYINIT
    );
  mac_control_bitcnt_104_LOGIC_ZERO_1561 : X_ZERO
    port map (
      O => mac_control_bitcnt_104_LOGIC_ZERO
    );
  mac_control_bitcnt_inst_cy_287_1562 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC1_30,
      IB => mac_control_bitcnt_104_LOGIC_ZERO,
      SEL => mac_control_Mshreg_scslll_103_rt,
      O => mac_control_bitcnt_inst_cy_287
    );
  mac_control_Mshreg_scslll_103_rt_1563 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => GLOBAL_LOGIC1_30,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_Mshreg_scslll_103,
      O => mac_control_Mshreg_scslll_103_rt
    );
  mac_control_bitcnt_inst_lut3_1861 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => GLOBAL_LOGIC0_44,
      ADR1 => mac_control_Mshreg_scslll_103,
      ADR2 => mac_control_bitcnt_104,
      ADR3 => VCC,
      O => mac_control_bitcnt_inst_lut3_186
    );
  mac_control_bitcnt_104_COUTUSED : X_BUF
    port map (
      I => mac_control_bitcnt_104_CYMUXG,
      O => mac_control_bitcnt_inst_cy_288
    );
  mac_control_bitcnt_inst_cy_288_1564 : X_MUX2
    port map (
      IA => GLOBAL_LOGIC0_44,
      IB => mac_control_bitcnt_inst_cy_287,
      SEL => mac_control_bitcnt_inst_lut3_186,
      O => mac_control_bitcnt_104_CYMUXG
    );
  mac_control_bitcnt_inst_sum_251_1565 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_inst_cy_287,
      I1 => mac_control_bitcnt_inst_lut3_186,
      O => mac_control_bitcnt_inst_sum_251
    );
  mac_control_bitcnt_105_LOGIC_ZERO_1566 : X_ZERO
    port map (
      O => mac_control_bitcnt_105_LOGIC_ZERO
    );
  mac_control_bitcnt_inst_cy_289_1567 : X_MUX2
    port map (
      IA => mac_control_bitcnt_105_LOGIC_ZERO,
      IB => mac_control_bitcnt_105_CYINIT,
      SEL => mac_control_bitcnt_inst_lut3_187,
      O => mac_control_bitcnt_inst_cy_289
    );
  mac_control_bitcnt_inst_sum_252_1568 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_105_CYINIT,
      I1 => mac_control_bitcnt_inst_lut3_187,
      O => mac_control_bitcnt_inst_sum_252
    );
  mac_control_bitcnt_inst_lut3_1871 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => mac_control_Mshreg_scslll_103,
      ADR1 => mac_control_bitcnt_105,
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_bitcnt_inst_lut3_187
    );
  mac_control_bitcnt_inst_lut3_1881 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => mac_control_bitcnt_106,
      ADR1 => VCC,
      ADR2 => mac_control_Mshreg_scslll_103,
      ADR3 => VCC,
      O => mac_control_bitcnt_inst_lut3_188
    );
  mac_control_bitcnt_105_COUTUSED : X_BUF
    port map (
      I => mac_control_bitcnt_105_CYMUXG,
      O => mac_control_bitcnt_inst_cy_290
    );
  mac_control_bitcnt_inst_cy_290_1569 : X_MUX2
    port map (
      IA => mac_control_bitcnt_105_LOGIC_ZERO,
      IB => mac_control_bitcnt_inst_cy_289,
      SEL => mac_control_bitcnt_inst_lut3_188,
      O => mac_control_bitcnt_105_CYMUXG
    );
  mac_control_bitcnt_inst_sum_253_1570 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_inst_cy_289,
      I1 => mac_control_bitcnt_inst_lut3_188,
      O => mac_control_bitcnt_inst_sum_253
    );
  mac_control_bitcnt_105_CYINIT_1571 : X_BUF
    port map (
      I => mac_control_bitcnt_inst_cy_288,
      O => mac_control_bitcnt_105_CYINIT
    );
  mac_control_bitcnt_107_LOGIC_ZERO_1572 : X_ZERO
    port map (
      O => mac_control_bitcnt_107_LOGIC_ZERO
    );
  mac_control_bitcnt_inst_cy_291_1573 : X_MUX2
    port map (
      IA => mac_control_bitcnt_107_LOGIC_ZERO,
      IB => mac_control_bitcnt_107_CYINIT,
      SEL => mac_control_bitcnt_inst_lut3_189,
      O => mac_control_bitcnt_inst_cy_291
    );
  mac_control_bitcnt_inst_sum_254_1574 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_107_CYINIT,
      I1 => mac_control_bitcnt_inst_lut3_189,
      O => mac_control_bitcnt_inst_sum_254
    );
  mac_control_bitcnt_inst_lut3_1891 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_bitcnt_107,
      ADR2 => VCC,
      ADR3 => mac_control_Mshreg_scslll_103,
      O => mac_control_bitcnt_inst_lut3_189
    );
  mac_control_bitcnt_inst_lut3_1901 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_bitcnt_108,
      ADR3 => mac_control_Mshreg_scslll_103,
      O => mac_control_bitcnt_inst_lut3_190
    );
  mac_control_bitcnt_107_COUTUSED : X_BUF
    port map (
      I => mac_control_bitcnt_107_CYMUXG,
      O => mac_control_bitcnt_inst_cy_292
    );
  mac_control_bitcnt_inst_cy_292_1575 : X_MUX2
    port map (
      IA => mac_control_bitcnt_107_LOGIC_ZERO,
      IB => mac_control_bitcnt_inst_cy_291,
      SEL => mac_control_bitcnt_inst_lut3_190,
      O => mac_control_bitcnt_107_CYMUXG
    );
  mac_control_bitcnt_inst_sum_255_1576 : X_XOR2
    port map (
      I0 => mac_control_bitcnt_inst_cy_291,
      I1 => mac_control_bitcnt_inst_lut3_190,
      O => mac_control_bitcnt_inst_sum_255
    );
  mac_control_bitcnt_107_CYINIT_1577 : X_BUF
    port map (
      I => mac_control_bitcnt_inst_cy_290,
      O => mac_control_bitcnt_107_CYINIT
    );
  tx_output_crc_loigc_Mxor_n0009_Result1 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_data(3),
      ADR3 => tx_output_crcl(28),
      O => tx_output_crc_loigc_n0115_0_FROM
    );
  tx_output_crc_loigc_Mxor_CO_15_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_Mxor_CO_13_Xo(2),
      ADR1 => tx_output_crcl(7),
      ADR2 => tx_output_crc_loigc_n0118(0),
      ADR3 => tx_output_crc_loigc_n0115(0),
      O => tx_output_crc_loigc_n0115_0_GROM
    );
  tx_output_crc_loigc_n0115_0_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0115_0_FROM,
      O => tx_output_crc_loigc_n0115(0)
    );
  tx_output_crc_loigc_n0115_0_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_n0115_0_GROM,
      O => tx_output_crc_15_Q
    );
  rx_input_memio_n0048_15_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_15_Q,
      O => rx_input_memio_n0048_15_1_O
    );
  rx_input_memio_n0048_12_1 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crc_12_Q,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => VCC,
      O => rx_input_memio_n0048_12_1_O
    );
  rx_input_memio_n0048_31_1 : X_LUT4
    generic map(
      INIT => X"EDDE"
    )
    port map (
      ADR0 => rx_input_memio_crcl(29),
      ADR1 => rx_input_memio_crcrst,
      ADR2 => rx_input_memio_datal(2),
      ADR3 => rx_input_memio_crcl(23),
      O => rx_input_memio_n0048_31_Q
    );
  rx_input_memio_n00341 : X_LUT4
    generic map(
      INIT => X"3330"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_RESET_1,
      ADR2 => rx_input_memio_crcen,
      ADR3 => rx_input_memio_crcrst,
      O => rx_input_memio_crcl_31_GROM
    );
  rx_input_memio_crcl_31_YUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_31_GROM,
      O => rx_input_memio_n0034
    );
  rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(30),
      ADR1 => rx_input_memio_crcl(4),
      ADR2 => rx_input_memio_datal(1),
      ADR3 => rx_input_memio_crccomb_n0115(0),
      O => rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O_FROM
    );
  rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0118(0),
      ADR1 => rx_input_memio_crccomb_Mxor_CO_23_Xo(0),
      ADR2 => rx_input_memio_crccomb_n0118(1),
      ADR3 => rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O,
      O => rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O_FROM,
      O => rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O
    );
  rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_12_Xo_3_1_SW0_O_GROM,
      O => rx_input_memio_crc_12_Q
    );
  rx_input_memio_cs_FFd15_In6 : X_LUT4
    generic map(
      INIT => X"F800"
    )
    port map (
      ADR0 => rx_input_memio_n0016,
      ADR1 => rx_input_memio_cs_FFd16_1,
      ADR2 => rx_input_memio_cs_FFd10,
      ADR3 => rx_input_memio_brdy,
      O => rx_input_memio_cs_FFd15_FROM
    );
  rx_input_memio_cs_FFd15_In7 : X_LUT4
    generic map(
      INIT => X"FF88"
    )
    port map (
      ADR0 => rx_input_invalid,
      ADR1 => rx_input_memio_cs_FFd15,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd15_In6_O,
      O => rx_input_memio_cs_FFd15_In7_O
    );
  rx_input_memio_cs_FFd15_XUSED : X_BUF
    port map (
      I => rx_input_memio_cs_FFd15_FROM,
      O => rx_input_memio_cs_FFd15_In6_O
    );
  rx_input_memio_cs_Out910 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd8,
      ADR1 => rx_input_memio_cs_FFd13,
      ADR2 => rx_input_memio_cs_FFd15,
      ADR3 => rx_input_memio_cs_FFd16_1,
      O => rx_input_memio_menl_FROM
    );
  rx_input_memio_cs_Out917 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd7,
      ADR1 => rx_input_memio_cs_FFd6,
      ADR2 => rx_input_memio_N80990,
      ADR3 => rx_input_memio_cs_Out910_O,
      O => rx_input_memio_menl_GROM
    );
  rx_input_memio_menl_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_menl_CEMUXNOT
    );
  rx_input_memio_menl_XUSED : X_BUF
    port map (
      I => rx_input_memio_menl_FROM,
      O => rx_input_memio_cs_Out910_O
    );
  rx_input_memio_menl_YUSED : X_BUF
    port map (
      I => rx_input_memio_menl_GROM,
      O => rx_input_memio_men
    );
  mac_control_PHY_status_n0019_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => mac_control_PHY_status_cs_FFd5,
      ADR2 => mac_control_PHY_status_cs_FFd2,
      ADR3 => mac_control_PHY_status_cs_FFd4,
      O => mac_control_PHY_status_n0019_SW0_O_FROM
    );
  mac_control_PHY_status_n0019_1578 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => mac_control_PHY_status_done,
      ADR1 => mac_control_PHY_status_cs_FFd6,
      ADR2 => mac_control_PHY_status_cs_FFd3,
      ADR3 => mac_control_PHY_status_n0019_SW0_O,
      O => mac_control_PHY_status_n0019_SW0_O_GROM
    );
  mac_control_PHY_status_n0019_SW0_O_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_n0019_SW0_O_FROM,
      O => mac_control_PHY_status_n0019_SW0_O
    );
  mac_control_PHY_status_n0019_SW0_O_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_n0019_SW0_O_GROM,
      O => mac_control_PHY_status_n0019
    );
  rx_input_memio_crccomb_Mxor_n0009_Result1 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_input_memio_crcl(28),
      ADR1 => rx_input_memio_datal(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_crccomb_n0115_0_FROM
    );
  rx_input_memio_crccomb_Mxor_CO_15_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(7),
      ADR1 => rx_input_memio_crccomb_n0118(0),
      ADR2 => rx_input_memio_crccomb_Mxor_CO_13_Xo(2),
      ADR3 => rx_input_memio_crccomb_n0115(0),
      O => rx_input_memio_crccomb_n0115_0_GROM
    );
  rx_input_memio_crccomb_n0115_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_n0115_0_FROM,
      O => rx_input_memio_crccomb_n0115(0)
    );
  rx_input_memio_crccomb_n0115_0_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_n0115_0_GROM,
      O => rx_input_memio_crc_15_Q
    );
  tx_input_Ker3585921 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => tx_input_CNT(8),
      ADR1 => tx_input_CNT(9),
      ADR2 => tx_input_CNT(10),
      ADR3 => tx_input_CNT(11),
      O => tx_input_Ker3585921_O_FROM
    );
  tx_input_Ker3585927 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_CHOICE1998,
      ADR2 => VCC,
      ADR3 => tx_input_Ker3585921_O,
      O => tx_input_Ker3585921_O_GROM
    );
  tx_input_Ker3585921_O_XUSED : X_BUF
    port map (
      I => tx_input_Ker3585921_O_FROM,
      O => tx_input_Ker3585921_O
    );
  tx_input_Ker3585921_O_YUSED : X_BUF
    port map (
      I => tx_input_Ker3585921_O_GROM,
      O => tx_input_CHOICE1999
    );
  rx_input_fifo_control_ldata_8_10 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_control_CHOICE1605,
      ADR2 => rx_input_fifo_control_CHOICE1602,
      ADR3 => VCC,
      O => rx_input_fifo_control_ldata(8)
    );
  rx_input_fifo_control_n00081 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => RESET_IBUF_2,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_ce,
      O => rx_input_endf_GROM
    );
  rx_input_endf_YUSED : X_BUF
    port map (
      I => rx_input_endf_GROM,
      O => rx_input_fifo_control_n0008
    );
  tx_output_n0034_15_1 : X_LUT4
    generic map(
      INIT => X"FAFA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => tx_output_crc_15_Q,
      ADR3 => VCC,
      O => tx_output_n0034_15_1_O
    );
  tx_output_n0034_5_1 : X_LUT4
    generic map(
      INIT => X"FAFA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => tx_output_crc_5_Q,
      ADR3 => VCC,
      O => tx_output_n0034_5_1_O
    );
  tx_input_Ker35859120 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => tx_input_N80947,
      ADR1 => tx_input_CHOICE2014,
      ADR2 => tx_input_CHOICE2029,
      ADR3 => tx_input_CHOICE2022,
      O => tx_input_Ker35859120_O_FROM
    );
  tx_input_Ker35859137 : X_LUT4
    generic map(
      INIT => X"FF80"
    )
    port map (
      ADR0 => tx_input_CHOICE1991,
      ADR1 => tx_input_CHOICE1988,
      ADR2 => tx_input_CHOICE1999,
      ADR3 => tx_input_Ker35859120_O,
      O => tx_input_Ker35859120_O_GROM
    );
  tx_input_Ker35859120_O_XUSED : X_BUF
    port map (
      I => tx_input_Ker35859120_O_FROM,
      O => tx_input_Ker35859120_O
    );
  tx_input_Ker35859120_O_YUSED : X_BUF
    port map (
      I => tx_input_Ker35859120_O_GROM,
      O => tx_input_N35861
    );
  rx_input_memio_n0048_22_1 : X_LUT4
    generic map(
      INIT => X"FF96"
    )
    port map (
      ADR0 => rx_input_memio_datal(7),
      ADR1 => rx_input_memio_crcl(24),
      ADR2 => rx_input_memio_crcl(14),
      ADR3 => rx_input_memio_crcrst,
      O => rx_input_memio_n0048_22_Q
    );
  rx_input_memio_n0048_5_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_5_Q,
      O => rx_input_memio_n0048_5_1_O
    );
  tx_output_crc_loigc_Mxor_n0005_Result1 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => tx_output_data(3),
      ADR1 => VCC,
      ADR2 => tx_output_crcl(28),
      ADR3 => tx_output_crc_0_Q,
      O => tx_output_crc_loigc_Mxor_n0005_Result1_O_FROM
    );
  tx_output_crc_loigc_Mxor_CO_5_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0124(1),
      ADR1 => tx_output_crc_loigc_Mxor_n0007_Xo(0),
      ADR2 => tx_output_crc_loigc_n0124(0),
      ADR3 => tx_output_crc_loigc_Mxor_n0005_Result1_O,
      O => tx_output_crc_loigc_Mxor_n0005_Result1_O_GROM
    );
  tx_output_crc_loigc_Mxor_n0005_Result1_O_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_n0005_Result1_O_FROM,
      O => tx_output_crc_loigc_Mxor_n0005_Result1_O
    );
  tx_output_crc_loigc_Mxor_n0005_Result1_O_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_n0005_Result1_O_GROM,
      O => tx_output_crc_5_Q
    );
  rx_output_n0046_10_SW0 : X_LUT4
    generic map(
      INIT => X"4747"
    )
    port map (
      ADR0 => rx_output_n0070(10),
      ADR1 => rx_output_len(1),
      ADR2 => rx_output_len(10),
      ADR3 => VCC,
      O => rx_output_lenr_10_FROM
    );
  rx_output_n0046_10_Q : X_LUT4
    generic map(
      INIT => X"C0CF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_n0060(10),
      ADR2 => rx_output_len(0),
      ADR3 => rx_output_n0046_10_SW0_O,
      O => rx_output_n0046_10_O
    );
  rx_output_lenr_10_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_10_CEMUXNOT
    );
  rx_output_lenr_10_XUSED : X_BUF
    port map (
      I => rx_output_lenr_10_FROM,
      O => rx_output_n0046_10_SW0_O
    );
  mac_control_PHY_status_MII_Interface_cs_FFd2_1579 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd2_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_cs_FFd2_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_cs_FFd2
    );
  mac_control_PHY_status_MII_Interface_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_MII_Interface_cs_FFd2_FFY_RST
    );
  rx_output_n0046_11_SW0 : X_LUT4
    generic map(
      INIT => X"505F"
    )
    port map (
      ADR0 => rx_output_n0070(11),
      ADR1 => VCC,
      ADR2 => rx_output_len(1),
      ADR3 => rx_output_len(11),
      O => rx_output_lenr_11_FROM
    );
  rx_output_n0046_11_Q : X_LUT4
    generic map(
      INIT => X"A0F5"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => VCC,
      ADR2 => rx_output_n0060(11),
      ADR3 => rx_output_n0046_11_SW0_O,
      O => rx_output_n0046_11_O
    );
  rx_output_lenr_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_11_CEMUXNOT
    );
  rx_output_lenr_11_XUSED : X_BUF
    port map (
      I => rx_output_lenr_11_FROM,
      O => rx_output_n0046_11_SW0_O
    );
  rx_output_n0046_12_SW0 : X_LUT4
    generic map(
      INIT => X"550F"
    )
    port map (
      ADR0 => rx_output_n0070(12),
      ADR1 => VCC,
      ADR2 => rx_output_len(12),
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_12_FROM
    );
  rx_output_n0046_12_Q : X_LUT4
    generic map(
      INIT => X"88DD"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => rx_output_n0060(12),
      ADR2 => VCC,
      ADR3 => rx_output_n0046_12_SW0_O,
      O => rx_output_n0046_12_O
    );
  rx_output_lenr_12_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_12_CEMUXNOT
    );
  rx_output_lenr_12_XUSED : X_BUF
    port map (
      I => rx_output_lenr_12_FROM,
      O => rx_output_n0046_12_SW0_O
    );
  rx_output_n0046_13_SW0 : X_LUT4
    generic map(
      INIT => X"5353"
    )
    port map (
      ADR0 => rx_output_n0070(13),
      ADR1 => rx_output_len(13),
      ADR2 => rx_output_len(1),
      ADR3 => VCC,
      O => rx_output_lenr_13_FROM
    );
  rx_output_n0046_13_Q : X_LUT4
    generic map(
      INIT => X"C0F3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(0),
      ADR2 => rx_output_n0060(13),
      ADR3 => rx_output_n0046_13_SW0_O,
      O => rx_output_n0046_13_O
    );
  rx_output_lenr_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_13_CEMUXNOT
    );
  rx_output_lenr_13_XUSED : X_BUF
    port map (
      I => rx_output_lenr_13_FROM,
      O => rx_output_n0046_13_SW0_O
    );
  rx_output_n0046_14_SW0 : X_LUT4
    generic map(
      INIT => X"550F"
    )
    port map (
      ADR0 => rx_output_n0070(14),
      ADR1 => VCC,
      ADR2 => rx_output_len(14),
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_14_FROM
    );
  rx_output_n0046_14_Q : X_LUT4
    generic map(
      INIT => X"88DD"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => rx_output_n0060(14),
      ADR2 => VCC,
      ADR3 => rx_output_n0046_14_SW0_O,
      O => rx_output_n0046_14_O
    );
  rx_output_lenr_14_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_14_CEMUXNOT
    );
  rx_output_lenr_14_XUSED : X_BUF
    port map (
      I => rx_output_lenr_14_FROM,
      O => rx_output_n0046_14_SW0_O
    );
  rx_output_n0046_15_SW0 : X_LUT4
    generic map(
      INIT => X"550F"
    )
    port map (
      ADR0 => rx_output_n0070(15),
      ADR1 => VCC,
      ADR2 => rx_output_len(15),
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_15_FROM
    );
  rx_output_n0046_15_Q : X_LUT4
    generic map(
      INIT => X"A0F5"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => VCC,
      ADR2 => rx_output_n0060(15),
      ADR3 => rx_output_n0046_15_SW0_O,
      O => rx_output_n0046_15_O
    );
  rx_output_lenr_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_15_CEMUXNOT
    );
  rx_output_lenr_15_XUSED : X_BUF
    port map (
      I => rx_output_lenr_15_FROM,
      O => rx_output_n0046_15_SW0_O
    );
  tx_input_Ker358701 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => RESET_IBUF_1,
      ADR1 => VCC,
      ADR2 => tx_input_den,
      ADR3 => VCC,
      O => tx_input_N35872_FROM
    );
  tx_input_n00201 : X_LUT4
    generic map(
      INIT => X"FE00"
    )
    port map (
      ADR0 => tx_input_cs_FFd11,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => tx_input_cs_FFd10,
      ADR3 => tx_input_N35872,
      O => tx_input_N35872_GROM
    );
  tx_input_N35872_XUSED : X_BUF
    port map (
      I => tx_input_N35872_FROM,
      O => tx_input_N35872
    );
  tx_input_N35872_YUSED : X_BUF
    port map (
      I => tx_input_N35872_GROM,
      O => tx_input_n0020
    );
  tx_output_crc_loigc_Mxor_CO_0_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(1),
      ADR1 => tx_output_crcl(30),
      ADR2 => tx_output_crcl(24),
      ADR3 => tx_output_data(7),
      O => tx_output_crc_0_FROM
    );
  tx_output_crc_loigc_Mxor_CO_1_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(0),
      ADR1 => tx_output_crc_0_Q,
      ADR2 => tx_output_crc_loigc_n0122(0),
      ADR3 => tx_output_crcl(31),
      O => tx_output_crc_0_GROM
    );
  tx_output_crc_0_XUSED : X_BUF
    port map (
      I => tx_output_crc_0_FROM,
      O => tx_output_crc_0_Q
    );
  tx_output_crc_0_YUSED : X_BUF
    port map (
      I => tx_output_crc_0_GROM,
      O => tx_output_crc_1_Q
    );
  rx_output_n0046_2_SW0 : X_LUT4
    generic map(
      INIT => X"303F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_n0070(2),
      ADR2 => rx_output_len(1),
      ADR3 => rx_output_len(2),
      O => rx_output_lenr_2_FROM
    );
  rx_output_n0046_2_Q : X_LUT4
    generic map(
      INIT => X"A0AF"
    )
    port map (
      ADR0 => rx_output_n0060(2),
      ADR1 => VCC,
      ADR2 => rx_output_len(0),
      ADR3 => rx_output_n0046_2_SW0_O,
      O => rx_output_n0046_2_O
    );
  rx_output_lenr_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_2_CEMUXNOT
    );
  rx_output_lenr_2_XUSED : X_BUF
    port map (
      I => rx_output_lenr_2_FROM,
      O => rx_output_n0046_2_SW0_O
    );
  rx_output_n0046_3_SW0 : X_LUT4
    generic map(
      INIT => X"0F33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(3),
      ADR2 => rx_output_n0070(3),
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_3_FROM
    );
  rx_output_n0046_3_Q : X_LUT4
    generic map(
      INIT => X"88BB"
    )
    port map (
      ADR0 => rx_output_n0060(3),
      ADR1 => rx_output_len(0),
      ADR2 => VCC,
      ADR3 => rx_output_n0046_3_SW0_O,
      O => rx_output_n0046_3_O
    );
  rx_output_lenr_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_3_CEMUXNOT
    );
  rx_output_lenr_3_XUSED : X_BUF
    port map (
      I => rx_output_lenr_3_FROM,
      O => rx_output_n0046_3_SW0_O
    );
  rx_output_n0046_4_SW0 : X_LUT4
    generic map(
      INIT => X"550F"
    )
    port map (
      ADR0 => rx_output_n0070(4),
      ADR1 => VCC,
      ADR2 => rx_output_len(4),
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_4_FROM
    );
  rx_output_n0046_4_Q : X_LUT4
    generic map(
      INIT => X"88DD"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => rx_output_n0060(4),
      ADR2 => VCC,
      ADR3 => rx_output_n0046_4_SW0_O,
      O => rx_output_n0046_4_O
    );
  rx_output_lenr_4_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_4_CEMUXNOT
    );
  rx_output_lenr_4_XUSED : X_BUF
    port map (
      I => rx_output_lenr_4_FROM,
      O => rx_output_n0046_4_SW0_O
    );
  rx_output_n0046_5_SW0 : X_LUT4
    generic map(
      INIT => X"0C3F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_len(1),
      ADR2 => rx_output_n0070(5),
      ADR3 => rx_output_len(5),
      O => rx_output_lenr_5_FROM
    );
  rx_output_n0046_5_Q : X_LUT4
    generic map(
      INIT => X"C0CF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_n0060(5),
      ADR2 => rx_output_len(0),
      ADR3 => rx_output_n0046_5_SW0_O,
      O => rx_output_n0046_5_O
    );
  rx_output_lenr_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_5_CEMUXNOT
    );
  rx_output_lenr_5_XUSED : X_BUF
    port map (
      I => rx_output_lenr_5_FROM,
      O => rx_output_n0046_5_SW0_O
    );
  tx_output_cs_Out151 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd5,
      ADR1 => tx_output_cs_FFd4,
      ADR2 => tx_output_cs_FFd6,
      ADR3 => tx_output_cs_FFd8,
      O => tx_output_crcenl_FROM
    );
  tx_output_n00331 : X_LUT4
    generic map(
      INIT => X"5544"
    )
    port map (
      ADR0 => RESET_IBUF_2,
      ADR1 => tx_output_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_output_decbcnt,
      O => tx_output_crcenl_GROM
    );
  tx_output_crcenl_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_crcenl_CEMUXNOT
    );
  tx_output_crcenl_XUSED : X_BUF
    port map (
      I => tx_output_crcenl_FROM,
      O => tx_output_decbcnt
    );
  tx_output_crcenl_YUSED : X_BUF
    port map (
      I => tx_output_crcenl_GROM,
      O => tx_output_n0033
    );
  rx_output_n0046_6_SW0 : X_LUT4
    generic map(
      INIT => X"5533"
    )
    port map (
      ADR0 => rx_output_n0070(6),
      ADR1 => rx_output_len(6),
      ADR2 => VCC,
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_6_FROM
    );
  rx_output_n0046_6_Q : X_LUT4
    generic map(
      INIT => X"88DD"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => rx_output_n0060(6),
      ADR2 => VCC,
      ADR3 => rx_output_n0046_6_SW0_O,
      O => rx_output_n0046_6_O
    );
  rx_output_lenr_6_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_6_CEMUXNOT
    );
  rx_output_lenr_6_XUSED : X_BUF
    port map (
      I => rx_output_lenr_6_FROM,
      O => rx_output_n0046_6_SW0_O
    );
  mac_control_MACADDR_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_1_FFY_RST,
      O => macaddr(0)
    );
  macaddr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_1_FFY_RST
    );
  rx_output_n0046_7_SW0 : X_LUT4
    generic map(
      INIT => X"0F55"
    )
    port map (
      ADR0 => rx_output_len(7),
      ADR1 => VCC,
      ADR2 => rx_output_n0070(7),
      ADR3 => rx_output_len(1),
      O => rx_output_lenr_7_FROM
    );
  rx_output_n0046_7_Q : X_LUT4
    generic map(
      INIT => X"C0CF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_n0060(7),
      ADR2 => rx_output_len(0),
      ADR3 => rx_output_n0046_7_SW0_O,
      O => rx_output_n0046_7_O
    );
  rx_output_lenr_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_7_CEMUXNOT
    );
  rx_output_lenr_7_XUSED : X_BUF
    port map (
      I => rx_output_lenr_7_FROM,
      O => rx_output_n0046_7_SW0_O
    );
  rx_output_n0046_8_SW0 : X_LUT4
    generic map(
      INIT => X"505F"
    )
    port map (
      ADR0 => rx_output_n0070(8),
      ADR1 => VCC,
      ADR2 => rx_output_len(1),
      ADR3 => rx_output_len(8),
      O => rx_output_lenr_8_FROM
    );
  rx_output_n0046_8_Q : X_LUT4
    generic map(
      INIT => X"88DD"
    )
    port map (
      ADR0 => rx_output_len(0),
      ADR1 => rx_output_n0060(8),
      ADR2 => VCC,
      ADR3 => rx_output_n0046_8_SW0_O,
      O => rx_output_n0046_8_O
    );
  rx_output_lenr_8_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_8_CEMUXNOT
    );
  rx_output_lenr_8_XUSED : X_BUF
    port map (
      I => rx_output_lenr_8_FROM,
      O => rx_output_n0046_8_SW0_O
    );
  rx_output_n0046_9_SW0 : X_LUT4
    generic map(
      INIT => X"0A5F"
    )
    port map (
      ADR0 => rx_output_len(1),
      ADR1 => VCC,
      ADR2 => rx_output_n0070(9),
      ADR3 => rx_output_len(9),
      O => rx_output_lenr_9_FROM
    );
  rx_output_n0046_9_Q : X_LUT4
    generic map(
      INIT => X"88BB"
    )
    port map (
      ADR0 => rx_output_n0060(9),
      ADR1 => rx_output_len(0),
      ADR2 => VCC,
      ADR3 => rx_output_n0046_9_SW0_O,
      O => rx_output_n0046_9_O
    );
  rx_output_lenr_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_lenr_9_CEMUXNOT
    );
  rx_output_lenr_9_XUSED : X_BUF
    port map (
      I => rx_output_lenr_9_FROM,
      O => rx_output_n0046_9_SW0_O
    );
  rx_input_memio_n001618 : X_LUT4
    generic map(
      INIT => X"0040"
    )
    port map (
      ADR0 => rx_input_data(3),
      ADR1 => rx_input_data(0),
      ADR2 => rx_input_data(2),
      ADR3 => rx_input_data(1),
      O => rx_input_memio_n001618_O_FROM
    );
  rx_input_memio_n001619 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_CHOICE1979,
      ADR2 => VCC,
      ADR3 => rx_input_memio_n001618_O,
      O => rx_input_memio_n001618_O_GROM
    );
  rx_input_memio_n001618_O_XUSED : X_BUF
    port map (
      I => rx_input_memio_n001618_O_FROM,
      O => rx_input_memio_n001618_O
    );
  rx_input_memio_n001618_O_YUSED : X_BUF
    port map (
      I => rx_input_memio_n001618_O_GROM,
      O => rx_input_memio_n0016
    );
  rx_output_n0043_SW1 : X_LUT4
    generic map(
      INIT => X"0005"
    )
    port map (
      ADR0 => rx_output_cs_FFd17,
      ADR1 => VCC,
      ADR2 => rx_output_cs_FFd5,
      ADR3 => rx_output_cs_FFd11,
      O => rx_output_n0043_SW1_O_FROM
    );
  rx_output_n0043_1580 : X_LUT4
    generic map(
      INIT => X"3233"
    )
    port map (
      ADR0 => rx_output_cs_FFd1,
      ADR1 => RESET_IBUF,
      ADR2 => rx_output_cs_FFd19,
      ADR3 => rx_output_n0043_SW1_O,
      O => rx_output_n0043_SW1_O_GROM
    );
  rx_output_n0043_SW1_O_XUSED : X_BUF
    port map (
      I => rx_output_n0043_SW1_O_FROM,
      O => rx_output_n0043_SW1_O
    );
  rx_output_n0043_SW1_O_YUSED : X_BUF
    port map (
      I => rx_output_n0043_SW1_O_GROM,
      O => rx_output_n0043
    );
  mac_control_n00851 : X_LUT4
    generic map(
      INIT => X"0A00"
    )
    port map (
      ADR0 => mac_control_addr(3),
      ADR1 => VCC,
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_N53132,
      O => mac_control_n0085_FROM
    );
  mac_control_n00421 : X_LUT4
    generic map(
      INIT => X"F5FF"
    )
    port map (
      ADR0 => mac_control_sclkdeltal,
      ADR1 => VCC,
      ADR2 => mac_control_addr(7),
      ADR3 => mac_control_n0085,
      O => mac_control_n0085_GROM
    );
  mac_control_n0085_XUSED : X_BUF
    port map (
      I => mac_control_n0085_FROM,
      O => mac_control_n0085
    );
  mac_control_n0085_YUSED : X_BUF
    port map (
      I => mac_control_n0085_GROM,
      O => mac_control_PHY_status_n00181_O
    );
  tx_input_cs_FFd6_In1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => tx_input_den,
      ADR1 => VCC,
      ADR2 => tx_input_cs_FFd7,
      ADR3 => VCC,
      O => tx_input_cs_FFd6_In
    );
  tx_input_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"FCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_cs_FFd4,
      ADR2 => tx_input_N35861,
      ADR3 => tx_input_cs_FFd6,
      O => tx_input_cs_FFd5_In1_O
    );
  mac_control_MACADDR_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_1_FFX_RST,
      O => macaddr(1)
    );
  macaddr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_1_FFX_RST
    );
  tx_input_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_input_N35861,
      ADR3 => tx_input_cs_FFd9,
      O => tx_input_cs_FFd8_In1_O
    );
  tx_input_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"4F44"
    )
    port map (
      ADR0 => tx_input_den,
      ADR1 => tx_input_cs_FFd7,
      ADR2 => tx_input_N35861,
      ADR3 => tx_input_cs_FFd9,
      O => tx_input_cs_FFd7_In1_O
    );
  rx_input_memio_crccomb_Mxor_CO_0_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_datal(7),
      ADR1 => rx_input_memio_crcl(30),
      ADR2 => rx_input_memio_crcl(24),
      ADR3 => rx_input_memio_datal(1),
      O => rx_input_memio_crc_0_FROM
    );
  rx_input_memio_crccomb_Mxor_CO_1_Result1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(31),
      ADR1 => rx_input_memio_crccomb_n0122(0),
      ADR2 => rx_input_memio_datal(0),
      ADR3 => rx_input_memio_crc_0_Q,
      O => rx_input_memio_crc_0_GROM
    );
  rx_input_memio_crc_0_XUSED : X_BUF
    port map (
      I => rx_input_memio_crc_0_FROM,
      O => rx_input_memio_crc_0_Q
    );
  rx_input_memio_crc_0_YUSED : X_BUF
    port map (
      I => rx_input_memio_crc_0_GROM,
      O => rx_input_memio_crc_1_Q
    );
  rx_input_memio_cs_Out8 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd14,
      ADR1 => rx_input_memio_cs_FFd12,
      ADR2 => rx_input_memio_N70855,
      ADR3 => rx_input_memio_cs_FFd16_1,
      O => rx_input_fifo_rd_en_FROM
    );
  rx_input_memio_n01021 : X_LUT4
    generic map(
      INIT => X"CDCC"
    )
    port map (
      ADR0 => rx_input_invalid,
      ADR1 => rx_input_memio_cs_FFd16,
      ADR2 => rx_input_endf,
      ADR3 => rx_input_ce,
      O => rx_input_fifo_rd_en_GROM
    );
  rx_input_fifo_rd_en_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_rd_en_CEMUXNOT
    );
  rx_input_fifo_rd_en_XUSED : X_BUF
    port map (
      I => rx_input_fifo_rd_en_FROM,
      O => rx_input_ce
    );
  rx_input_fifo_rd_en_YUSED : X_BUF
    port map (
      I => rx_input_fifo_rd_en_GROM,
      O => rx_input_memio_n0102
    );
  mac_control_PHY_status_n00171 : X_LUT4
    generic map(
      INIT => X"0F05"
    )
    port map (
      ADR0 => mac_control_PHY_status_n00181_O,
      ADR1 => VCC,
      ADR2 => RESET_IBUF,
      ADR3 => mac_control_PHY_status_cs_FFd1,
      O => mac_control_phyaddr_31_GROM
    );
  mac_control_phyaddr_31_YUSED : X_BUF
    port map (
      I => mac_control_phyaddr_31_GROM,
      O => mac_control_PHY_status_n00171_O
    );
  tx_output_addrinc_SW0 : X_LUT4
    generic map(
      INIT => X"EEEE"
    )
    port map (
      ADR0 => tx_output_cs_FFd16,
      ADR1 => tx_output_cs_FFd7,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_output_addrinc_SW0_O_FROM
    );
  tx_output_addrinc_1581 : X_LUT4
    generic map(
      INIT => X"FEFC"
    )
    port map (
      ADR0 => tx_output_cs_FFd8,
      ADR1 => tx_output_addrinc_SW0_O,
      ADR2 => tx_output_cs_FFd12,
      ADR3 => tx_output_n0035,
      O => tx_output_addrinc_SW0_O_GROM
    );
  tx_output_addrinc_SW0_O_XUSED : X_BUF
    port map (
      I => tx_output_addrinc_SW0_O_FROM,
      O => tx_output_addrinc_SW0_O
    );
  tx_output_addrinc_SW0_O_YUSED : X_BUF
    port map (
      I => tx_output_addrinc_SW0_O_GROM,
      O => tx_output_addrinc
    );
  tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(1),
      ADR1 => tx_output_crcl(30),
      ADR2 => tx_output_crcl(4),
      ADR3 => tx_output_crc_loigc_n0115(0),
      O => tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O_FROM
    );
  tx_output_crc_loigc_Mxor_CO_12_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0118(1),
      ADR1 => tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O,
      ADR2 => tx_output_crc_loigc_Mxor_CO_23_Xo(0),
      ADR3 => tx_output_crc_loigc_n0118(0),
      O => tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O_GROM
    );
  tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O_XUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O_FROM,
      O => tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O
    );
  tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O_YUSED : X_BUF
    port map (
      I => tx_output_crc_loigc_Mxor_CO_12_Xo_3_1_SW0_O_GROM,
      O => tx_output_crc_12_Q
    );
  rx_input_memio_crccomb_Mxor_n0005_Result1 : X_LUT4
    generic map(
      INIT => X"C33C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_datal(3),
      ADR2 => rx_input_memio_crcl(28),
      ADR3 => rx_input_memio_crc_0_Q,
      O => rx_input_memio_crccomb_Mxor_n0005_Result1_O_FROM
    );
  rx_input_memio_crccomb_Mxor_CO_5_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0124(0),
      ADR1 => rx_input_memio_crccomb_n0124(1),
      ADR2 => rx_input_memio_crccomb_Mxor_n0007_Xo(0),
      ADR3 => rx_input_memio_crccomb_Mxor_n0005_Result1_O,
      O => rx_input_memio_crccomb_Mxor_n0005_Result1_O_GROM
    );
  rx_input_memio_crccomb_Mxor_n0005_Result1_O_XUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_n0005_Result1_O_FROM,
      O => rx_input_memio_crccomb_Mxor_n0005_Result1_O
    );
  rx_input_memio_crccomb_Mxor_n0005_Result1_O_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_n0005_Result1_O_GROM,
      O => rx_input_memio_crc_5_Q
    );
  mac_control_n00461 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => mac_control_N53194,
      ADR1 => mac_control_din(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_n0046
    );
  mac_control_n00481 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => mac_control_N53194,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_din(2),
      O => mac_control_n0048
    );
  mac_control_txf_rst_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_rst_CEMUXNOT
    );
  rx_input_memio_addrchk_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"00E4"
    )
    port map (
      ADR0 => rx_input_memio_brdy,
      ADR1 => rx_input_memio_addrchk_cs_FFd4,
      ADR2 => rx_input_memio_addrchk_cs_FFd5,
      ADR3 => rx_input_memio_cs_FFd16_1,
      O => rx_input_memio_addrchk_cs_FFd4_In
    );
  rx_input_memio_addrchk_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"00E4"
    )
    port map (
      ADR0 => rx_input_memio_brdy,
      ADR1 => rx_input_memio_addrchk_cs_FFd3,
      ADR2 => rx_input_memio_addrchk_cs_FFd4,
      ADR3 => rx_input_memio_cs_FFd16_1,
      O => rx_input_memio_addrchk_cs_FFd3_In
    );
  rx_input_memio_cs_FFd10_In1 : X_LUT4
    generic map(
      INIT => X"DC10"
    )
    port map (
      ADR0 => rx_input_endf,
      ADR1 => rx_input_invalid,
      ADR2 => rx_input_memio_cs_FFd12,
      ADR3 => rx_input_memio_cs_FFd10,
      O => rx_input_memio_cs_FFd10_In
    );
  rx_input_memio_cs_FFd9_In1 : X_LUT4
    generic map(
      INIT => X"FF08"
    )
    port map (
      ADR0 => rx_input_endf,
      ADR1 => rx_input_memio_cs_FFd12,
      ADR2 => rx_input_invalid,
      ADR3 => rx_input_memio_cs_FFd11,
      O => rx_input_memio_cs_FFd9_In
    );
  mac_control_PHY_status_MII_Interface_n0014_1_1 : X_LUT4
    generic map(
      INIT => X"4404"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR1 => mac_control_PHY_status_MII_Interface_n0076(1),
      ADR2 => mac_control_PHY_status_MII_Interface_N38617,
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE1101,
      O => mac_control_PHY_status_MII_Interface_n0014(1)
    );
  mac_control_PHY_status_MII_Interface_n0014_0_1 : X_LUT4
    generic map(
      INIT => X"000F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      O => mac_control_PHY_status_MII_Interface_n0014(0)
    );
  mac_control_PHY_status_MII_Interface_n0014_3_1 : X_LUT4
    generic map(
      INIT => X"00D0"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_N38617,
      ADR1 => mac_control_PHY_status_MII_Interface_CHOICE1101,
      ADR2 => mac_control_PHY_status_MII_Interface_n0076(3),
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      O => mac_control_PHY_status_MII_Interface_n0014(3)
    );
  mac_control_PHY_status_MII_Interface_n0014_2_1 : X_LUT4
    generic map(
      INIT => X"3100"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_N38617,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR2 => mac_control_PHY_status_MII_Interface_CHOICE1101,
      ADR3 => mac_control_PHY_status_MII_Interface_n0076(2),
      O => mac_control_PHY_status_MII_Interface_n0014(2)
    );
  mac_control_PHY_status_MII_Interface_n0014_5_1 : X_LUT4
    generic map(
      INIT => X"0A02"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_n0076(5),
      ADR1 => mac_control_PHY_status_MII_Interface_N38617,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE1101,
      O => mac_control_PHY_status_MII_Interface_n0014(5)
    );
  mac_control_PHY_status_MII_Interface_n0014_4_1 : X_LUT4
    generic map(
      INIT => X"2030"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_CHOICE1101,
      ADR1 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      ADR2 => mac_control_PHY_status_MII_Interface_n0076(4),
      ADR3 => mac_control_PHY_status_MII_Interface_N38617,
      O => mac_control_PHY_status_MII_Interface_n0014(4)
    );
  mac_control_MACADDR_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_3_FFX_RST,
      O => macaddr(3)
    );
  macaddr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_3_FFX_RST
    );
  rx_input_memio_Mmux_lma_Result_1_1 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_71,
      ADR3 => rx_input_memio_bpl(1),
      O => rx_input_memio_lma(1)
    );
  rx_input_memio_Mmux_lma_Result_0_1 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_70,
      ADR3 => rx_input_memio_bpl(0),
      O => rx_input_memio_lma(0)
    );
  rx_input_memio_Mmux_lma_Result_3_1 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => rx_input_memio_macnt_73,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bpl(3),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(3)
    );
  rx_input_memio_Mmux_lma_Result_2_1 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => rx_input_memio_macnt_72,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bpl(2),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(2)
    );
  mac_control_PHY_status_MII_Interface_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"FE00"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd8,
      ADR1 => mac_control_PHY_status_cs_FFd3,
      ADR2 => mac_control_PHY_status_cs_FFd6,
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd6,
      O => mac_control_PHY_status_MII_Interface_cs_FFd5_In
    );
  mac_control_PHY_status_MII_Interface_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"FFD0"
    )
    port map (
      ADR0 => MDC_OBUF,
      ADR1 => mac_control_PHY_status_MII_Interface_mdccnt_37,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd4,
      ADR3 => mac_control_PHY_status_MII_Interface_cs_FFd5,
      O => mac_control_PHY_status_MII_Interface_cs_FFd4_In
    );
  rx_input_memio_Mmux_lma_Result_5_1 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bpl(5),
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_75,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(5)
    );
  rx_input_memio_Mmux_lma_Result_4_1 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => rx_input_memio_macnt_74,
      ADR1 => rx_input_memio_wbpl,
      ADR2 => rx_input_memio_bpl(4),
      ADR3 => VCC,
      O => rx_input_memio_lma(4)
    );
  rx_input_memio_Mmux_lma_Result_7_1 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bpl(7),
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_77,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(7)
    );
  rx_input_memio_Mmux_lma_Result_6_1 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => rx_input_memio_macnt_76,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bpl(6),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(6)
    );
  rx_input_memio_Mmux_lma_Result_9_1 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_79,
      ADR3 => rx_input_memio_bpl(9),
      O => rx_input_memio_lma(9)
    );
  rx_input_memio_Mmux_lma_Result_8_1 : X_LUT4
    generic map(
      INIT => X"F3C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_wbpl,
      ADR2 => rx_input_memio_bpl(8),
      ADR3 => rx_input_memio_macnt_78,
      O => rx_input_memio_lma(8)
    );
  rx_input_memio_Mmux_lmd_Result_15_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_bcntl(15),
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(15),
      O => rx_input_memio_lmd(15)
    );
  rx_input_memio_Mmux_lmd_Result_0_1 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcntl(0),
      ADR3 => rx_input_memio_doutl(0),
      O => rx_input_memio_lmd(0)
    );
  rx_input_memio_Mmux_lmd_Result_14_1 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => rx_input_memio_doutl(14),
      ADR1 => rx_input_memio_wbpl,
      ADR2 => rx_input_memio_bcntl(14),
      ADR3 => VCC,
      O => rx_input_memio_lmd(14)
    );
  rx_input_memio_Mmux_lmd_Result_1_1 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(1),
      ADR1 => rx_input_memio_wbpl,
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(1),
      O => rx_input_memio_lmd(1)
    );
  rx_input_memio_Mmux_lmd_Result_3_1 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(3),
      ADR1 => rx_input_memio_doutl(3),
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lmd(3)
    );
  rx_input_memio_Mmux_lmd_Result_2_1 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_bcntl(2),
      ADR2 => rx_input_memio_doutl(2),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(2)
    );
  rx_input_memio_Mmux_lmd_Result_5_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_bcntl(5),
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(5),
      O => rx_input_memio_lmd(5)
    );
  rx_input_memio_Mmux_lmd_Result_4_1 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcntl(4),
      ADR3 => rx_input_memio_doutl(4),
      O => rx_input_memio_lmd(4)
    );
  rx_input_memio_Mmux_lmd_Result_7_1 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bcntl(7),
      ADR3 => rx_input_memio_doutl(7),
      O => rx_input_memio_lmd(7)
    );
  rx_input_memio_Mmux_lmd_Result_6_1 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(6),
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(6),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(6)
    );
  mac_control_MACADDR_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_5_FFX_RST,
      O => macaddr(5)
    );
  macaddr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_5_FFX_RST
    );
  rx_input_memio_Mmux_lmd_Result_9_1 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => rx_input_memio_doutl(9),
      ADR1 => rx_input_memio_bcntl(9),
      ADR2 => VCC,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(9)
    );
  rx_input_memio_Mmux_lmd_Result_8_1 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(8),
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(8),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(8)
    );
  mac_control_MACADDR_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_7_FFY_RST,
      O => macaddr(6)
    );
  macaddr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_7_FFY_RST
    );
  rx_input_memio_n0048_21_1 : X_LUT4
    generic map(
      INIT => X"EBBE"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => rx_input_memio_crcl(29),
      ADR2 => rx_input_memio_datal(2),
      ADR3 => rx_input_memio_crcl(13),
      O => rx_input_memio_n0048_21_Q
    );
  rx_input_memio_n0048_20_1 : X_LUT4
    generic map(
      INIT => X"EBBE"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => rx_input_memio_crcl(28),
      ADR2 => rx_input_memio_datal(3),
      ADR3 => rx_input_memio_crcl(12),
      O => rx_input_memio_n0048_20_Q
    );
  memcontroller_clknum_1_2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_1_2_FFY_RST
    );
  memcontroller_clknum_1_1_1582 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_1_2_GROM,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_clknum_1_2_FFY_RST,
      O => memcontroller_clknum_1_1
    );
  memcontroller_n01491 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_0_1,
      ADR3 => memcontroller_clknum_1_2,
      O => memcontroller_clknum_1_2_GROM
    );
  memcontroller_clknum_1_2_YUSED : X_BUF
    port map (
      I => memcontroller_clknum_1_2_GROM,
      O => memcontroller_n0149
    );
  rx_input_memio_cs_FFd12_In1 : X_LUT4
    generic map(
      INIT => X"CE02"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd14,
      ADR1 => rx_input_invalid,
      ADR2 => rx_input_endf,
      ADR3 => rx_input_memio_cs_FFd12,
      O => rx_input_memio_cs_FFd12_In
    );
  rx_input_memio_cs_FFd11_In1 : X_LUT4
    generic map(
      INIT => X"4040"
    )
    port map (
      ADR0 => rx_input_invalid,
      ADR1 => rx_input_memio_cs_FFd14,
      ADR2 => rx_input_endf,
      ADR3 => VCC,
      O => rx_input_memio_cs_FFd11_In
    );
  rx_input_memio_cs_FFd14_In1 : X_LUT4
    generic map(
      INIT => X"AE04"
    )
    port map (
      ADR0 => rx_input_invalid,
      ADR1 => rx_input_memio_cs_FFd15,
      ADR2 => rx_input_endf,
      ADR3 => rx_input_memio_cs_FFd14,
      O => rx_input_memio_cs_FFd14_In
    );
  rx_input_memio_cs_FFd13_In1 : X_LUT4
    generic map(
      INIT => X"FF40"
    )
    port map (
      ADR0 => rx_input_invalid,
      ADR1 => rx_input_memio_cs_FFd15,
      ADR2 => rx_input_endf,
      ADR3 => rx_input_memio_cs_FFd8,
      O => rx_input_memio_cs_FFd13_In
    );
  rx_input_memio_cs_FFd16_In13 : X_LUT4
    generic map(
      INIT => X"EFCC"
    )
    port map (
      ADR0 => rx_input_memio_CHOICE1113,
      ADR1 => rx_input_memio_CHOICE1112,
      ADR2 => rx_input_memio_n0016,
      ADR3 => rx_input_memio_cs_FFd16_1,
      O => rx_input_memio_cs_FFd16_1_GROM
    );
  rx_input_memio_cs_FFd16_1_YUSED : X_BUF
    port map (
      I => rx_input_memio_cs_FFd16_1_GROM,
      O => rx_input_memio_cs_FFd16_In
    );
  mac_control_n00491 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => mac_control_N53194,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_din(3),
      O => mac_control_n0049
    );
  mac_control_n00511 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => mac_control_N53194,
      ADR1 => VCC,
      ADR2 => mac_control_din(5),
      ADR3 => VCC,
      O => mac_control_n0051
    );
  mac_control_rxfifowerr_rst_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxfifowerr_rst_CEMUXNOT
    );
  mac_control_n00471 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_din(1),
      ADR3 => mac_control_N53194,
      O => mac_control_n0047
    );
  mac_control_rxf_rst_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_rst_CEMUXNOT
    );
  rx_input_memio_Mmux_lma_Result_11_1 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => rx_input_memio_macnt_81,
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_bpl(11),
      O => rx_input_memio_lma(11)
    );
  rx_input_memio_Mmux_lma_Result_10_1 : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_macnt_80,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_bpl(10),
      O => rx_input_memio_lma(10)
    );
  rx_input_memio_Mmux_lma_Result_13_1 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_macnt_83,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bpl(13),
      O => rx_input_memio_lma(13)
    );
  rx_input_memio_Mmux_lma_Result_12_1 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bpl(12),
      ADR1 => VCC,
      ADR2 => rx_input_memio_macnt_82,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(12)
    );
  rx_input_memio_Mmux_lma_Result_15_1 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_macnt_85,
      ADR2 => VCC,
      ADR3 => rx_input_memio_bpl(15),
      O => rx_input_memio_lma(15)
    );
  rx_input_memio_Mmux_lma_Result_14_1 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => rx_input_memio_macnt_84,
      ADR1 => VCC,
      ADR2 => rx_input_memio_bpl(14),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lma(14)
    );
  mac_control_MACADDR_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_7_FFX_RST,
      O => macaddr(7)
    );
  macaddr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_7_FFX_RST
    );
  rx_input_memio_Mmux_lmd_Result_11_1 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => rx_input_memio_doutl(11),
      ADR1 => rx_input_memio_bcntl(11),
      ADR2 => VCC,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(11)
    );
  rx_input_memio_Mmux_lmd_Result_10_1 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(10),
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(10),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(10)
    );
  rx_input_memio_Mmux_lmd_Result_21_1 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(21),
      O => rx_input_memio_lmd(21)
    );
  rx_input_memio_Mmux_lmd_Result_20_1 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_wbpl,
      ADR2 => rx_input_memio_doutl(20),
      ADR3 => VCC,
      O => rx_input_memio_lmd(20)
    );
  rx_input_memio_Mmux_lmd_Result_13_1 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => rx_input_memio_bcntl(13),
      ADR1 => rx_input_memio_doutl(13),
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lmd(13)
    );
  rx_input_memio_Mmux_lmd_Result_12_1 : X_LUT4
    generic map(
      INIT => X"D8D8"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => rx_input_memio_bcntl(12),
      ADR2 => rx_input_memio_doutl(12),
      ADR3 => VCC,
      O => rx_input_memio_lmd(12)
    );
  rx_input_memio_Mmux_lmd_Result_31_1 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rx_input_memio_doutl(31),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(31)
    );
  rx_input_memio_Mmux_lmd_Result_30_1 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(30),
      O => rx_input_memio_lmd(30)
    );
  rx_input_memio_Mmux_lmd_Result_23_1 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_doutl(23),
      ADR2 => VCC,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(23)
    );
  rx_input_memio_Mmux_lmd_Result_22_1 : X_LUT4
    generic map(
      INIT => X"5500"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(22),
      O => rx_input_memio_lmd(22)
    );
  rx_input_memio_Mmux_lmd_Result_25_1 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_doutl(25),
      O => rx_input_memio_lmd(25)
    );
  rx_input_memio_Mmux_lmd_Result_24_1 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(24),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(24)
    );
  rx_input_memio_Mmux_lmd_Result_17_1 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_doutl(17),
      ADR2 => VCC,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(17)
    );
  rx_input_memio_Mmux_lmd_Result_16_1 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => rx_input_memio_wbpl,
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(16),
      ADR3 => VCC,
      O => rx_input_memio_lmd(16)
    );
  rx_input_memio_Mmux_lmd_Result_27_1 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_wbpl,
      ADR3 => rx_input_memio_doutl(27),
      O => rx_input_memio_lmd(27)
    );
  rx_input_memio_Mmux_lmd_Result_26_1 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_doutl(26),
      ADR2 => rx_input_memio_wbpl,
      ADR3 => VCC,
      O => rx_input_memio_lmd(26)
    );
  rx_input_memio_Mmux_lmd_Result_19_1 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_doutl(19),
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(19)
    );
  rx_input_memio_Mmux_lmd_Result_18_1 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rx_input_memio_doutl(18),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_wbpl,
      O => rx_input_memio_lmd(18)
    );
  rx_input_memio_Mmux_lmd_Result_29_1 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => rx_input_memio_doutl(29),
      ADR1 => rx_input_memio_wbpl,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_lmd(29)
    );
  rx_input_memio_Mmux_lmd_Result_28_1 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_wbpl,
      ADR2 => VCC,
      ADR3 => rx_input_memio_doutl(28),
      O => rx_input_memio_lmd(28)
    );
  rx_output_Mmux_lma_Result_11_1 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => rx_output_mdl(27),
      ADR1 => VCC,
      ADR2 => rx_output_lmasell,
      ADR3 => rx_output_mdl(11),
      O => rx_output_lma(11)
    );
  rx_output_Mmux_lma_Result_10_1 : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_mdl(10),
      ADR2 => rx_output_lmasell,
      ADR3 => rx_output_mdl(26),
      O => rx_output_lma(10)
    );
  rx_output_fifodin_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_11_CEMUXNOT
    );
  mac_control_MACADDR_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_9_FFX_RST,
      O => macaddr(9)
    );
  macaddr_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_9_FFX_RST
    );
  rx_output_Mmux_lma_Result_13_1 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_lmasell,
      ADR2 => rx_output_mdl(13),
      ADR3 => rx_output_mdl(29),
      O => rx_output_lma(13)
    );
  rx_output_Mmux_lma_Result_12_1 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => rx_output_mdl(28),
      ADR1 => rx_output_lmasell,
      ADR2 => VCC,
      ADR3 => rx_output_mdl(12),
      O => rx_output_lma(12)
    );
  rx_output_fifodin_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_13_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_15_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => rx_output_mdl(31),
      ADR2 => VCC,
      ADR3 => rx_output_mdl(15),
      O => rx_output_lma(15)
    );
  rx_output_Mmux_lma_Result_14_1 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => rx_output_lmasell,
      ADR1 => rx_output_mdl(30),
      ADR2 => VCC,
      ADR3 => rx_output_mdl(14),
      O => rx_output_lma(14)
    );
  rx_output_fifodin_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_15_CEMUXNOT
    );
  tx_input_enableintl_LOGIC_ONE_1583 : X_ONE
    port map (
      O => tx_input_enableintl_LOGIC_ONE
    );
  tx_input_srl16_enable_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_21,
      A1 => GLOBAL_LOGIC0_21,
      A2 => GLOBAL_LOGIC1_13,
      A3 => GLOBAL_LOGIC0_21,
      D => tx_input_enable,
      CE => tx_input_enableintl_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_enableintl_GSHIFT
    );
  tx_input_enableintl_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_enableintl_CEMUXNOT
    );
  tx_input_enableintl_YUSED : X_BUF
    port map (
      I => tx_input_enableintl_GSHIFT,
      O => tx_input_enableint
    );
  mac_control_PHY_status_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"F3F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_done,
      ADR2 => mac_control_PHY_status_cs_FFd3,
      ADR3 => mac_control_PHY_status_cs_FFd2,
      O => mac_control_PHY_status_cs_FFd2_In
    );
  mac_control_PHY_status_cs_FFd1_In1 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => mac_control_PHY_status_done,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_cs_FFd2,
      O => mac_control_PHY_status_cs_FFd1_In
    );
  mac_control_PHY_status_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_cs_FFd5,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_done,
      O => mac_control_PHY_status_cs_FFd4_In
    );
  mac_control_PHY_status_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_cs_FFd4,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_phyaddrws,
      O => mac_control_PHY_status_cs_FFd3_In
    );
  mac_control_PHY_status_cs_FFd6_In1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd7,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_done,
      ADR3 => VCC,
      O => mac_control_PHY_status_cs_FFd6_In
    );
  mac_control_PHY_status_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"F4F4"
    )
    port map (
      ADR0 => mac_control_PHY_status_done,
      ADR1 => mac_control_PHY_status_cs_FFd5,
      ADR2 => mac_control_PHY_status_cs_FFd6,
      ADR3 => VCC,
      O => mac_control_PHY_status_cs_FFd5_In
    );
  mac_control_PHY_status_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"BABA"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd1,
      ADR1 => mac_control_PHY_status_phyaddrws,
      ADR2 => mac_control_PHY_status_cs_FFd4,
      ADR3 => VCC,
      O => mac_control_PHY_status_cs_FFd8_In
    );
  mac_control_PHY_status_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"F2F2"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd7,
      ADR1 => mac_control_PHY_status_done,
      ADR2 => mac_control_PHY_status_cs_FFd8,
      ADR3 => VCC,
      O => mac_control_PHY_status_cs_FFd7_In
    );
  rx_input_memio_n00491 : X_LUT4
    generic map(
      INIT => X"0030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_invalid,
      ADR2 => rx_input_ce,
      ADR3 => rx_input_endf,
      O => rx_input_memio_n0049
    );
  rx_input_memio_crcen_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcen_CEMUXNOT
    );
  tx_input_Mxor_lden_Result1 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_enableint,
      ADR2 => tx_input_enableintl,
      ADR3 => VCC,
      O => tx_input_lden
    );
  tx_input_den_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_den_CEMUXNOT
    );
  tx_output_crcl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_7_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_7_FFY_RST,
      O => tx_output_crcl(7)
    );
  tx_output_crcl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_7_FFY_RST
    );
  tx_input_Mmux_n0032_Result_1_1 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => tx_input_n0074(1),
      ADR1 => tx_input_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_input_dinint(1),
      O => tx_input_n0032(1)
    );
  tx_input_Mmux_n0032_Result_0_1 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => tx_input_n0074(0),
      ADR1 => VCC,
      ADR2 => tx_input_cs_FFd12,
      ADR3 => tx_input_dinint(0),
      O => tx_input_n0032(0)
    );
  tx_input_Mmux_n0032_Result_3_1 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => tx_input_n0074(3),
      ADR1 => tx_input_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_input_dinint(3),
      O => tx_input_n0032(3)
    );
  tx_input_Mmux_n0032_Result_2_1 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_cs_FFd12,
      ADR2 => tx_input_n0074(2),
      ADR3 => tx_input_dinint(2),
      O => tx_input_n0032(2)
    );
  tx_input_Mmux_n0032_Result_5_1 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => tx_input_dinint(5),
      ADR1 => tx_input_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_input_n0074(5),
      O => tx_input_n0032(5)
    );
  tx_input_Mmux_n0032_Result_4_1 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => tx_input_n0074(4),
      ADR1 => tx_input_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_input_dinint(4),
      O => tx_input_n0032(4)
    );
  tx_input_Mmux_n0032_Result_7_1 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_n0074(7),
      ADR2 => tx_input_dinint(7),
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(7)
    );
  tx_input_Mmux_n0032_Result_6_1 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => tx_input_n0074(6),
      ADR1 => VCC,
      ADR2 => tx_input_dinint(6),
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(6)
    );
  tx_input_Mmux_n0032_Result_9_1 : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => tx_input_dinint(9),
      ADR1 => tx_input_n0074(9),
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(9)
    );
  tx_input_Mmux_n0032_Result_8_1 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => tx_input_dinint(8),
      ADR1 => VCC,
      ADR2 => tx_input_n0074(8),
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(8)
    );
  rx_input_GMII_dvdelta1 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_GMII_rx_dvl,
      ADR2 => VCC,
      ADR3 => rx_input_GMII_rx_dvll,
      O => rx_input_endfin_FROM
    );
  rx_input_GMII_endf1 : X_LUT4
    generic map(
      INIT => X"FFF3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_GMII_rx_dvl,
      ADR2 => rx_input_GMII_rx_of,
      ADR3 => rx_input_GMII_rx_erl,
      O => rx_input_endfin_GROM
    );
  rx_input_endfin_XUSED : X_BUF
    port map (
      I => rx_input_endfin_FROM,
      O => rx_input_GMII_dvdelta
    );
  rx_input_endfin_YUSED : X_BUF
    port map (
      I => rx_input_endfin_GROM,
      O => rx_input_GMII_endf
    );
  rx_output_fifo_BU16 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_denll,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_empty,
      O => rx_output_invalid_FROM
    );
  rx_output_fifo_BU29 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => rx_output_denll,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_empty,
      ADR3 => VCC,
      O => rx_output_fifo_N1835
    );
  rx_output_invalid_XUSED : X_BUF
    port map (
      I => rx_output_invalid_FROM,
      O => rx_output_fifo_N1515
    );
  rx_output_fifo_BU90 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N16,
      ADR3 => rx_output_fifo_N17,
      O => rx_output_fifo_N2259
    );
  rx_output_fifo_BU97 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N16,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N15,
      O => rx_output_fifo_N2299
    );
  tx_output_n0034_1_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_1_Q,
      O => tx_output_n0034_1_Q
    );
  tx_output_n0034_0_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16,
      ADR3 => tx_output_crc_0_Q,
      O => tx_output_n0034_0_Q
    );
  mac_control_lsclkdelta1 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => mac_control_sclkl,
      ADR1 => VCC,
      ADR2 => mac_control_sclkll,
      ADR3 => VCC,
      O => mac_control_lsclkdelta
    );
  mac_control_sclkdelta_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_sclkdelta_CEMUXNOT
    );
  rx_input_memio_n0048_1_1 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crc_1_Q,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => VCC,
      O => rx_input_memio_n0048_1_Q
    );
  rx_input_memio_n0048_0_1 : X_LUT4
    generic map(
      INIT => X"FCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crc_0_Q,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => VCC,
      O => rx_input_memio_n0048_0_Q
    );
  tx_output_cs_FFd16_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd16_FFY_RST
    );
  tx_output_cs_FFd16_1_1584 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd16_GROM,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd16_FFY_RST,
      O => tx_output_cs_FFd16_1
    );
  tx_output_cs_FFd16_In1 : X_LUT4
    generic map(
      INIT => X"0200"
    )
    port map (
      ADR0 => tx_output_cs_FFd17,
      ADR1 => memcontroller_clknum_1_1,
      ADR2 => tx_output_n0006,
      ADR3 => memcontroller_clknum_0_1,
      O => tx_output_cs_FFd16_GROM
    );
  tx_output_cs_FFd16_YUSED : X_BUF
    port map (
      I => tx_output_cs_FFd16_GROM,
      O => tx_output_cs_FFd16_In
    );
  mac_control_n00501 : X_LUT4
    generic map(
      INIT => X"8888"
    )
    port map (
      ADR0 => mac_control_N53194,
      ADR1 => mac_control_din(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => mac_control_n0050
    );
  mac_control_rxphyerr_rst_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_rst_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_1_1 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => rx_output_mdl(17),
      ADR1 => rx_output_lmasell,
      ADR2 => VCC,
      ADR3 => rx_output_mdl(1),
      O => rx_output_lma(1)
    );
  rx_output_Mmux_lma_Result_0_1 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => rx_output_mdl(0),
      ADR1 => VCC,
      ADR2 => rx_output_mdl(16),
      ADR3 => rx_output_lmasell,
      O => rx_output_lma(0)
    );
  rx_output_fifodin_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_1_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_3_1 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => rx_output_mdl(3),
      ADR1 => VCC,
      ADR2 => rx_output_lmasell,
      ADR3 => rx_output_mdl(19),
      O => rx_output_lma(3)
    );
  rx_output_Mmux_lma_Result_2_1 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => rx_output_mdl(2),
      ADR1 => rx_output_lmasell,
      ADR2 => rx_output_mdl(18),
      ADR3 => VCC,
      O => rx_output_lma(2)
    );
  rx_output_fifodin_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_3_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_5_1 : X_LUT4
    generic map(
      INIT => X"B8B8"
    )
    port map (
      ADR0 => rx_output_mdl(21),
      ADR1 => rx_output_lmasell,
      ADR2 => rx_output_mdl(5),
      ADR3 => VCC,
      O => rx_output_lma(5)
    );
  rx_output_Mmux_lma_Result_4_1 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_mdl(20),
      ADR2 => rx_output_lmasell,
      ADR3 => rx_output_mdl(4),
      O => rx_output_lma(4)
    );
  rx_output_fifodin_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_5_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_7_1 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => rx_output_mdl(23),
      ADR1 => rx_output_mdl(7),
      ADR2 => rx_output_lmasell,
      ADR3 => VCC,
      O => rx_output_lma(7)
    );
  rx_output_Mmux_lma_Result_6_1 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_mdl(6),
      ADR2 => rx_output_mdl(22),
      ADR3 => rx_output_lmasell,
      O => rx_output_lma(6)
    );
  rx_output_fifodin_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_7_CEMUXNOT
    );
  rx_output_Mmux_lma_Result_9_1 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_lmasell,
      ADR2 => rx_output_mdl(9),
      ADR3 => rx_output_mdl(25),
      O => rx_output_lma(9)
    );
  rx_output_Mmux_lma_Result_8_1 : X_LUT4
    generic map(
      INIT => X"B8B8"
    )
    port map (
      ADR0 => rx_output_mdl(24),
      ADR1 => rx_output_lmasell,
      ADR2 => rx_output_mdl(8),
      ADR3 => VCC,
      O => rx_output_lma(8)
    );
  rx_output_fifodin_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifodin_9_CEMUXNOT
    );
  rx_output_n00511 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rx_output_fifo_wrcount(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_wrcount(0),
      O => rx_output_n0051
    );
  rx_output_fifo_full_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_fifo_full_CEMUXNOT
    );
  rx_input_GMII_lfifoin_0_11 : X_LUT4
    generic map(
      INIT => X"00C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_GMII_rx_dvl,
      ADR2 => rx_input_GMII_rxdl(0),
      ADR3 => rx_input_GMII_rx_of,
      O => rx_input_GMII_N79913
    );
  rx_input_GMII_lfifoin_1_11 : X_LUT4
    generic map(
      INIT => X"2020"
    )
    port map (
      ADR0 => rx_input_GMII_rxdl(1),
      ADR1 => rx_input_GMII_rx_erl,
      ADR2 => rx_input_GMII_rx_dvl,
      ADR3 => VCC,
      O => rx_input_GMII_N79916
    );
  rx_input_GMII_lfifoin_3_11 : X_LUT4
    generic map(
      INIT => X"0808"
    )
    port map (
      ADR0 => rx_input_GMII_rxdl(3),
      ADR1 => rx_input_GMII_rx_dvl,
      ADR2 => rx_input_GMII_rx_erl,
      ADR3 => VCC,
      O => rx_input_GMII_N79922
    );
  rx_input_GMII_lfifoin_2_11 : X_LUT4
    generic map(
      INIT => X"FAAA"
    )
    port map (
      ADR0 => rx_input_GMII_rx_erl,
      ADR1 => VCC,
      ADR2 => rx_input_GMII_rx_dvl,
      ADR3 => rx_input_GMII_rxdl(2),
      O => rx_input_GMII_N79919
    );
  rx_input_GMII_lfifoin_5_11 : X_LUT4
    generic map(
      INIT => X"0808"
    )
    port map (
      ADR0 => rx_input_GMII_rx_dvl,
      ADR1 => rx_input_GMII_rxdl(5),
      ADR2 => rx_input_GMII_rx_erl,
      ADR3 => VCC,
      O => rx_input_GMII_N79901
    );
  rx_input_GMII_lfifoin_4_11 : X_LUT4
    generic map(
      INIT => X"4400"
    )
    port map (
      ADR0 => rx_input_GMII_rx_erl,
      ADR1 => rx_input_GMII_rxdl(4),
      ADR2 => VCC,
      ADR3 => rx_input_GMII_rx_dvl,
      O => rx_input_GMII_N79910
    );
  rx_input_GMII_lfifoin_7_11 : X_LUT4
    generic map(
      INIT => X"2020"
    )
    port map (
      ADR0 => rx_input_GMII_rx_dvl,
      ADR1 => rx_input_GMII_rx_erl,
      ADR2 => rx_input_GMII_rxdl(7),
      ADR3 => VCC,
      O => rx_input_GMII_N79907
    );
  rx_input_GMII_lfifoin_6_11 : X_LUT4
    generic map(
      INIT => X"2200"
    )
    port map (
      ADR0 => rx_input_GMII_rx_dvl,
      ADR1 => rx_input_GMII_rx_erl,
      ADR2 => VCC,
      ADR3 => rx_input_GMII_rxdl(6),
      O => rx_input_GMII_N79904
    );
  tx_input_dinint_11_LOGIC_ONE_1585 : X_ONE
    port map (
      O => tx_input_dinint_11_LOGIC_ONE
    );
  tx_input_srl16_din_bit11_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_30,
      A1 => GLOBAL_LOGIC0_30,
      A2 => GLOBAL_LOGIC1_22,
      A3 => GLOBAL_LOGIC0_35,
      D => tx_input_dinl(11),
      CE => tx_input_dinint_11_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(11)
    );
  tx_input_srl16_din_bit10_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_30,
      A1 => GLOBAL_LOGIC0_30,
      A2 => GLOBAL_LOGIC1_22,
      A3 => GLOBAL_LOGIC0_35,
      D => tx_input_dinl(10),
      CE => tx_input_dinint_11_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(10)
    );
  tx_input_dinint_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_11_CEMUXNOT
    );
  tx_input_dinint_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_13_FFY_RST
    );
  tx_input_dinint_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(12),
      CE => tx_input_dinint_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_13_FFY_RST,
      O => tx_input_dinint(12)
    );
  tx_input_dinint_13_LOGIC_ONE_1586 : X_ONE
    port map (
      O => tx_input_dinint_13_LOGIC_ONE
    );
  tx_input_srl16_din_bit13_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_35,
      A1 => GLOBAL_LOGIC0_35,
      A2 => GLOBAL_LOGIC1_20,
      A3 => GLOBAL_LOGIC0_29,
      D => tx_input_dinl(13),
      CE => tx_input_dinint_13_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(13)
    );
  tx_input_srl16_din_bit12_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_35,
      A1 => GLOBAL_LOGIC0_35,
      A2 => GLOBAL_LOGIC1_20,
      A3 => GLOBAL_LOGIC0_29,
      D => tx_input_dinl(12),
      CE => tx_input_dinint_13_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(12)
    );
  tx_input_dinint_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_13_CEMUXNOT
    );
  tx_input_dinint_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_15_FFY_RST
    );
  tx_input_dinint_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(14),
      CE => tx_input_dinint_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_15_FFY_RST,
      O => tx_input_dinint(14)
    );
  tx_input_dinint_15_LOGIC_ONE_1587 : X_ONE
    port map (
      O => tx_input_dinint_15_LOGIC_ONE
    );
  tx_input_srl16_din_bit15_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_38,
      A1 => GLOBAL_LOGIC0_38,
      A2 => GLOBAL_LOGIC1_21,
      A3 => GLOBAL_LOGIC0_34,
      D => tx_input_dinl(15),
      CE => tx_input_dinint_15_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(15)
    );
  tx_input_srl16_din_bit14_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_38,
      A1 => GLOBAL_LOGIC0_38,
      A2 => GLOBAL_LOGIC1_21,
      A3 => GLOBAL_LOGIC0_34,
      D => tx_input_dinl(14),
      CE => tx_input_dinint_15_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(14)
    );
  tx_input_dinint_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_15_CEMUXNOT
    );
  memcontroller_oe_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_oe_FFY_RST
    );
  memcontroller_oe_1588 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_wen,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_oe_FFY_RST,
      O => memcontroller_oe
    );
  memcontroller_n00111 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => memcontroller_clknum_0_1,
      ADR1 => VCC,
      ADR2 => memcontroller_clknum_1_2,
      ADR3 => VCC,
      O => memcontroller_wen
    );
  rx_input_memio_n00611 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => rxfifofull,
      ADR1 => rx_input_memio_cs_FFd5,
      ADR2 => rx_input_memio_endbyte(2),
      ADR3 => rx_input_memio_crcequal,
      O => rx_input_memio_n0061
    );
  rx_input_memio_n00601 : X_LUT4
    generic map(
      INIT => X"1010"
    )
    port map (
      ADR0 => rx_input_memio_endbyte(2),
      ADR1 => rx_input_memio_crcequal,
      ADR2 => rx_input_memio_cs_FFd5,
      ADR3 => VCC,
      O => rx_input_memio_n0060
    );
  rxfifowerr_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxfifowerr_CEMUXNOT
    );
  rx_output_cs_FFd17_In1 : X_LUT4
    generic map(
      INIT => X"0008"
    )
    port map (
      ADR0 => rx_output_cs_FFd18,
      ADR1 => memcontroller_clknum(1),
      ADR2 => memcontroller_clknum(0),
      ADR3 => rx_output_n0017,
      O => rx_output_cs_FFd17_In
    );
  rx_output_cs_FFd4_In1 : X_LUT4
    generic map(
      INIT => X"CC80"
    )
    port map (
      ADR0 => rx_output_n0018,
      ADR1 => rx_output_nf,
      ADR2 => rx_output_cs_FFd5,
      ADR3 => rx_output_cs_FFd4,
      O => rx_output_cs_FFd4_In
    );
  rx_output_cs_FFd19_In1 : X_LUT4
    generic map(
      INIT => X"FCDC"
    )
    port map (
      ADR0 => rx_output_nf,
      ADR1 => rx_output_cs_FFd10,
      ADR2 => rx_output_cs_FFd19,
      ADR3 => rx_output_nfl,
      O => rx_output_cs_FFd19_In
    );
  mac_control_dout_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(1),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_1_FFY_RST,
      O => mac_control_dout(1)
    );
  mac_control_dout_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_1_FFY_RST
    );
  rx_input_memio_n00581 : X_LUT4
    generic map(
      INIT => X"2000"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd5,
      ADR1 => rx_input_memio_endbyte(0),
      ADR2 => rx_input_memio_endbyte(2),
      ADR3 => rx_input_memio_endbyte(1),
      O => rx_input_memio_n0058
    );
  rx_input_memio_n00571 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => rx_input_memio_endbyte(1),
      ADR1 => rx_input_memio_endbyte(0),
      ADR2 => rx_input_memio_endbyte(2),
      ADR3 => rx_input_memio_cs_FFd5,
      O => rx_input_memio_n0057
    );
  rxoferr_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxoferr_CEMUXNOT
    );
  tx_input_cs_FFd10_In_SW0 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_den,
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd10,
      O => tx_input_cs_FFd11_FROM
    );
  tx_input_cs_FFd11_In1 : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_den,
      ADR2 => tx_input_cs_FFd12,
      ADR3 => tx_input_newfint,
      O => tx_input_cs_FFd11_In
    );
  tx_input_cs_FFd11_XUSED : X_BUF
    port map (
      I => tx_input_cs_FFd11_FROM,
      O => tx_input_N70883
    );
  tx_output_TXF1 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_ltxen3,
      ADR2 => VCC,
      ADR3 => tx_output_ltxen2,
      O => mac_control_txf_cross_GROM
    );
  mac_control_txf_cross_YUSED : X_BUF
    port map (
      I => mac_control_txf_cross_GROM,
      O => txf
    );
  tx_input_Mmux_n0032_Result_11_1 : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => tx_input_dinint(11),
      ADR1 => tx_input_n0074(11),
      ADR2 => VCC,
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(11)
    );
  tx_input_Mmux_n0032_Result_10_1 : X_LUT4
    generic map(
      INIT => X"F0AA"
    )
    port map (
      ADR0 => tx_input_n0074(10),
      ADR1 => VCC,
      ADR2 => tx_input_dinint(10),
      ADR3 => tx_input_cs_FFd12,
      O => tx_input_n0032(10)
    );
  tx_input_Mmux_n0032_Result_13_1 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => tx_input_n0074(13),
      ADR1 => tx_input_cs_FFd12,
      ADR2 => VCC,
      ADR3 => tx_input_dinint(13),
      O => tx_input_n0032(13)
    );
  tx_input_Mmux_n0032_Result_12_1 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => tx_input_cs_FFd12,
      ADR1 => tx_input_n0074(12),
      ADR2 => tx_input_dinint(12),
      ADR3 => VCC,
      O => tx_input_n0032(12)
    );
  tx_input_Mmux_n0032_Result_15_1 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => tx_input_n0074(15),
      ADR1 => tx_input_cs_FFd12,
      ADR2 => tx_input_dinint(15),
      ADR3 => VCC,
      O => tx_input_n0032(15)
    );
  tx_input_Mmux_n0032_Result_14_1 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_dinint(14),
      ADR2 => tx_input_cs_FFd12,
      ADR3 => tx_input_n0074(14),
      O => tx_input_n0032(14)
    );
  tx_output_cs_FFd5_In1 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_n0007,
      ADR3 => tx_output_cs_FFd6_1,
      O => tx_output_cs_FFd5_GROM
    );
  tx_output_cs_FFd5_YUSED : X_BUF
    port map (
      I => tx_output_cs_FFd5_GROM,
      O => tx_output_cs_FFd5_In
    );
  tx_output_cs_FFd6_In1 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd8,
      ADR3 => tx_output_n0007,
      O => tx_output_cs_FFd6_GROM
    );
  tx_output_cs_FFd6_YUSED : X_BUF
    port map (
      I => tx_output_cs_FFd6_GROM,
      O => tx_output_cs_FFd6_In
    );
  tx_input_dinint_1_LOGIC_ONE_1589 : X_ONE
    port map (
      O => tx_input_dinint_1_LOGIC_ONE
    );
  tx_input_srl16_din_bit1_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_27,
      A1 => GLOBAL_LOGIC0_26,
      A2 => GLOBAL_LOGIC1_18,
      A3 => GLOBAL_LOGIC0_26,
      D => tx_input_dinl(1),
      CE => tx_input_dinint_1_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(1)
    );
  tx_input_srl16_din_bit0_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_27,
      A1 => GLOBAL_LOGIC0_26,
      A2 => GLOBAL_LOGIC1_18,
      A3 => GLOBAL_LOGIC0_26,
      D => tx_input_dinl(0),
      CE => tx_input_dinint_1_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(0)
    );
  tx_input_dinint_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_1_CEMUXNOT
    );
  tx_input_dinint_3_LOGIC_ONE_1590 : X_ONE
    port map (
      O => tx_input_dinint_3_LOGIC_ONE
    );
  tx_input_srl16_din_bit3_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_33,
      A1 => GLOBAL_LOGIC0_33,
      A2 => GLOBAL_LOGIC1_25,
      A3 => GLOBAL_LOGIC0_39,
      D => tx_input_dinl(3),
      CE => tx_input_dinint_3_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(3)
    );
  tx_input_srl16_din_bit2_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_33,
      A1 => GLOBAL_LOGIC0_33,
      A2 => GLOBAL_LOGIC1_25,
      A3 => GLOBAL_LOGIC0_39,
      D => tx_input_dinl(2),
      CE => tx_input_dinint_3_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(2)
    );
  tx_input_dinint_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_3_CEMUXNOT
    );
  tx_input_dinint_5_LOGIC_ONE_1591 : X_ONE
    port map (
      O => tx_input_dinint_5_LOGIC_ONE
    );
  tx_input_srl16_din_bit5_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_32,
      A1 => GLOBAL_LOGIC0_32,
      A2 => GLOBAL_LOGIC1_23,
      A3 => GLOBAL_LOGIC0_36,
      D => tx_input_dinl(5),
      CE => tx_input_dinint_5_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(5)
    );
  tx_input_srl16_din_bit4_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_32,
      A1 => GLOBAL_LOGIC0_32,
      A2 => GLOBAL_LOGIC1_23,
      A3 => GLOBAL_LOGIC0_36,
      D => tx_input_dinl(4),
      CE => tx_input_dinint_5_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(4)
    );
  tx_input_dinint_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_5_CEMUXNOT
    );
  tx_input_dinint_7_LOGIC_ONE_1592 : X_ONE
    port map (
      O => tx_input_dinint_7_LOGIC_ONE
    );
  tx_input_srl16_din_bit7_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_36,
      A1 => GLOBAL_LOGIC0_32,
      A2 => GLOBAL_LOGIC1_23,
      A3 => GLOBAL_LOGIC0_32,
      D => tx_input_dinl(7),
      CE => tx_input_dinint_7_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(7)
    );
  tx_input_srl16_din_bit6_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_36,
      A1 => GLOBAL_LOGIC0_32,
      A2 => GLOBAL_LOGIC1_23,
      A3 => GLOBAL_LOGIC0_32,
      D => tx_input_dinl(6),
      CE => tx_input_dinint_7_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(6)
    );
  tx_input_dinint_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_7_CEMUXNOT
    );
  tx_input_dinint_9_LOGIC_ONE_1593 : X_ONE
    port map (
      O => tx_input_dinint_9_LOGIC_ONE
    );
  tx_input_srl16_din_bit9_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_31,
      A1 => GLOBAL_LOGIC0_31,
      A2 => GLOBAL_LOGIC1_22,
      A3 => GLOBAL_LOGIC0_35,
      D => tx_input_dinl(9),
      CE => tx_input_dinint_9_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(9)
    );
  tx_input_srl16_din_bit8_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_31,
      A1 => GLOBAL_LOGIC0_31,
      A2 => GLOBAL_LOGIC1_22,
      A3 => GLOBAL_LOGIC0_35,
      D => tx_input_dinl(8),
      CE => tx_input_dinint_9_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_ldinint(8)
    );
  tx_input_dinint_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_dinint_9_CEMUXNOT
    );
  rx_input_fifo_control_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_ce,
      ADR3 => rx_input_fifo_control_cs_FFd3,
      O => rx_input_fifo_control_cs_FFd2_In
    );
  rx_input_fifo_control_cs_FFd1_In1 : X_LUT4
    generic map(
      INIT => X"CCC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_ce,
      ADR2 => rx_input_fifo_control_cs_FFd1,
      ADR3 => rx_input_fifo_control_cs_FFd2,
      O => rx_input_fifo_control_cs_FFd1_In
    );
  mac_control_PHY_status_din_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(2),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_3_FFY_RST,
      O => mac_control_PHY_status_din(2)
    );
  mac_control_PHY_status_din_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_3_FFY_RST
    );
  rx_output_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"AA00"
    )
    port map (
      ADR0 => rx_output_cs_FFd3,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_nf,
      O => rx_output_cs_FFd2_In
    );
  rx_output_cs_FFd1_In1 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_cs_FFd2,
      ADR3 => rx_output_nf,
      O => rx_output_cs_FFd1_In
    );
  rx_output_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_cs_FFd9,
      ADR2 => VCC,
      ADR3 => rx_output_nf,
      O => rx_output_cs_FFd8_In
    );
  rx_output_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_nf,
      ADR2 => rx_output_cs_FFd8,
      ADR3 => VCC,
      O => rx_output_cs_FFd7_In
    );
  rx_input_GMII_lince1 : X_LUT4
    generic map(
      INIT => X"CCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_GMII_ro,
      ADR2 => rx_input_GMII_rx_dvl,
      ADR3 => rx_input_GMII_rx_dvll,
      O => rx_input_GMII_lince
    );
  tx_input_cs_FFd2_In1 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_input_fifofulll,
      ADR3 => tx_input_cs_FFd5,
      O => tx_input_cs_FFd2_In
    );
  tx_input_cs_FFd3_In1 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_input_cs_FFd5,
      ADR3 => tx_input_fifofulll,
      O => tx_input_cs_FFd3_In
    );
  tx_input_cs_FFd10_In : X_LUT4
    generic map(
      INIT => X"FFF2"
    )
    port map (
      ADR0 => tx_input_cs_FFd6,
      ADR1 => tx_input_N35861,
      ADR2 => tx_input_cs_FFd11,
      ADR3 => tx_input_N70883,
      O => tx_input_cs_FFd10_In_O
    );
  tx_input_cs_FFd9_In1 : X_LUT4
    generic map(
      INIT => X"C0C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_input_den,
      ADR2 => tx_input_cs_FFd10,
      ADR3 => VCC,
      O => tx_input_cs_FFd9_In
    );
  mac_control_PHY_status_din_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(1),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_1_FFX_RST,
      O => mac_control_PHY_status_din(1)
    );
  mac_control_PHY_status_din_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_1_FFX_RST
    );
  rx_input_memio_Mshreg_lbpout4_10_srl_5 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_2,
      A1 => GLOBAL_LOGIC1_0,
      A2 => GLOBAL_LOGIC0_2,
      A3 => GLOBAL_LOGIC0_2,
      D => rx_input_memio_bp(10),
      CE => rx_input_memio_Mshreg_lbpout4_10_59_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_10_net14
    );
  rx_input_memio_Mshreg_lbpout4_10_59_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_10_59_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_10_59_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_10_59_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_11_srl_4 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_4,
      A1 => GLOBAL_LOGIC1_5,
      A2 => GLOBAL_LOGIC0_5,
      A3 => GLOBAL_LOGIC0_4,
      D => rx_input_memio_bp(11),
      CE => rx_input_memio_Mshreg_lbpout4_11_58_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_11_net12
    );
  rx_input_memio_Mshreg_lbpout4_11_58_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_11_58_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_11_58_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_11_58_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_12_srl_3 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_10,
      A1 => GLOBAL_LOGIC1_1,
      A2 => GLOBAL_LOGIC0_10,
      A3 => GLOBAL_LOGIC0_10,
      D => rx_input_memio_bp(12),
      CE => rx_input_memio_Mshreg_lbpout4_12_57_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_12_net10
    );
  rx_input_memio_Mshreg_lbpout4_12_57_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_12_57_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_12_57_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_12_57_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_13_srl_2 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_12,
      A1 => GLOBAL_LOGIC1_3,
      A2 => GLOBAL_LOGIC0_12,
      A3 => GLOBAL_LOGIC0_12,
      D => rx_input_memio_bp(13),
      CE => rx_input_memio_Mshreg_lbpout4_13_56_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_13_net8
    );
  rx_input_memio_Mshreg_lbpout4_13_56_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_13_56_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_13_56_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_13_56_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_14_srl_1 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_12,
      A1 => GLOBAL_LOGIC1_3,
      A2 => GLOBAL_LOGIC0_12,
      A3 => GLOBAL_LOGIC0_12,
      D => rx_input_memio_bp(14),
      CE => rx_input_memio_Mshreg_lbpout4_14_55_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_14_net6
    );
  rx_input_memio_Mshreg_lbpout4_14_55_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_14_55_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_14_55_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_14_55_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_15_srl_0 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_9,
      A1 => GLOBAL_LOGIC1_0,
      A2 => GLOBAL_LOGIC0_9,
      A3 => GLOBAL_LOGIC0_9,
      D => rx_input_memio_bp(15),
      CE => rx_input_memio_Mshreg_lbpout4_15_54_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_15_net4
    );
  rx_input_memio_Mshreg_lbpout4_15_54_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_15_54_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_15_54_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_15_54_SRMUX_OUTPUTNOT
    );
  mac_control_Mshreg_sinlll_srl_16 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC1_26,
      A1 => GLOBAL_LOGIC0_41,
      A2 => GLOBAL_LOGIC0_41,
      A3 => GLOBAL_LOGIC0_41,
      D => SIN_IBUF,
      CE => mac_control_Mshreg_sinlll_102_SRMUX_OUTPUTNOT,
      CLK => mac_control_CLKSL_4,
      Q => mac_control_Mshreg_sinlll_net185
    );
  mac_control_Mshreg_sinlll_102_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_Mshreg_sinlll_102_CEMUXNOT
    );
  mac_control_Mshreg_sinlll_102_SRMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_Mshreg_sinlll_102_SRMUX_OUTPUTNOT
    );
  rx_output_fifo_BU104 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N15,
      ADR2 => rx_output_fifo_N14,
      ADR3 => VCC,
      O => rx_output_fifo_N2339
    );
  rx_output_fifo_BU111 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N14,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N13,
      O => rx_output_fifo_N2379
    );
  rx_output_fifo_BU118 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N12,
      ADR2 => rx_output_fifo_N13,
      ADR3 => VCC,
      O => rx_output_fifo_N2419
    );
  rx_output_fifo_BU125 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_fifo_N11,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N12,
      O => rx_output_fifo_N2459
    );
  rx_output_fifo_BU265 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_output_fifo_N6,
      ADR3 => rx_output_fifo_N7,
      O => rx_output_fifo_N3267
    );
  rx_output_fifo_BU272 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N5,
      ADR2 => rx_output_fifo_N6,
      ADR3 => VCC,
      O => rx_output_fifo_N3307
    );
  mac_control_PHY_status_din_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(3),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_3_FFX_RST,
      O => mac_control_PHY_status_din(3)
    );
  mac_control_PHY_status_din_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_3_FFX_RST
    );
  rx_output_fifo_BU251 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_fifo_N8,
      ADR1 => rx_output_fifo_N9,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N3187
    );
  rx_output_fifo_BU258 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N8,
      ADR2 => rx_output_fifo_N7,
      ADR3 => VCC,
      O => rx_output_fifo_N3227
    );
  rx_output_fifo_BU279 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_fifo_N4,
      ADR1 => rx_output_fifo_N5,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N3347
    );
  rx_output_fifo_BU286 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rx_output_fifo_N3,
      ADR1 => rx_output_fifo_N4,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_output_fifo_N3387
    );
  rx_output_fifo_BU422 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_output_fifo_N1579,
      ADR1 => rx_output_fifo_N1581,
      ADR2 => rx_output_fifo_N1580,
      ADR3 => rx_output_fifo_N1578,
      O => rx_output_fifo_N1589_FROM
    );
  rx_output_fifo_BU428 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rx_output_fifo_N1582,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N3959,
      O => rx_output_fifo_N3971
    );
  rx_output_fifo_N1589_XUSED : X_BUF
    port map (
      I => rx_output_fifo_N1589_FROM,
      O => rx_output_fifo_N3959
    );
  rx_output_fifo_BU416 : X_LUT4
    generic map(
      INIT => X"C33C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N1579,
      ADR2 => rx_output_fifo_N1578,
      ADR3 => rx_output_fifo_N1580,
      O => rx_output_fifo_N3973
    );
  rx_output_fifo_BU452 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_fifo_N3958,
      ADR2 => VCC,
      ADR3 => rx_output_fifo_N3959,
      O => rx_output_fifo_N3968
    );
  rx_output_fifo_BU440 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_output_fifo_N1583,
      ADR1 => rx_output_fifo_N1582,
      ADR2 => rx_output_fifo_N1584,
      ADR3 => rx_output_fifo_N3959,
      O => rx_output_fifo_N3969
    );
  tx_output_cs_FFd8_In1 : X_LUT4
    generic map(
      INIT => X"CFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd9,
      ADR2 => tx_output_n0007,
      ADR3 => tx_output_cs_FFd4_1,
      O => tx_output_cs_FFd8_In
    );
  tx_output_cs_FFd7_In1 : X_LUT4
    generic map(
      INIT => X"A0A0"
    )
    port map (
      ADR0 => tx_output_decbcnt,
      ADR1 => VCC,
      ADR2 => tx_output_n0007,
      ADR3 => VCC,
      O => tx_output_cs_FFd7_In
    );
  rx_input_memio_Mshreg_lbpout4_0_srl_15 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_4,
      A1 => GLOBAL_LOGIC1_5,
      A2 => GLOBAL_LOGIC0_5,
      A3 => GLOBAL_LOGIC0_4,
      D => rx_input_memio_bp(0),
      CE => rx_input_memio_Mshreg_lbpout4_0_69_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_0_net34
    );
  rx_input_memio_Mshreg_lbpout4_0_69_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_0_69_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_0_69_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_0_69_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_1_srl_14 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_5,
      A1 => GLOBAL_LOGIC1_33,
      A2 => GLOBAL_LOGIC0_5,
      A3 => GLOBAL_LOGIC0_6,
      D => rx_input_memio_bp(1),
      CE => rx_input_memio_Mshreg_lbpout4_1_68_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_1_net32
    );
  rx_input_memio_Mshreg_lbpout4_1_68_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_1_68_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_1_68_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_1_68_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_2_srl_13 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0,
      A1 => GLOBAL_LOGIC1,
      A2 => GLOBAL_LOGIC0_8,
      A3 => GLOBAL_LOGIC0_8,
      D => rx_input_memio_bp(2),
      CE => rx_input_memio_Mshreg_lbpout4_2_67_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_2_net30
    );
  rx_input_memio_Mshreg_lbpout4_2_67_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_2_67_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_2_67_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_2_67_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_3_srl_12 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_8,
      A1 => GLOBAL_LOGIC1,
      A2 => GLOBAL_LOGIC0_8,
      A3 => GLOBAL_LOGIC0_8,
      D => rx_input_memio_bp(3),
      CE => rx_input_memio_Mshreg_lbpout4_3_66_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_3_net28
    );
  rx_input_memio_Mshreg_lbpout4_3_66_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_3_66_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_3_66_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_3_66_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_4_srl_11 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_5,
      A1 => GLOBAL_LOGIC1_5,
      A2 => GLOBAL_LOGIC0_5,
      A3 => GLOBAL_LOGIC0_5,
      D => rx_input_memio_bp(4),
      CE => rx_input_memio_Mshreg_lbpout4_4_65_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_4_net26
    );
  rx_input_memio_Mshreg_lbpout4_4_65_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_4_65_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_4_65_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_4_65_SRMUX_OUTPUTNOT
    );
  mac_control_PHY_status_din_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(5),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_5_FFX_RST,
      O => mac_control_PHY_status_din(5)
    );
  mac_control_PHY_status_din_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_5_FFX_RST
    );
  rx_input_memio_Mshreg_lbpout4_5_srl_10 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_5,
      A1 => GLOBAL_LOGIC1_5,
      A2 => GLOBAL_LOGIC0_13,
      A3 => GLOBAL_LOGIC0_5,
      D => rx_input_memio_bp(5),
      CE => rx_input_memio_Mshreg_lbpout4_5_64_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_5_net24
    );
  rx_input_memio_Mshreg_lbpout4_5_64_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_5_64_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_5_64_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_5_64_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_6_srl_9 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_13,
      A1 => GLOBAL_LOGIC1_4,
      A2 => GLOBAL_LOGIC0_13,
      A3 => GLOBAL_LOGIC0_13,
      D => rx_input_memio_bp(6),
      CE => rx_input_memio_Mshreg_lbpout4_6_63_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_6_net22
    );
  rx_input_memio_Mshreg_lbpout4_6_63_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_6_63_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_6_63_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_6_63_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_7_srl_8 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_13,
      A1 => GLOBAL_LOGIC1_4,
      A2 => GLOBAL_LOGIC0_13,
      A3 => GLOBAL_LOGIC0_13,
      D => rx_input_memio_bp(7),
      CE => rx_input_memio_Mshreg_lbpout4_7_62_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_7_net20
    );
  rx_input_memio_Mshreg_lbpout4_7_62_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_7_62_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_7_62_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_7_62_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_8_srl_7 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_8,
      A1 => GLOBAL_LOGIC1,
      A2 => GLOBAL_LOGIC0_8,
      A3 => GLOBAL_LOGIC0_8,
      D => rx_input_memio_bp(8),
      CE => rx_input_memio_Mshreg_lbpout4_8_61_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_8_net18
    );
  rx_input_memio_Mshreg_lbpout4_8_61_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_8_61_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_8_61_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_8_61_SRMUX_OUTPUTNOT
    );
  rx_input_memio_Mshreg_lbpout4_9_srl_6 : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_9,
      A1 => GLOBAL_LOGIC1_1,
      A2 => GLOBAL_LOGIC0_9,
      A3 => GLOBAL_LOGIC0_9,
      D => rx_input_memio_bp(9),
      CE => rx_input_memio_Mshreg_lbpout4_9_60_SRMUX_OUTPUTNOT,
      CLK => GTX_CLK_OBUF,
      Q => rx_input_memio_Mshreg_lbpout4_9_net16
    );
  rx_input_memio_Mshreg_lbpout4_9_60_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_9_60_CEMUXNOT
    );
  rx_input_memio_Mshreg_lbpout4_9_60_SRMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_Mshreg_lbpout4_9_60_SRMUX_OUTPUTNOT
    );
  tx_input_newfint_LOGIC_ONE_1594 : X_ONE
    port map (
      O => tx_input_newfint_LOGIC_ONE
    );
  tx_input_srl16_newframe_SRL16E : X_SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => GLOBAL_LOGIC0_26,
      A1 => GLOBAL_LOGIC0_26,
      A2 => GLOBAL_LOGIC1_18,
      A3 => GLOBAL_LOGIC0_27,
      D => tx_input_newframel,
      CE => tx_input_newfint_LOGIC_ONE,
      CLK => GTX_CLK_OBUF,
      Q => tx_input_lnewfint
    );
  tx_input_newfint_CEMUX : X_INV
    port map (
      I => RESET_IBUF_1,
      O => tx_input_newfint_CEMUXNOT
    );
  tx_output_n0034_21_1 : X_LUT4
    generic map(
      INIT => X"F9F6"
    )
    port map (
      ADR0 => tx_output_data(2),
      ADR1 => tx_output_crcl(29),
      ADR2 => tx_output_cs_FFd16_1,
      ADR3 => tx_output_crcl(13),
      O => tx_output_n0034_21_Q
    );
  tx_output_n0034_20_1 : X_LUT4
    generic map(
      INIT => X"EBBE"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => tx_output_crcl(28),
      ADR2 => tx_output_data(3),
      ADR3 => tx_output_crcl(12),
      O => tx_output_n0034_20_Q
    );
  mac_control_PHY_status_din_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(8),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_9_FFY_RST,
      O => mac_control_PHY_status_din(8)
    );
  mac_control_PHY_status_din_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_9_FFY_RST
    );
  tx_output_crc_loigc_Mxor_CO_23_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(25),
      ADR1 => tx_output_data(7),
      ADR2 => tx_output_crcl(24),
      ADR3 => tx_output_data(6),
      O => tx_output_crcl_22_FROM
    );
  tx_output_n0034_22_1 : X_LUT4
    generic map(
      INIT => X"F9F6"
    )
    port map (
      ADR0 => tx_output_crcl(14),
      ADR1 => tx_output_data(7),
      ADR2 => tx_output_cs_FFd16_1,
      ADR3 => tx_output_crcl(24),
      O => tx_output_n0034_22_Q
    );
  tx_output_crcl_22_XUSED : X_BUF
    port map (
      I => tx_output_crcl_22_FROM,
      O => tx_output_crc_loigc_Mxor_CO_23_Xo(0)
    );
  tx_output_crc_loigc_Mxor_n0007_Xo_0_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(2),
      ADR1 => tx_output_crcl(29),
      ADR2 => tx_output_crcl(25),
      ADR3 => tx_output_data(6),
      O => tx_output_crcl_31_FROM
    );
  tx_output_n0034_31_1 : X_LUT4
    generic map(
      INIT => X"EDDE"
    )
    port map (
      ADR0 => tx_output_data(2),
      ADR1 => tx_output_cs_FFd16_1,
      ADR2 => tx_output_crcl(23),
      ADR3 => tx_output_crcl(29),
      O => tx_output_n0034_31_Q
    );
  tx_output_crcl_31_XUSED : X_BUF
    port map (
      I => tx_output_crcl_31_FROM,
      O => tx_output_crc_loigc_Mxor_n0007_Xo(0)
    );
  mac_control_PHY_status_din_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(7),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_7_FFX_RST,
      O => mac_control_PHY_status_din(7)
    );
  mac_control_PHY_status_din_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_7_FFX_RST
    );
  tx_output_crc_loigc_Mxor_CO_13_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(4),
      ADR1 => tx_output_data(0),
      ADR2 => tx_output_crcl(27),
      ADR3 => tx_output_crcl(31),
      O => tx_output_crcl_19_FROM
    );
  tx_output_n0034_19_1 : X_LUT4
    generic map(
      INIT => X"F5FA"
    )
    port map (
      ADR0 => tx_output_crcl(11),
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16_1,
      ADR3 => tx_output_crc_loigc_Mxor_CO_13_Xo(2),
      O => tx_output_n0034_19_Q
    );
  tx_output_crcl_19_XUSED : X_BUF
    port map (
      I => tx_output_crcl_19_FROM,
      O => tx_output_crc_loigc_Mxor_CO_13_Xo(2)
    );
  tx_output_crc_loigc_Mxor_CO_13_Xo_5_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_Mxor_CO_18_Xo(0),
      ADR1 => tx_output_crc_loigc_Mxor_n0007_Xo(0),
      ADR2 => tx_output_crcl(5),
      ADR3 => tx_output_crc_loigc_Mxor_CO_13_Xo(2),
      O => tx_output_crcl_13_FROM
    );
  tx_output_n0034_13_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16_1,
      ADR3 => tx_output_crc_13_Q,
      O => tx_output_n0034_13_Q
    );
  tx_output_crcl_13_XUSED : X_BUF
    port map (
      I => tx_output_crcl_13_FROM,
      O => tx_output_crc_13_Q
    );
  rx_input_memio_crccomb_Mxor_CO_6_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_Mxor_CO_18_Xo(0),
      ADR1 => rx_input_memio_crccomb_n0124(0),
      ADR2 => rx_input_memio_crccomb_Mxor_n0007_Xo(0),
      ADR3 => rx_input_memio_crccomb_n0115(0),
      O => rx_input_memio_crcl_6_FROM
    );
  rx_input_memio_n0048_6_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_6_Q,
      O => rx_input_memio_n0048_6_1_O
    );
  rx_input_memio_crcl_6_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_6_FROM,
      O => rx_input_memio_crc_6_Q
    );
  tx_output_crcsell_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_crcsell_3_CEMUXNOT
    );
  memcontroller_dnl2_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_1_CEMUXNOT
    );
  mac_control_PHY_status_din_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(9),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_9_FFX_RST,
      O => mac_control_PHY_status_din(9)
    );
  mac_control_PHY_status_din_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_9_FFX_RST
    );
  memcontroller_dnl2_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_3_CEMUXNOT
    );
  tx_output_crc_loigc_Mxor_CO_30_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_data(0),
      ADR1 => tx_output_crcl(22),
      ADR2 => tx_output_crcl(31),
      ADR3 => tx_output_crc_loigc_n0115(0),
      O => tx_output_crcl_30_FROM
    );
  tx_output_n0034_30_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16_1,
      ADR2 => VCC,
      ADR3 => tx_output_crc_30_Q,
      O => tx_output_n0034_30_1_O
    );
  tx_output_crcl_30_XUSED : X_BUF
    port map (
      I => tx_output_crcl_30_FROM,
      O => tx_output_crc_30_Q
    );
  memcontroller_dnl2_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_5_CEMUXNOT
    );
  memcontroller_dnl2_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_7_CEMUXNOT
    );
  memcontroller_dnl2_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_9_CEMUXNOT
    );
  tx_output_crc_loigc_Mxor_CO_14_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_Mxor_CO_13_Xo(2),
      ADR1 => tx_output_crc_loigc_n0104(0),
      ADR2 => tx_output_crcl(26),
      ADR3 => tx_output_crc_loigc_N81257,
      O => tx_output_crcl_14_FROM
    );
  tx_output_n0034_14_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_14_Q,
      O => tx_output_n0034_14_Q
    );
  tx_output_crcl_14_XUSED : X_BUF
    port map (
      I => tx_output_crcl_14_FROM,
      O => tx_output_crc_14_Q
    );
  mac_control_sclkdeltal_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_sclkdeltal_CEMUXNOT
    );
  rx_input_memio_crccomb_Mxor_CO_7_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0124(0),
      ADR1 => rx_input_memio_crccomb_Mxor_CO_7_Xo(1),
      ADR2 => rx_input_memio_crccomb_n0118(0),
      ADR3 => rx_input_memio_crccomb_n0118(1),
      O => rx_input_memio_crcl_7_FROM
    );
  rx_input_memio_n0048_7_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_7_Q,
      O => rx_input_memio_n0048_7_Q
    );
  rx_input_memio_crcl_7_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_7_FROM,
      O => rx_input_memio_crc_7_Q
    );
  rx_input_fifo_control_cs_FFd4_In_SW0 : X_LUT4
    generic map(
      INIT => X"FAFA"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd1,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_cs_FFd2,
      ADR3 => VCC,
      O => rx_input_fifo_control_cs_FFd4_FROM
    );
  rx_input_fifo_control_cs_FFd4_In_1595 : X_LUT4
    generic map(
      INIT => X"0F0E"
    )
    port map (
      ADR0 => rx_input_fifo_control_cs_FFd4,
      ADR1 => rx_input_fifo_control_cs_FFd3,
      ADR2 => rx_input_ce,
      ADR3 => rx_input_fifo_control_N70466,
      O => rx_input_fifo_control_cs_FFd4_In
    );
  rx_input_fifo_control_cs_FFd4_XUSED : X_BUF
    port map (
      I => rx_input_fifo_control_cs_FFd4_FROM,
      O => rx_input_fifo_control_N70466
    );
  mac_control_txfifowerr_cntl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_1_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_3_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_5_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_7_CEMUXNOT
    );
  mac_control_txfifowerr_cntl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txfifowerr_cntl_9_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(21),
      CE => mac_control_rxfifowerr_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_21_FFX_RST,
      O => mac_control_rxfifowerr_cntl(21)
    );
  mac_control_rxfifowerr_cntl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_21_FFX_RST
    );
  tx_output_crc_loigc_Mxor_CO_23_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_Mxor_CO_23_Xo(0),
      ADR1 => tx_output_crcl(30),
      ADR2 => tx_output_data(1),
      ADR3 => tx_output_crcl(15),
      O => tx_output_crcl_23_FROM
    );
  tx_output_n0034_23_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16_1,
      ADR3 => tx_output_crc_23_Q,
      O => tx_output_n0034_23_Q
    );
  tx_output_crcl_23_XUSED : X_BUF
    port map (
      I => tx_output_crcl_23_FROM,
      O => tx_output_crc_23_Q
    );
  rx_input_memio_crccomb_Mxor_CO_10_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_Mxor_CO_7_Xo(1),
      ADR1 => rx_input_memio_crcl(2),
      ADR2 => rx_input_memio_crccomb_n0118(1),
      ADR3 => rx_input_memio_crccomb_n0118(0),
      O => rx_input_memio_crcl_10_FROM
    );
  rx_input_memio_n0048_10_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_10_Q,
      O => rx_input_memio_n0048_10_Q
    );
  rx_input_memio_crcl_10_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_10_FROM,
      O => rx_input_memio_crc_10_Q
    );
  rx_input_memio_crccomb_Mxor_CO_8_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0115(0),
      ADR1 => rx_input_memio_crccomb_n0122(0),
      ADR2 => rx_input_memio_crcl(0),
      ADR3 => rx_input_memio_crccomb_Mxor_CO_7_Xo(1),
      O => rx_input_memio_crcl_8_FROM
    );
  rx_input_memio_n0048_8_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_8_Q,
      O => rx_input_memio_n0048_8_1_O
    );
  rx_input_memio_crcl_8_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_8_FROM,
      O => rx_input_memio_crc_8_Q
    );
  memcontroller_dnl2_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_11_CEMUXNOT
    );
  memcontroller_dnl2_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_21_CEMUXNOT
    );
  memcontroller_dnl2_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_13_CEMUXNOT
    );
  memcontroller_dnl2_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_23_CEMUXNOT
    );
  mac_control_rxfifowerr_cntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(13),
      CE => mac_control_rxfifowerr_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_13_FFX_RST,
      O => mac_control_rxfifowerr_cntl(13)
    );
  mac_control_rxfifowerr_cntl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_13_FFX_RST
    );
  memcontroller_dnl2_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_15_CEMUXNOT
    );
  memcontroller_dnl2_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_31_CEMUXNOT
    );
  memcontroller_dnl2_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_25_CEMUXNOT
    );
  memcontroller_dnl2_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_17_CEMUXNOT
    );
  memcontroller_dnl2_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_27_CEMUXNOT
    );
  memcontroller_dnl2_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_19_CEMUXNOT
    );
  memcontroller_dnl2_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_dnl2_29_CEMUXNOT
    );
  rx_input_memio_datal_1_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_datal_1_CEMUXNOT
    );
  rx_input_memio_datal_3_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_datal_3_CEMUXNOT
    );
  rx_input_memio_datal_5_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_datal_5_CEMUXNOT
    );
  rx_input_memio_datal_7_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_datal_7_CEMUXNOT
    );
  rx_input_memio_addrchk_lmaceq_0_rt_1596 : X_XOR2
    port map (
      I0 => rx_input_memio_addrchk_maceq_0_CYINIT,
      I1 => rx_input_memio_addrchk_maceq_0_FROM,
      O => rx_input_memio_addrchk_lmaceq_0_rt
    );
  rx_input_memio_addrchk_maceq_0_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_maceq_0_FROM
    );
  rx_input_memio_addrchk_maceq_0_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_maceq_0_CEMUXNOT
    );
  rx_input_memio_addrchk_maceq_0_CYINIT_1597 : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq(0),
      O => rx_input_memio_addrchk_maceq_0_CYINIT
    );
  rx_input_memio_addrchk_maceq_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_2_FFY_RST
    );
  rx_input_memio_addrchk_maceq_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq(3),
      CE => rx_input_memio_addrchk_maceq_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_2_FFY_RST,
      O => rx_input_memio_addrchk_maceq(3)
    );
  rx_input_memio_addrchk_lmaceq_2_rt_1598 : X_XOR2
    port map (
      I0 => rx_input_memio_addrchk_maceq_2_CYINIT,
      I1 => rx_input_memio_addrchk_maceq_2_FROM,
      O => rx_input_memio_addrchk_lmaceq_2_rt
    );
  rx_input_memio_addrchk_maceq_2_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_maceq_2_FROM
    );
  rx_input_memio_addrchk_maceq_2_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_maceq_2_CEMUXNOT
    );
  rx_input_memio_addrchk_maceq_2_CYINIT_1599 : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq(2),
      O => rx_input_memio_addrchk_maceq_2_CYINIT
    );
  mac_control_rxfifowerr_cntl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(31),
      CE => mac_control_rxfifowerr_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_31_FFX_RST,
      O => mac_control_rxfifowerr_cntl(31)
    );
  mac_control_rxfifowerr_cntl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_31_FFX_RST
    );
  rx_input_memio_addrchk_maceq_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_4_FFY_RST
    );
  rx_input_memio_addrchk_maceq_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq(5),
      CE => rx_input_memio_addrchk_maceq_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_4_FFY_RST,
      O => rx_input_memio_addrchk_maceq(5)
    );
  rx_input_memio_addrchk_lmaceq_4_rt_1600 : X_XOR2
    port map (
      I0 => rx_input_memio_addrchk_maceq_4_CYINIT,
      I1 => rx_input_memio_addrchk_maceq_4_FROM,
      O => rx_input_memio_addrchk_lmaceq_4_rt
    );
  rx_input_memio_addrchk_maceq_4_F : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_maceq_4_FROM
    );
  rx_input_memio_addrchk_maceq_4_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_maceq_4_CEMUXNOT
    );
  rx_input_memio_addrchk_maceq_4_CYINIT_1601 : X_BUF
    port map (
      I => rx_input_memio_addrchk_lmaceq(4),
      O => rx_input_memio_addrchk_maceq_4_CYINIT
    );
  mac_control_PHY_status_done_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_done_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd2,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_done_FFY_RST,
      O => mac_control_PHY_status_done
    );
  tx_output_crc_loigc_Mxor_CO_24_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0124(0),
      ADR1 => tx_output_crc_loigc_n0122(0),
      ADR2 => tx_output_crc_loigc_n0118(1),
      ADR3 => tx_output_crcl(16),
      O => tx_output_crcl_24_FROM
    );
  tx_output_n0034_24_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16_1,
      ADR3 => tx_output_crc_24_Q,
      O => tx_output_n0034_24_Q
    );
  tx_output_crcl_24_XUSED : X_BUF
    port map (
      I => tx_output_crcl_24_FROM,
      O => tx_output_crc_24_Q
    );
  tx_output_crc_loigc_Mxor_CO_16_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0118(0),
      ADR1 => tx_output_crcl(8),
      ADR2 => tx_output_crc_loigc_n0115(0),
      ADR3 => tx_output_crc_loigc_n0122(1),
      O => tx_output_crcl_16_FROM
    );
  tx_output_n0034_16_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16_1,
      ADR2 => VCC,
      ADR3 => tx_output_crc_16_Q,
      O => tx_output_n0034_16_1_O
    );
  tx_output_crcl_16_XUSED : X_BUF
    port map (
      I => tx_output_crcl_16_FROM,
      O => tx_output_crc_16_Q
    );
  rx_input_memio_crccomb_Mxor_CO_11_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_Mxor_CO_23_Xo(0),
      ADR1 => rx_input_memio_crcl(3),
      ADR2 => rx_input_memio_crccomb_n0115(0),
      ADR3 => rx_input_memio_crccomb_n0124(1),
      O => rx_input_memio_crcl_11_FROM
    );
  rx_input_memio_n0048_11_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_11_Q,
      O => rx_input_memio_n0048_11_1_O
    );
  rx_input_memio_crcl_11_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_11_FROM,
      O => rx_input_memio_crc_11_Q
    );
  mac_control_PHY_status_n00111 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => RESET_IBUF,
      ADR2 => VCC,
      ADR3 => mac_control_PHY_status_cs_FFd4,
      O => mac_control_PHY_status_n0011_GROM
    );
  mac_control_PHY_status_n0011_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_n0011_GROM,
      O => mac_control_PHY_status_n0011
    );
  mac_control_PHY_status_miiaddr_1_1 : X_LUT4
    generic map(
      INIT => X"FFF8"
    )
    port map (
      ADR0 => mac_control_PHY_status_N43105,
      ADR1 => mac_control_PHY_status_addrl(1),
      ADR2 => mac_control_PHY_status_cs_FFd6,
      ADR3 => mac_control_PHY_status_cs_FFd5,
      O => mac_control_PHY_status_miiaddr_1_FROM
    );
  mac_control_PHY_status_n00201 : X_LUT4
    generic map(
      INIT => X"5040"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => mac_control_PHY_status_cs_FFd6,
      ADR2 => mac_control_PHY_status_done,
      ADR3 => mac_control_PHY_status_cs_FFd5,
      O => mac_control_PHY_status_miiaddr_1_GROM
    );
  mac_control_PHY_status_miiaddr_1_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_1_FROM,
      O => mac_control_PHY_status_miiaddr(1)
    );
  mac_control_PHY_status_miiaddr_1_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_1_GROM,
      O => mac_control_PHY_status_n0020
    );
  rx_input_memio_crccomb_Mxor_CO_9_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(1),
      ADR1 => rx_input_memio_crccomb_n0118(1),
      ADR2 => rx_input_memio_crccomb_n0118(0),
      ADR3 => rx_input_memio_crccomb_Mxor_CO_9_Xo(0),
      O => rx_input_memio_crcl_9_FROM
    );
  rx_input_memio_n0048_9_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_9_Q,
      O => rx_input_memio_n0048_9_Q
    );
  rx_input_memio_crcl_9_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_9_FROM,
      O => rx_input_memio_crc_9_Q
    );
  mac_control_sclkdeltall_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_sclkdeltall_CEMUXNOT
    );
  mac_control_phyaddr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_13_FFY_RST
    );
  mac_control_phyaddr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_13_FFY_RST,
      O => mac_control_phyaddr(12)
    );
  mac_control_phyaddr_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_21_FFY_RST
    );
  mac_control_phyaddr_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(20),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_21_FFY_RST,
      O => mac_control_phyaddr(20)
    );
  mac_control_phyaddr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_15_FFY_RST
    );
  mac_control_phyaddr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_15_FFY_RST,
      O => mac_control_phyaddr(14)
    );
  mac_control_rxfifowerr_cntl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(23),
      CE => mac_control_rxfifowerr_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_23_FFX_RST,
      O => mac_control_rxfifowerr_cntl(23)
    );
  mac_control_rxfifowerr_cntl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_23_FFX_RST
    );
  mac_control_phyaddr_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_30_FFY_RST
    );
  mac_control_phyaddr_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(30),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_30_FFY_RST,
      O => mac_control_phyaddr(30)
    );
  mac_control_phyaddr_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_25_FFY_RST
    );
  mac_control_phyaddr_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(24),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_25_FFY_RST,
      O => mac_control_phyaddr(24)
    );
  mac_control_phyaddr_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_19_FFY_RST
    );
  mac_control_phyaddr_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(18),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_19_FFY_RST,
      O => mac_control_phyaddr(18)
    );
  mac_control_phyaddr_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_27_FFY_RST
    );
  mac_control_phyaddr_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(26),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_27_FFY_RST,
      O => mac_control_phyaddr(26)
    );
  mac_control_phyaddr_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_29_FFY_RST
    );
  mac_control_phyaddr_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(28),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_29_FFY_RST,
      O => mac_control_phyaddr(28)
    );
  rx_input_memio_addrchk_datal_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_11_FFY_RST
    );
  rx_input_memio_addrchk_datal_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_11_FFY_RST,
      O => rx_input_memio_addrchk_datal(10)
    );
  mac_control_rxfifowerr_cntl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(24),
      CE => mac_control_rxfifowerr_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_25_FFY_RST,
      O => mac_control_rxfifowerr_cntl(24)
    );
  mac_control_rxfifowerr_cntl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_25_FFY_RST
    );
  mac_control_rxfifowerr_cntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(15),
      CE => mac_control_rxfifowerr_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_15_FFX_RST,
      O => mac_control_rxfifowerr_cntl(15)
    );
  mac_control_rxfifowerr_cntl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_15_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_35_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_34 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(34),
      CE => rx_input_memio_addrchk_macaddrl_35_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_35_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(34)
    );
  rx_input_memio_addrchk_macaddrl_35_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_35_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_27_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(26),
      CE => rx_input_memio_addrchk_macaddrl_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_27_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(26)
    );
  rx_input_memio_addrchk_macaddrl_27_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_27_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_19_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_19_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_45_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_44 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(44),
      CE => rx_input_memio_addrchk_macaddrl_45_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_45_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(44)
    );
  rx_input_memio_addrchk_macaddrl_45_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_45_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_37_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_37_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_36 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(36),
      CE => rx_input_memio_addrchk_macaddrl_37_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_37_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(36)
    );
  rx_input_memio_addrchk_macaddrl_37_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_37_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_29_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(28),
      CE => rx_input_memio_addrchk_macaddrl_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_29_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(28)
    );
  rx_input_memio_addrchk_macaddrl_29_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_29_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_47_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_46 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(46),
      CE => rx_input_memio_addrchk_macaddrl_47_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_47_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(46)
    );
  rx_input_memio_addrchk_macaddrl_47_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_47_CEMUXNOT
    );
  rx_input_memio_addrchk_macaddrl_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_39_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_38 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(38),
      CE => rx_input_memio_addrchk_macaddrl_39_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_39_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(38)
    );
  rx_input_memio_addrchk_macaddrl_39_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_macaddrl_39_CEMUXNOT
    );
  mac_control_Mmux_n0016_Result_10_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0062,
      ADR1 => mac_control_rxf_cntl(10),
      ADR2 => mac_control_txf_cntl(10),
      ADR3 => mac_control_n0061,
      O => mac_control_CHOICE2745_FROM
    );
  mac_control_Mmux_n0016_Result_10_48_SW0 : X_LUT4
    generic map(
      INIT => X"FFEC"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cntl(10),
      ADR1 => mac_control_n0056,
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_CHOICE2745,
      O => mac_control_CHOICE2745_GROM
    );
  mac_control_CHOICE2745_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2745_FROM,
      O => mac_control_CHOICE2745
    );
  mac_control_CHOICE2745_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2745_GROM,
      O => mac_control_N81058
    );
  mac_control_Mmux_n0016_Result_17_30 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_phyaddr(17),
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_n00851_1,
      ADR3 => mac_control_txfifowerr_cntl(17),
      O => mac_control_CHOICE2348_FROM
    );
  mac_control_Mmux_n0016_Result_10_30 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_txfifowerr_cntl(10),
      ADR3 => mac_control_phyaddr(10),
      O => mac_control_CHOICE2348_GROM
    );
  mac_control_CHOICE2348_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2348_FROM,
      O => mac_control_CHOICE2348
    );
  mac_control_CHOICE2348_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2348_GROM,
      O => mac_control_CHOICE2750
    );
  mac_control_Mmux_n0016_Result_19_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txfifowerr_cntl(19),
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_rxfifowerr_cntl(19),
      ADR3 => mac_control_n0064,
      O => mac_control_CHOICE2085_FROM
    );
  mac_control_Mmux_n0016_Result_11_10 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cntl(11),
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_txfifowerr_cntl(11),
      ADR3 => mac_control_n0064,
      O => mac_control_CHOICE2085_GROM
    );
  mac_control_CHOICE2085_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2085_FROM,
      O => mac_control_CHOICE2085
    );
  mac_control_CHOICE2085_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2085_GROM,
      O => mac_control_CHOICE2486
    );
  mac_control_Mmux_n0016_Result_26_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_phyaddr(26),
      ADR2 => mac_control_n0065,
      ADR3 => mac_control_rxphyerr_cntl(26),
      O => mac_control_CHOICE2181_FROM
    );
  mac_control_Mmux_n0016_Result_11_22 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_phyaddr(11),
      ADR1 => mac_control_rxphyerr_cntl(11),
      ADR2 => mac_control_n00851_1,
      ADR3 => mac_control_n0065,
      O => mac_control_CHOICE2181_GROM
    );
  mac_control_CHOICE2181_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2181_FROM,
      O => mac_control_CHOICE2181
    );
  mac_control_CHOICE2181_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2181_GROM,
      O => mac_control_CHOICE2490
    );
  mac_control_Mmux_n0016_Result_10_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2741,
      ADR1 => mac_control_CHOICE2750,
      ADR2 => mac_control_CHOICE2738,
      ADR3 => mac_control_N81058,
      O => mac_control_CHOICE2753_FROM
    );
  mac_control_Mmux_n0016_Result_10_60 : X_LUT4
    generic map(
      INIT => X"FF88"
    )
    port map (
      ADR0 => mac_control_phystat(10),
      ADR1 => mac_control_n0057,
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2753,
      O => mac_control_CHOICE2753_GROM
    );
  mac_control_CHOICE2753_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2753_FROM,
      O => mac_control_CHOICE2753
    );
  mac_control_CHOICE2753_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2753_GROM,
      O => mac_control_CHOICE2755
    );
  mac_control_Mmux_n0016_Result_15_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0063,
      ADR1 => mac_control_n0064,
      ADR2 => mac_control_txfifowerr_cntl(15),
      ADR3 => mac_control_rxfifowerr_cntl(15),
      O => mac_control_CHOICE2586_FROM
    );
  mac_control_Mmux_n0016_Result_20_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_txfifowerr_cntl(20),
      ADR2 => mac_control_rxfifowerr_cntl(20),
      ADR3 => mac_control_n0063,
      O => mac_control_CHOICE2586_GROM
    );
  mac_control_CHOICE2586_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2586_FROM,
      O => mac_control_CHOICE2586
    );
  mac_control_CHOICE2586_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2586_GROM,
      O => mac_control_CHOICE2131
    );
  mac_control_Mmux_n0016_Result_11_28 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0061,
      ADR1 => mac_control_n0066,
      ADR2 => mac_control_txf_cntl(11),
      ADR3 => mac_control_rxoferr_cntl(11),
      O => mac_control_CHOICE2494_FROM
    );
  mac_control_Mmux_n0016_Result_11_45_SW0 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_n0059,
      ADR1 => VCC,
      ADR2 => mac_control_phydi(11),
      ADR3 => mac_control_CHOICE2494,
      O => mac_control_CHOICE2494_GROM
    );
  mac_control_CHOICE2494_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2494_FROM,
      O => mac_control_CHOICE2494
    );
  mac_control_CHOICE2494_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2494_GROM,
      O => mac_control_N81110
    );
  mac_control_Mmux_n0016_Result_11_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_N81110,
      ADR1 => mac_control_CHOICE2483,
      ADR2 => mac_control_CHOICE2486,
      ADR3 => mac_control_CHOICE2490,
      O => mac_control_CHOICE2497_FROM
    );
  mac_control_Mmux_n0016_Result_11_56 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_phystat(11),
      ADR1 => VCC,
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_CHOICE2497,
      O => mac_control_CHOICE2497_GROM
    );
  mac_control_CHOICE2497_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2497_FROM,
      O => mac_control_CHOICE2497
    );
  mac_control_CHOICE2497_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2497_GROM,
      O => mac_control_CHOICE2499
    );
  mac_control_Mmux_n0016_Result_19_22 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_phyaddr(19),
      ADR1 => mac_control_rxphyerr_cntl(19),
      ADR2 => mac_control_n00851_1,
      ADR3 => mac_control_n0065,
      O => mac_control_CHOICE2089_FROM
    );
  mac_control_Mmux_n0016_Result_20_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0065,
      ADR1 => mac_control_n00851_1,
      ADR2 => mac_control_phyaddr(20),
      ADR3 => mac_control_rxphyerr_cntl(20),
      O => mac_control_CHOICE2089_GROM
    );
  mac_control_CHOICE2089_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2089_FROM,
      O => mac_control_CHOICE2089
    );
  mac_control_CHOICE2089_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2089_GROM,
      O => mac_control_CHOICE2135
    );
  tx_output_crc_loigc_Mxor_CO_28_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(20),
      ADR1 => tx_output_crc_loigc_n0118(1),
      ADR2 => tx_output_crc_loigc_n0118(0),
      ADR3 => tx_output_crc_loigc_n0104(0),
      O => tx_output_crcl_28_FROM
    );
  tx_output_n0034_28_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_output_cs_FFd16_1,
      ADR2 => VCC,
      ADR3 => tx_output_crc_28_Q,
      O => tx_output_n0034_28_Q
    );
  tx_output_crcl_28_XUSED : X_BUF
    port map (
      I => tx_output_crcl_28_FROM,
      O => tx_output_crc_28_Q
    );
  mac_control_Mmux_n0016_Result_16_10 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phydi(16),
      ADR1 => mac_control_n0066,
      ADR2 => mac_control_rxoferr_cntl(16),
      ADR3 => mac_control_n0059,
      O => mac_control_CHOICE2315_FROM
    );
  mac_control_Mmux_n0016_Result_21_10 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0066,
      ADR1 => mac_control_n0059,
      ADR2 => mac_control_phydi(21),
      ADR3 => mac_control_rxoferr_cntl(21),
      O => mac_control_CHOICE2315_GROM
    );
  mac_control_CHOICE2315_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2315_FROM,
      O => mac_control_CHOICE2315
    );
  mac_control_CHOICE2315_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2315_GROM,
      O => mac_control_CHOICE2363
    );
  tx_output_crcl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_8_1_O,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_8_FFY_RST,
      O => tx_output_crcl(8)
    );
  tx_output_crcl_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_8_FFY_RST
    );
  mac_control_Mmux_n0016_Result_18_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_rxfifowerr_cntl(18),
      ADR3 => mac_control_txfifowerr_cntl(18),
      O => mac_control_CHOICE2062_FROM
    );
  mac_control_Mmux_n0016_Result_13_10 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxfifowerr_cntl(13),
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_txfifowerr_cntl(13),
      ADR3 => mac_control_n0064,
      O => mac_control_CHOICE2062_GROM
    );
  mac_control_CHOICE2062_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2062_FROM,
      O => mac_control_CHOICE2062
    );
  mac_control_CHOICE2062_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2062_GROM,
      O => mac_control_CHOICE2561
    );
  mac_control_Mmux_n0016_Result_12_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxoferr_cntl(12),
      ADR1 => mac_control_n0066,
      ADR2 => mac_control_txf_cntl(12),
      ADR3 => mac_control_n0061,
      O => mac_control_CHOICE2544_FROM
    );
  mac_control_Mmux_n0016_Result_12_45_SW0 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_n0059,
      ADR1 => VCC,
      ADR2 => mac_control_phydi(12),
      ADR3 => mac_control_CHOICE2544,
      O => mac_control_CHOICE2544_GROM
    );
  mac_control_CHOICE2544_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2544_FROM,
      O => mac_control_CHOICE2544
    );
  mac_control_CHOICE2544_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2544_GROM,
      O => mac_control_N81138
    );
  mac_control_Mmux_n0016_Result_12_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_N81138,
      ADR1 => mac_control_CHOICE2536,
      ADR2 => mac_control_CHOICE2540,
      ADR3 => mac_control_CHOICE2533,
      O => mac_control_CHOICE2547_FROM
    );
  mac_control_Mmux_n0016_Result_12_56 : X_LUT4
    generic map(
      INIT => X"FFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_phystat(12),
      ADR2 => mac_control_n0057,
      ADR3 => mac_control_CHOICE2547,
      O => mac_control_CHOICE2547_GROM
    );
  mac_control_CHOICE2547_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2547_FROM,
      O => mac_control_CHOICE2547
    );
  mac_control_CHOICE2547_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2547_GROM,
      O => mac_control_CHOICE2549
    );
  mac_control_Mmux_n0016_Result_17_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cntl(17),
      ADR1 => mac_control_n0061,
      ADR2 => mac_control_rxf_cntl(17),
      ADR3 => mac_control_n0062,
      O => mac_control_CHOICE2343_FROM
    );
  mac_control_Mmux_n0016_Result_21_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cntl(21),
      ADR1 => mac_control_n0061,
      ADR2 => mac_control_n0062,
      ADR3 => mac_control_rxf_cntl(21),
      O => mac_control_CHOICE2343_GROM
    );
  mac_control_CHOICE2343_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2343_FROM,
      O => mac_control_CHOICE2343
    );
  mac_control_CHOICE2343_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2343_GROM,
      O => mac_control_CHOICE2367
    );
  mac_control_Mmux_n0016_Result_15_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cntl(15),
      ADR1 => mac_control_n0065,
      ADR2 => mac_control_phyaddr(15),
      ADR3 => mac_control_n00851_1,
      O => mac_control_CHOICE2590_FROM
    );
  mac_control_Mmux_n0016_Result_13_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cntl(13),
      ADR1 => mac_control_n00851_1,
      ADR2 => mac_control_phyaddr(13),
      ADR3 => mac_control_n0065,
      O => mac_control_CHOICE2590_GROM
    );
  mac_control_CHOICE2590_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2590_FROM,
      O => mac_control_CHOICE2590
    );
  mac_control_CHOICE2590_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2590_GROM,
      O => mac_control_CHOICE2565
    );
  mac_control_Mmux_n0016_Result_17_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0066,
      ADR1 => mac_control_phydi(17),
      ADR2 => mac_control_rxoferr_cntl(17),
      ADR3 => mac_control_n0059,
      O => mac_control_CHOICE2339_FROM
    );
  mac_control_Mmux_n0016_Result_14_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phydi(14),
      ADR1 => mac_control_n0059,
      ADR2 => mac_control_rxoferr_cntl(14),
      ADR3 => mac_control_n0066,
      O => mac_control_CHOICE2339_GROM
    );
  mac_control_CHOICE2339_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2339_FROM,
      O => mac_control_CHOICE2339
    );
  mac_control_CHOICE2339_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2339_GROM,
      O => mac_control_CHOICE2767
    );
  mac_control_Mmux_n0016_Result_13_28 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0061,
      ADR1 => mac_control_n0066,
      ADR2 => mac_control_txf_cntl(13),
      ADR3 => mac_control_rxoferr_cntl(13),
      O => mac_control_CHOICE2569_FROM
    );
  mac_control_Mmux_n0016_Result_13_45_SW0 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_n0059,
      ADR1 => VCC,
      ADR2 => mac_control_phydi(13),
      ADR3 => mac_control_CHOICE2569,
      O => mac_control_CHOICE2569_GROM
    );
  mac_control_CHOICE2569_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2569_FROM,
      O => mac_control_CHOICE2569
    );
  mac_control_CHOICE2569_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2569_GROM,
      O => mac_control_N81082
    );
  mac_control_Mmux_n0016_Result_13_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2558,
      ADR1 => mac_control_N81082,
      ADR2 => mac_control_CHOICE2561,
      ADR3 => mac_control_CHOICE2565,
      O => mac_control_CHOICE2572_FROM
    );
  mac_control_Mmux_n0016_Result_13_56 : X_LUT4
    generic map(
      INIT => X"FF88"
    )
    port map (
      ADR0 => mac_control_n0057,
      ADR1 => mac_control_phystat(13),
      ADR2 => VCC,
      ADR3 => mac_control_CHOICE2572,
      O => mac_control_CHOICE2572_GROM
    );
  mac_control_CHOICE2572_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2572_FROM,
      O => mac_control_CHOICE2572
    );
  mac_control_CHOICE2572_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2572_GROM,
      O => mac_control_CHOICE2574
    );
  mac_control_Mmux_n0016_Result_14_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0062,
      ADR1 => mac_control_txf_cntl(14),
      ADR2 => mac_control_n0061,
      ADR3 => mac_control_rxf_cntl(14),
      O => mac_control_CHOICE2771_FROM
    );
  mac_control_Mmux_n0016_Result_14_48_SW0 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_n0056,
      ADR1 => mac_control_rxcrcerr_cntl(14),
      ADR2 => mac_control_n0067,
      ADR3 => mac_control_CHOICE2771,
      O => mac_control_CHOICE2771_GROM
    );
  mac_control_CHOICE2771_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2771_FROM,
      O => mac_control_CHOICE2771
    );
  mac_control_CHOICE2771_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2771_GROM,
      O => mac_control_N81042
    );
  mac_control_Mmux_n0016_Result_23_10 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_txfifowerr_cntl(23),
      ADR3 => mac_control_rxfifowerr_cntl(23),
      O => mac_control_CHOICE2154_FROM
    );
  mac_control_Mmux_n0016_Result_14_30 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0063,
      ADR1 => mac_control_n00851_1,
      ADR2 => mac_control_phyaddr(14),
      ADR3 => mac_control_txfifowerr_cntl(14),
      O => mac_control_CHOICE2154_GROM
    );
  mac_control_CHOICE2154_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2154_FROM,
      O => mac_control_CHOICE2154
    );
  mac_control_CHOICE2154_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2154_GROM,
      O => mac_control_CHOICE2776
    );
  mac_control_Mmux_n0016_Result_18_22 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_rxphyerr_cntl(18),
      ADR2 => mac_control_phyaddr(18),
      ADR3 => mac_control_n0065,
      O => mac_control_CHOICE2066_FROM
    );
  mac_control_Mmux_n0016_Result_22_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0065,
      ADR1 => mac_control_rxphyerr_cntl(22),
      ADR2 => mac_control_phyaddr(22),
      ADR3 => mac_control_n00851_1,
      O => mac_control_CHOICE2066_GROM
    );
  mac_control_CHOICE2066_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2066_FROM,
      O => mac_control_CHOICE2066
    );
  mac_control_CHOICE2066_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2066_GROM,
      O => mac_control_CHOICE2112
    );
  mac_control_Mmux_n0016_Result_27_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_n0063,
      ADR2 => mac_control_rxfifowerr_cntl(27),
      ADR3 => mac_control_txfifowerr_cntl(27),
      O => mac_control_CHOICE2223_FROM
    );
  mac_control_Mmux_n0016_Result_31_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0062,
      ADR1 => mac_control_txfifowerr_cntl(31),
      ADR2 => mac_control_rxf_cntl(31),
      ADR3 => mac_control_n0063,
      O => mac_control_CHOICE2223_GROM
    );
  mac_control_CHOICE2223_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2223_FROM,
      O => mac_control_CHOICE2223
    );
  mac_control_CHOICE2223_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2223_GROM,
      O => mac_control_CHOICE2039
    );
  mac_control_Mmux_n0016_Result_19_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cntl(19),
      ADR1 => mac_control_n0061,
      ADR2 => mac_control_rxoferr_cntl(19),
      ADR3 => mac_control_n0066,
      O => mac_control_CHOICE2093_FROM
    );
  mac_control_Mmux_n0016_Result_22_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0061,
      ADR1 => mac_control_txf_cntl(22),
      ADR2 => mac_control_n0066,
      ADR3 => mac_control_rxoferr_cntl(22),
      O => mac_control_CHOICE2093_GROM
    );
  mac_control_CHOICE2093_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2093_FROM,
      O => mac_control_CHOICE2093
    );
  mac_control_CHOICE2093_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2093_GROM,
      O => mac_control_CHOICE2116
    );
  mac_control_Mmux_n0016_Result_18_28 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_txf_cntl(18),
      ADR1 => mac_control_rxoferr_cntl(18),
      ADR2 => mac_control_n0066,
      ADR3 => mac_control_n0061,
      O => mac_control_CHOICE2070_FROM
    );
  mac_control_Mmux_n0016_Result_30_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0066,
      ADR1 => mac_control_rxoferr_cntl(30),
      ADR2 => mac_control_n0061,
      ADR3 => mac_control_txf_cntl(30),
      O => mac_control_CHOICE2070_GROM
    );
  mac_control_CHOICE2070_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2070_FROM,
      O => mac_control_CHOICE2070
    );
  mac_control_CHOICE2070_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2070_GROM,
      O => mac_control_CHOICE2300
    );
  mac_control_Mmux_n0016_Result_27_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_phyaddr(27),
      ADR2 => mac_control_n0065,
      ADR3 => mac_control_rxphyerr_cntl(27),
      O => mac_control_CHOICE2227_FROM
    );
  mac_control_Mmux_n0016_Result_23_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n00851_1,
      ADR1 => mac_control_n0065,
      ADR2 => mac_control_rxphyerr_cntl(23),
      ADR3 => mac_control_phyaddr(23),
      O => mac_control_CHOICE2227_GROM
    );
  mac_control_CHOICE2227_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2227_FROM,
      O => mac_control_CHOICE2227
    );
  mac_control_CHOICE2227_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2227_GROM,
      O => mac_control_CHOICE2158
    );
  mac_control_Mmux_n0016_Result_14_48 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_N81042,
      ADR1 => mac_control_CHOICE2767,
      ADR2 => mac_control_CHOICE2776,
      ADR3 => mac_control_CHOICE2764,
      O => mac_control_CHOICE2779_FROM
    );
  mac_control_Mmux_n0016_Result_14_60 : X_LUT4
    generic map(
      INIT => X"FFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0057,
      ADR2 => mac_control_phystat(14),
      ADR3 => mac_control_CHOICE2779,
      O => mac_control_CHOICE2779_GROM
    );
  mac_control_CHOICE2779_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2779_FROM,
      O => mac_control_CHOICE2779
    );
  mac_control_CHOICE2779_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2779_GROM,
      O => mac_control_CHOICE2781
    );
  mac_control_Mmux_n0016_Result_27_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_txf_cntl(27),
      ADR1 => mac_control_n0061,
      ADR2 => mac_control_n0066,
      ADR3 => mac_control_rxoferr_cntl(27),
      O => mac_control_CHOICE2231_FROM
    );
  mac_control_Mmux_n0016_Result_31_27 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxcrcerr_cntl(31),
      ADR1 => mac_control_n0067,
      ADR2 => mac_control_n0066,
      ADR3 => mac_control_rxoferr_cntl(31),
      O => mac_control_CHOICE2231_GROM
    );
  mac_control_CHOICE2231_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2231_FROM,
      O => mac_control_CHOICE2231
    );
  mac_control_CHOICE2231_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2231_GROM,
      O => mac_control_CHOICE2046
    );
  mac_control_Mmux_n0016_Result_15_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxoferr_cntl(15),
      ADR1 => mac_control_n0066,
      ADR2 => mac_control_n0061,
      ADR3 => mac_control_txf_cntl(15),
      O => mac_control_CHOICE2594_FROM
    );
  mac_control_Mmux_n0016_Result_15_45_SW0 : X_LUT4
    generic map(
      INIT => X"FFA0"
    )
    port map (
      ADR0 => mac_control_n0059,
      ADR1 => VCC,
      ADR2 => mac_control_phydi(15),
      ADR3 => mac_control_CHOICE2594,
      O => mac_control_CHOICE2594_GROM
    );
  mac_control_CHOICE2594_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2594_FROM,
      O => mac_control_CHOICE2594
    );
  mac_control_CHOICE2594_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2594_GROM,
      O => mac_control_N81118
    );
  mac_control_Mmux_n0016_Result_29_28 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0066,
      ADR1 => mac_control_txf_cntl(29),
      ADR2 => mac_control_rxoferr_cntl(29),
      ADR3 => mac_control_n0061,
      O => mac_control_CHOICE2277_FROM
    );
  mac_control_Mmux_n0016_Result_23_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0061,
      ADR1 => mac_control_txf_cntl(23),
      ADR2 => mac_control_n0066,
      ADR3 => mac_control_rxoferr_cntl(23),
      O => mac_control_CHOICE2277_GROM
    );
  mac_control_CHOICE2277_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2277_FROM,
      O => mac_control_CHOICE2277
    );
  mac_control_CHOICE2277_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2277_GROM,
      O => mac_control_CHOICE2162
    );
  mac_control_Mmux_n0016_Result_31_36 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2039,
      ADR1 => mac_control_CHOICE2046,
      ADR2 => mac_control_CHOICE2043,
      ADR3 => mac_control_N80963,
      O => mac_control_CHOICE2048_FROM
    );
  mac_control_Mmux_n0016_Result_31_85_SW0 : X_LUT4
    generic map(
      INIT => X"FFEA"
    )
    port map (
      ADR0 => mac_control_N81417,
      ADR1 => mac_control_n0057,
      ADR2 => mac_control_phystat(31),
      ADR3 => mac_control_CHOICE2048,
      O => mac_control_CHOICE2048_GROM
    );
  mac_control_CHOICE2048_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2048_FROM,
      O => mac_control_CHOICE2048
    );
  mac_control_CHOICE2048_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2048_GROM,
      O => mac_control_N81176
    );
  mac_control_Mmux_n0016_Result_15_45 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE2586,
      ADR1 => mac_control_CHOICE2583,
      ADR2 => mac_control_N81118,
      ADR3 => mac_control_CHOICE2590,
      O => mac_control_CHOICE2597_FROM
    );
  mac_control_Mmux_n0016_Result_15_56 : X_LUT4
    generic map(
      INIT => X"FFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_n0057,
      ADR2 => mac_control_phystat(15),
      ADR3 => mac_control_CHOICE2597,
      O => mac_control_CHOICE2597_GROM
    );
  mac_control_CHOICE2597_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2597_FROM,
      O => mac_control_CHOICE2597
    );
  mac_control_CHOICE2597_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2597_GROM,
      O => mac_control_CHOICE2599
    );
  mac_control_Mmux_n0016_Result_25_28 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0061,
      ADR1 => mac_control_txf_cntl(25),
      ADR2 => mac_control_rxoferr_cntl(25),
      ADR3 => mac_control_n0066,
      O => mac_control_CHOICE2208_FROM
    );
  mac_control_Mmux_n0016_Result_24_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_n0061,
      ADR1 => mac_control_n0062,
      ADR2 => mac_control_rxf_cntl(24),
      ADR3 => mac_control_txf_cntl(24),
      O => mac_control_CHOICE2208_GROM
    );
  mac_control_CHOICE2208_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2208_FROM,
      O => mac_control_CHOICE2208
    );
  mac_control_CHOICE2208_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2208_GROM,
      O => mac_control_CHOICE2391
    );
  mac_control_Mmux_n0016_Result_29_10 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_n0063,
      ADR1 => mac_control_txfifowerr_cntl(29),
      ADR2 => mac_control_n0064,
      ADR3 => mac_control_rxfifowerr_cntl(29),
      O => mac_control_CHOICE2269_FROM
    );
  mac_control_Mmux_n0016_Result_25_10 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0064,
      ADR1 => mac_control_txfifowerr_cntl(25),
      ADR2 => mac_control_rxfifowerr_cntl(25),
      ADR3 => mac_control_n0063,
      O => mac_control_CHOICE2269_GROM
    );
  mac_control_CHOICE2269_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2269_FROM,
      O => mac_control_CHOICE2269
    );
  mac_control_CHOICE2269_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2269_GROM,
      O => mac_control_CHOICE2200
    );
  mac_control_rxfifowerr_cntl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(25),
      CE => mac_control_rxfifowerr_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_25_FFX_RST,
      O => mac_control_rxfifowerr_cntl(25)
    );
  mac_control_rxfifowerr_cntl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_25_FFX_RST
    );
  rx_input_memio_crcll_1_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_1_CEMUXNOT
    );
  rx_input_memio_crcll_3_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_3_CEMUXNOT
    );
  rx_input_memio_crcll_5_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_5_CEMUXNOT
    );
  rx_input_memio_crcll_7_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_7_CEMUXNOT
    );
  rx_input_memio_crcll_9_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_9_CEMUXNOT
    );
  tx_output_ltxd_3_1 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => tx_output_outselll(0),
      ADR1 => tx_output_ncrcbytel(4),
      ADR2 => tx_output_outselll(3),
      ADR3 => tx_output_datal(3),
      O => tx_output_ltxd_3_FROM
    );
  tx_output_ltxd_1_1 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => tx_output_ncrcbytel(6),
      ADR1 => tx_output_outselll(3),
      ADR2 => tx_output_datal(1),
      ADR3 => tx_output_outselll(0),
      O => tx_output_ltxd_3_GROM
    );
  tx_output_ltxd_3_XUSED : X_BUF
    port map (
      I => tx_output_ltxd_3_FROM,
      O => tx_output_ltxd(3)
    );
  tx_output_ltxd_3_YUSED : X_BUF
    port map (
      I => tx_output_ltxd_3_GROM,
      O => tx_output_ltxd(1)
    );
  tx_output_ltxd_5_1 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => tx_output_outselll(0),
      ADR1 => tx_output_outselll(3),
      ADR2 => tx_output_ncrcbytel(2),
      ADR3 => tx_output_datal(5),
      O => tx_output_ltxd_5_GROM
    );
  tx_output_ltxd_5_YUSED : X_BUF
    port map (
      I => tx_output_ltxd_5_GROM,
      O => tx_output_ltxd(5)
    );
  tx_output_crc_loigc_Mxor_CO_25_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crcl(26),
      ADR1 => tx_output_data(5),
      ADR2 => tx_output_crcl(17),
      ADR3 => tx_output_crc_loigc_n0124(1),
      O => tx_output_crcl_25_FROM
    );
  tx_output_n0034_25_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_crc_25_Q,
      ADR3 => tx_output_cs_FFd16_1,
      O => tx_output_n0034_25_Q
    );
  tx_output_crcl_25_XUSED : X_BUF
    port map (
      I => tx_output_crcl_25_FROM,
      O => tx_output_crc_25_Q
    );
  mac_control_rxfifowerr_cntl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(17),
      CE => mac_control_rxfifowerr_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_17_FFX_RST,
      O => mac_control_rxfifowerr_cntl(17)
    );
  mac_control_rxfifowerr_cntl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_17_FFX_RST
    );
  tx_output_crc_loigc_Mxor_CO_17_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0118(0),
      ADR1 => tx_output_crc_loigc_n0104(0),
      ADR2 => tx_output_crc_loigc_n0122(0),
      ADR3 => tx_output_crcl(9),
      O => tx_output_crcl_17_FROM
    );
  tx_output_n0034_17_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => tx_output_cs_FFd16_1,
      ADR3 => tx_output_crc_17_Q,
      O => tx_output_n0034_17_Q
    );
  tx_output_crcl_17_XUSED : X_BUF
    port map (
      I => tx_output_crcl_17_FROM,
      O => tx_output_crc_17_Q
    );
  memcontroller_clknum_0_1_BYMUX : X_INV
    port map (
      I => memcontroller_clknum_0_1,
      O => memcontroller_clknum_0_1_BYMUXNOT
    );
  rx_input_memio_dout_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_21_FFY_RST
    );
  rx_input_memio_dout_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_21_FFY_RST,
      O => rx_input_memio_dout(20)
    );
  rx_input_memio_dout_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_13_FFY_RST
    );
  rx_input_memio_dout_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_13_FFY_RST,
      O => rx_input_memio_dout(12)
    );
  mac_control_PHY_status_MII_Interface_dreg_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_12_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(10),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_12_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(11)
    );
  mac_control_rxfifowerr_cntl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(18),
      CE => mac_control_rxfifowerr_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_19_FFY_RST,
      O => mac_control_rxfifowerr_cntl(18)
    );
  mac_control_rxfifowerr_cntl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_19_FFY_RST
    );
  rx_input_memio_dout_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_23_FFY_RST
    );
  rx_input_memio_dout_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_23_FFY_RST,
      O => rx_input_memio_dout(22)
    );
  rx_input_memio_dout_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_15_FFY_RST
    );
  rx_input_memio_dout_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_15_FFY_RST,
      O => rx_input_memio_dout(14)
    );
  mac_control_rxfifowerr_cntl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(27),
      CE => mac_control_rxfifowerr_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_27_FFX_RST,
      O => mac_control_rxfifowerr_cntl(27)
    );
  mac_control_rxfifowerr_cntl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_27_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_14_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(12),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_14_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(13)
    );
  rx_input_memio_dout_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_17_FFY_RST
    );
  rx_input_memio_dout_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_17_FFY_RST,
      O => rx_input_memio_dout(16)
    );
  mac_control_PHY_status_MII_Interface_dreg_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_15_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(14),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_15_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(15)
    );
  rx_input_memio_dout_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_19_FFY_RST
    );
  rx_input_memio_dout_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_19_FFY_RST,
      O => rx_input_memio_dout(18)
    );
  rx_input_memio_dout_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_29_FFY_RST
    );
  rx_input_memio_dout_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_29_FFY_RST,
      O => rx_input_memio_dout(28)
    );
  rx_input_memio_addrchk_validbcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_validbcast_FFY_RST
    );
  rx_input_memio_addrchk_validbcast_1602 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_n0051,
      CE => rx_input_memio_addrchk_validbcast_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_validbcast_FFY_RST,
      O => rx_input_memio_addrchk_validbcast
    );
  rx_input_memio_addrchk_n0051_SW0 : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_addrchk_bcast(3),
      ADR2 => rx_input_memio_addrchk_bcast(5),
      ADR3 => rx_input_memio_addrchk_bcast(4),
      O => rx_input_memio_addrchk_validbcast_FROM
    );
  rx_input_memio_addrchk_n0051_1603 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_bcast(1),
      ADR1 => rx_input_memio_addrchk_bcast(2),
      ADR2 => rx_input_memio_addrchk_bcast(0),
      ADR3 => rx_input_memio_addrchk_N70362,
      O => rx_input_memio_addrchk_n0051
    );
  rx_input_memio_addrchk_validbcast_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_validbcast_CEMUXNOT
    );
  rx_input_memio_addrchk_validbcast_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_validbcast_FROM,
      O => rx_input_memio_addrchk_N70362
    );
  mac_control_rxoferr_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(20),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(20)
    );
  mac_control_rxoferr_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(22),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(22)
    );
  mac_control_rxoferr_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(25),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(25)
    );
  mac_control_rxoferr_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(29),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(29)
    );
  mac_control_rxoferr_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(24),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(24)
    );
  mac_control_rxoferr_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(27),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(27)
    );
  mac_control_rxoferr_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(2),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(2)
    );
  mac_control_rxoferr_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(4),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(4)
    );
  mac_control_rxoferr_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(7),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(7)
    );
  mac_control_rxoferr_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(11),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(11)
    );
  mac_control_rxoferr_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(6),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(6)
    );
  mac_control_rxoferr_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(9),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(9)
    );
  mac_control_rxoferr_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(5),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(5)
    );
  rx_input_memio_bp_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(12),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_12_FFX_RST,
      O => rx_input_memio_bp(12)
    );
  rx_input_memio_bp_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_12_FFX_RST
    );
  rx_input_memio_bp_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(14),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_14_FFX_RST,
      O => rx_input_memio_bp(14)
    );
  rx_input_memio_bp_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_14_FFX_RST
    );
  mac_control_rxoferr_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(3),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(3)
    );
  mac_control_rxoferr_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_Madd_n0000_inst_lut2_16,
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(0)
    );
  mac_control_rxphyerr_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(10),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(10)
    );
  mac_control_rxphyerr_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(12),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(12)
    );
  mac_control_rxphyerr_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(19),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(19)
    );
  mac_control_rxphyerr_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(14),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(14)
    );
  mac_control_rxphyerr_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(17),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(17)
    );
  mac_control_rxphyerr_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(21),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(21)
    );
  mac_control_rxfifowerr_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(4),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(4)
    );
  mac_control_rxfifowerr_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(11),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(11)
    );
  mac_control_rxfifowerr_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(6),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(6)
    );
  mac_control_rxfifowerr_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(9),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(9)
    );
  mac_control_rxfifowerr_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(13),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(13)
    );
  mac_control_rxfifowerr_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(8),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(8)
    );
  mac_control_txfifowerr_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(2),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(2)
    );
  mac_control_txfifowerr_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(4),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(4)
    );
  mac_control_txfifowerr_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(7),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(7)
    );
  mac_control_txfifowerr_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(11),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(11)
    );
  mac_control_txfifowerr_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(6),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(6)
    );
  mac_control_txfifowerr_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(9),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(9)
    );
  mac_control_rxoferr_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(26),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(26)
    );
  mac_control_rxoferr_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(28),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(28)
    );
  mac_control_rxoferr_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(31),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(31)
    );
  mac_control_ledrx_cnt_156_1604 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_303,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_155_FFY_RST,
      O => mac_control_ledrx_cnt_156
    );
  mac_control_ledrx_cnt_155_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_155_FFY_RST
    );
  mac_control_rxoferr_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(30),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(30)
    );
  mac_control_ledrx_cnt_154_1605 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_301,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_154_FFY_RST,
      O => mac_control_ledrx_cnt_154
    );
  mac_control_ledrx_cnt_154_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_154_FFY_RST
    );
  mac_control_rxphyerr_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(1),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(1)
    );
  mac_control_rxphyerr_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_Madd_n0000_inst_lut2_16,
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(0)
    );
  mac_control_rxphyerr_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(7),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(7)
    );
  mac_control_rxphyerr_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(2),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(2)
    );
  mac_control_rxphyerr_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(5),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(5)
    );
  mac_control_rxphyerr_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(9),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(9)
    );
  mac_control_rxphyerr_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(22),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(22)
    );
  mac_control_rxphyerr_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(24),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(24)
    );
  mac_control_rxphyerr_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(31),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(31)
    );
  mac_control_rxphyerr_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(26),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(26)
    );
  mac_control_rxphyerr_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(29),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(29)
    );
  mac_control_rxfifowerr_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(1),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(1)
    );
  rx_fifocheck_diff_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_0_FFY_RST,
      O => rx_fifocheck_diff(1)
    );
  rx_fifocheck_diff_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_0_FFY_RST
    );
  rx_fifocheck_diff_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_4_FFY_RST,
      O => rx_fifocheck_diff(5)
    );
  rx_fifocheck_diff_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_4_FFY_RST
    );
  rx_fifocheck_diff_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_0_FFX_RST,
      O => rx_fifocheck_diff(0)
    );
  rx_fifocheck_diff_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_0_FFX_RST
    );
  rx_fifocheck_diff_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_2_FFY_RST,
      O => rx_fifocheck_diff(3)
    );
  rx_fifocheck_diff_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_2_FFY_RST
    );
  rx_output_bp_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(1),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_0_FFY_RST,
      O => rx_output_bp(1)
    );
  rx_output_bp_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_0_FFY_RST
    );
  rx_output_bp_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(3),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_2_FFY_RST,
      O => rx_output_bp(3)
    );
  rx_output_bp_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_2_FFY_RST
    );
  rx_output_bp_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(0),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_0_FFX_RST,
      O => rx_output_bp(0)
    );
  rx_output_bp_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_0_FFX_RST
    );
  rx_output_bp_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(7),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_6_FFY_RST,
      O => rx_output_bp(7)
    );
  rx_output_bp_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_6_FFY_RST
    );
  rx_output_bp_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(2),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_2_FFX_RST,
      O => rx_output_bp(2)
    );
  rx_output_bp_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_2_FFX_RST
    );
  rx_output_bp_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(5),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_4_FFY_RST,
      O => rx_output_bp(5)
    );
  rx_output_bp_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_4_FFY_RST
    );
  mac_control_ledrx_cnt_155_1606 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_302,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_155_FFX_RST,
      O => mac_control_ledrx_cnt_155
    );
  mac_control_ledrx_cnt_155_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_155_FFX_RST
    );
  mac_control_ledrx_cnt_158_1607 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_305,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_157_FFY_RST,
      O => mac_control_ledrx_cnt_158
    );
  mac_control_ledrx_cnt_157_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_157_FFY_RST
    );
  mac_control_ledrx_cnt_162_1608 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_309,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_161_FFY_RST,
      O => mac_control_ledrx_cnt_162
    );
  mac_control_ledrx_cnt_161_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_161_FFY_RST
    );
  mac_control_ledrx_cnt_157_1609 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_304,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_157_FFX_RST,
      O => mac_control_ledrx_cnt_157
    );
  mac_control_ledrx_cnt_157_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_157_FFX_RST
    );
  mac_control_ledrx_cnt_160_1610 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_307,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_159_FFY_RST,
      O => mac_control_ledrx_cnt_160
    );
  mac_control_ledrx_cnt_159_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_159_FFY_RST
    );
  mac_control_Mmux_n0016_Result_29_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_phyaddr(29),
      ADR1 => mac_control_n00851_1,
      ADR2 => mac_control_n0065,
      ADR3 => mac_control_rxphyerr_cntl(29),
      O => mac_control_CHOICE2273_FROM
    );
  mac_control_Mmux_n0016_Result_25_22 : X_LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      ADR0 => mac_control_rxphyerr_cntl(25),
      ADR1 => mac_control_n0065,
      ADR2 => mac_control_n00851_1,
      ADR3 => mac_control_phyaddr(25),
      O => mac_control_CHOICE2273_GROM
    );
  mac_control_CHOICE2273_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE2273_FROM,
      O => mac_control_CHOICE2273
    );
  mac_control_CHOICE2273_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2273_GROM,
      O => mac_control_CHOICE2204
    );
  rx_input_memio_crccomb_Mxor_CO_23_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_Mxor_CO_23_Xo(0),
      ADR1 => rx_input_memio_crcl(15),
      ADR2 => rx_input_memio_crcl(30),
      ADR3 => rx_input_memio_datal(1),
      O => rx_input_memio_crcl_23_FROM
    );
  rx_input_memio_n0048_23_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_23_Q,
      O => rx_input_memio_n0048_23_Q
    );
  rx_input_memio_crcl_23_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_23_FROM,
      O => rx_input_memio_crc_23_Q
    );
  mac_control_Mmux_n0016_Result_28_28 : X_LUT4
    generic map(
      INIT => X"ECA0"
    )
    port map (
      ADR0 => mac_control_n0066,
      ADR1 => mac_control_txf_cntl(28),
      ADR2 => mac_control_rxoferr_cntl(28),
      ADR3 => mac_control_n0061,
      O => mac_control_CHOICE2254_GROM
    );
  mac_control_CHOICE2254_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE2254_GROM,
      O => mac_control_CHOICE2254
    );
  rx_input_memio_addrchk_rxallfl_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_rxallfl_CEMUXNOT
    );
  rx_input_memio_cs_FFd16_In0 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_cs_FFd3,
      O => rx_input_memio_CHOICE1112_GROM
    );
  rx_input_memio_CHOICE1112_YUSED : X_BUF
    port map (
      I => rx_input_memio_CHOICE1112_GROM,
      O => rx_input_memio_CHOICE1112
    );
  tx_output_crc_loigc_Mxor_CO_29_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0124(0),
      ADR1 => tx_output_crc_loigc_n0124(1),
      ADR2 => tx_output_crcl(21),
      ADR3 => tx_output_crc_loigc_n0104(0),
      O => tx_output_crcl_29_FROM
    );
  tx_output_n0034_29_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_29_Q,
      O => tx_output_n0034_29_Q
    );
  tx_output_crcl_29_XUSED : X_BUF
    port map (
      I => tx_output_crcl_29_FROM,
      O => tx_output_crc_29_Q
    );
  rx_input_memio_crcll_11_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_11_CEMUXNOT
    );
  rx_input_memio_crcll_13_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_13_CEMUXNOT
    );
  rx_input_memio_crcll_21_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_21_CEMUXNOT
    );
  rx_input_memio_crcll_15_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_15_CEMUXNOT
    );
  rx_input_memio_crcll_31_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_31_CEMUXNOT
    );
  rx_input_memio_crcll_23_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_23_CEMUXNOT
    );
  rx_input_memio_crcll_17_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_17_CEMUXNOT
    );
  rx_input_memio_crcll_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_25_FFY_RST
    );
  rx_input_memio_crcll_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(24),
      CE => rx_input_memio_crcll_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_25_FFY_RST,
      O => rx_input_memio_crcll(24)
    );
  rx_input_memio_crcll_25_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_25_CEMUXNOT
    );
  rx_input_memio_crcll_27_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_27_CEMUXNOT
    );
  rx_input_memio_crcll_19_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_19_CEMUXNOT
    );
  rx_input_memio_crcll_29_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_crcll_29_CEMUXNOT
    );
  rx_input_memio_crccomb_Mxor_CO_24_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0118(1),
      ADR1 => rx_input_memio_crccomb_n0124(0),
      ADR2 => rx_input_memio_crccomb_n0122(0),
      ADR3 => rx_input_memio_crcl(16),
      O => rx_input_memio_crcl_24_FROM
    );
  rx_input_memio_n0048_24_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_24_Q,
      O => rx_input_memio_n0048_24_Q
    );
  rx_input_memio_crcl_24_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_24_FROM,
      O => rx_input_memio_crc_24_Q
    );
  rx_input_memio_crccomb_Mxor_CO_16_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0118(0),
      ADR1 => rx_input_memio_crcl(8),
      ADR2 => rx_input_memio_crccomb_n0115(0),
      ADR3 => rx_input_memio_crccomb_n0122(1),
      O => rx_input_memio_crcl_16_FROM
    );
  rx_input_memio_n0048_16_1 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_memio_crcrst,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_16_Q,
      O => rx_input_memio_n0048_16_1_O
    );
  rx_input_memio_crcl_16_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_16_FROM,
      O => rx_input_memio_crc_16_Q
    );
  mac_control_Ker531301 : X_LUT4
    generic map(
      INIT => X"0003"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_addr(4),
      ADR2 => mac_control_addr(1),
      ADR3 => mac_control_addr(2),
      O => mac_control_N53132_FROM
    );
  mac_control_n00591 : X_LUT4
    generic map(
      INIT => X"C000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_addr(3),
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_N53132,
      O => mac_control_N53132_GROM
    );
  mac_control_N53132_XUSED : X_BUF
    port map (
      I => mac_control_N53132_FROM,
      O => mac_control_N53132
    );
  mac_control_N53132_YUSED : X_BUF
    port map (
      I => mac_control_N53132_GROM,
      O => mac_control_n0059
    );
  mac_control_Ker532021 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_addr(0),
      ADR3 => mac_control_addr(1),
      O => mac_control_N53204_FROM
    );
  mac_control_n00621 : X_LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      ADR0 => mac_control_addr(2),
      ADR1 => mac_control_addr(3),
      ADR2 => mac_control_addr(4),
      ADR3 => mac_control_N53204,
      O => mac_control_N53204_GROM
    );
  mac_control_N53204_XUSED : X_BUF
    port map (
      I => mac_control_N53204_FROM,
      O => mac_control_N53204
    );
  mac_control_N53204_YUSED : X_BUF
    port map (
      I => mac_control_N53204_GROM,
      O => mac_control_n0062
    );
  mac_control_Ker531231 : X_LUT4
    generic map(
      INIT => X"0030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_addr(3),
      ADR2 => mac_control_addr(4),
      ADR3 => mac_control_addr(2),
      O => mac_control_N53125_FROM
    );
  mac_control_n00611 : X_LUT4
    generic map(
      INIT => X"4400"
    )
    port map (
      ADR0 => mac_control_addr(1),
      ADR1 => mac_control_addr(0),
      ADR2 => VCC,
      ADR3 => mac_control_N53125,
      O => mac_control_N53125_GROM
    );
  mac_control_N53125_XUSED : X_BUF
    port map (
      I => mac_control_N53125_FROM,
      O => mac_control_N53125
    );
  mac_control_N53125_YUSED : X_BUF
    port map (
      I => mac_control_N53125_GROM,
      O => mac_control_n0061
    );
  mac_control_Ker531161 : X_LUT4
    generic map(
      INIT => X"0088"
    )
    port map (
      ADR0 => mac_control_addr(2),
      ADR1 => mac_control_addr(4),
      ADR2 => VCC,
      ADR3 => mac_control_addr(3),
      O => mac_control_N53118_FROM
    );
  mac_control_n00671 : X_LUT4
    generic map(
      INIT => X"A000"
    )
    port map (
      ADR0 => mac_control_addr(0),
      ADR1 => VCC,
      ADR2 => mac_control_addr(1),
      ADR3 => mac_control_N53118,
      O => mac_control_N53118_GROM
    );
  mac_control_N53118_XUSED : X_BUF
    port map (
      I => mac_control_N53118_FROM,
      O => mac_control_N53118
    );
  mac_control_N53118_YUSED : X_BUF
    port map (
      I => mac_control_N53118_GROM,
      O => mac_control_n0067
    );
  mac_control_Ker531521 : X_LUT4
    generic map(
      INIT => X"0005"
    )
    port map (
      ADR0 => mac_control_bitcnt_109,
      ADR1 => VCC,
      ADR2 => mac_control_bitcnt_108,
      ADR3 => mac_control_bitcnt_107,
      O => mac_control_N53154_FROM
    );
  mac_control_n00111 : X_LUT4
    generic map(
      INIT => X"0050"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => mac_control_sclkdelta,
      ADR3 => mac_control_N53154,
      O => mac_control_N53154_GROM
    );
  mac_control_N53154_XUSED : X_BUF
    port map (
      I => mac_control_N53154_FROM,
      O => mac_control_N53154
    );
  mac_control_N53154_YUSED : X_BUF
    port map (
      I => mac_control_N53154_GROM,
      O => mac_control_n0011
    );
  mac_control_Ker531471 : X_LUT4
    generic map(
      INIT => X"8080"
    )
    port map (
      ADR0 => mac_control_sclkdeltal,
      ADR1 => mac_control_addr(7),
      ADR2 => mac_control_n0085,
      ADR3 => VCC,
      O => mac_control_PHY_status_phyaddrws_FROM
    );
  mac_control_PHY_status_n00151 : X_LUT4
    generic map(
      INIT => X"5550"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_cs_FFd1,
      ADR3 => mac_control_phyaddrw,
      O => mac_control_PHY_status_phyaddrws_GROM
    );
  mac_control_PHY_status_phyaddrws_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_phyaddrws_FROM,
      O => mac_control_phyaddrw
    );
  mac_control_PHY_status_phyaddrws_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_phyaddrws_GROM,
      O => mac_control_PHY_status_n00151_O
    );
  mac_control_PHY_status_phyaddrws_BYMUX : X_INV
    port map (
      I => mac_control_PHY_status_cs_FFd1,
      O => mac_control_PHY_status_phyaddrws_BYMUXNOT
    );
  mac_control_Ker531571 : X_LUT4
    generic map(
      INIT => X"4040"
    )
    port map (
      ADR0 => mac_control_addr(5),
      ADR1 => mac_control_n0086,
      ADR2 => mac_control_sclkdeltall,
      ADR3 => VCC,
      O => mac_control_dout_31_FROM
    );
  mac_control_Mmux_n0016_Result_31_85 : X_LUT4
    generic map(
      INIT => X"F222"
    )
    port map (
      ADR0 => mac_control_dout(30),
      ADR1 => mac_control_n0044,
      ADR2 => mac_control_N81176,
      ADR3 => mac_control_N53159,
      O => mac_control_n0016(31)
    );
  mac_control_dout_31_XUSED : X_BUF
    port map (
      I => mac_control_dout_31_FROM,
      O => mac_control_N53159
    );
  mac_control_Ker531921 : X_LUT4
    generic map(
      INIT => X"0008"
    )
    port map (
      ADR0 => mac_control_N53125,
      ADR1 => mac_control_sclkdeltal,
      ADR2 => mac_control_addr_0_1,
      ADR3 => mac_control_addr(1),
      O => mac_control_rxcrcerr_rst_FROM
    );
  mac_control_n00521 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_din(6),
      ADR3 => mac_control_N53194,
      O => mac_control_n0052
    );
  mac_control_rxcrcerr_rst_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_rst_CEMUXNOT
    );
  mac_control_rxcrcerr_rst_XUSED : X_BUF
    port map (
      I => mac_control_rxcrcerr_rst_FROM,
      O => mac_control_N53194
    );
  mac_control_PHY_status_MII_Interface_sout361 : X_LUT4
    generic map(
      INIT => X"0ACC"
    )
    port map (
      ADR0 => mac_control_PHY_status_din(5),
      ADR1 => mac_control_PHY_status_miiaddr(3),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(4),
      O => mac_control_PHY_status_MII_Interface_CHOICE963_FROM
    );
  mac_control_PHY_status_MII_Interface_sout365 : X_LUT4
    generic map(
      INIT => X"FF8A"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR1 => mac_control_PHY_status_din(1),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE963,
      O => mac_control_PHY_status_MII_Interface_CHOICE963_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE963_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE963_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE963
    );
  mac_control_PHY_status_MII_Interface_CHOICE963_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE963_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE964
    );
  rx_input_memio_crcequal_1611 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0059,
      CE => rx_input_memio_crcequal_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcequal_FFY_RST,
      O => rx_input_memio_crcequal
    );
  rx_input_memio_crcequal_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcequal_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_sout442 : X_LUT4
    generic map(
      INIT => X"5540"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR2 => mac_control_PHY_status_MII_Interface_CHOICE964,
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE977,
      O => mac_control_PHY_status_MII_Interface_CHOICE980_FROM
    );
  mac_control_PHY_status_MII_Interface_sout498_SW0 : X_LUT4
    generic map(
      INIT => X"F808"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR1 => mac_control_PHY_status_MII_Interface_CHOICE902,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(1),
      ADR3 => mac_control_PHY_status_MII_Interface_CHOICE980,
      O => mac_control_PHY_status_MII_Interface_CHOICE980_GROM
    );
  mac_control_PHY_status_MII_Interface_CHOICE980_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE980_FROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE980
    );
  mac_control_PHY_status_MII_Interface_CHOICE980_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_CHOICE980_GROM,
      O => mac_control_PHY_status_MII_Interface_N81411
    );
  tx_output_bpl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bpl_1_CEMUXNOT
    );
  tx_output_bpl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bpl_3_CEMUXNOT
    );
  tx_output_bpl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bpl_5_CEMUXNOT
    );
  tx_output_bpl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bpl_7_CEMUXNOT
    );
  tx_output_bpl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bpl_9_CEMUXNOT
    );
  macaddr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_13_FFY_RST
    );
  mac_control_MACADDR_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_13_FFY_RST,
      O => macaddr(12)
    );
  macaddr_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_21_FFY_RST
    );
  mac_control_MACADDR_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(20),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_21_FFY_RST,
      O => macaddr(20)
    );
  macaddr_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_31_FFY_RST
    );
  mac_control_MACADDR_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(30),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_31_FFY_RST,
      O => macaddr(30)
    );
  macaddr_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_23_FFY_RST
    );
  mac_control_MACADDR_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(22),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_23_FFY_RST,
      O => macaddr(22)
    );
  macaddr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_15_FFY_RST
    );
  mac_control_MACADDR_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_15_FFY_RST,
      O => macaddr(14)
    );
  macaddr_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_33_FFY_RST
    );
  mac_control_MACADDR_32 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(32),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_33_FFY_RST,
      O => macaddr(32)
    );
  macaddr_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_41_FFY_RST
    );
  mac_control_MACADDR_40 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(40),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_41_FFY_RST,
      O => macaddr(40)
    );
  mac_control_dout_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(4),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_4_FFY_RST,
      O => mac_control_dout(4)
    );
  mac_control_dout_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_4_FFY_RST
    );
  macaddr_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_25_FFY_RST
    );
  mac_control_MACADDR_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(24),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_25_FFY_RST,
      O => macaddr(24)
    );
  macaddr_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_17_FFY_RST
    );
  mac_control_MACADDR_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(16),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_17_FFY_RST,
      O => macaddr(16)
    );
  macaddr_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_27_FFY_RST
    );
  mac_control_MACADDR_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(26),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_27_FFY_RST,
      O => macaddr(26)
    );
  macaddr_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_35_FFY_RST
    );
  mac_control_MACADDR_34 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(34),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_35_FFY_RST,
      O => macaddr(34)
    );
  macaddr_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_19_FFY_RST
    );
  mac_control_MACADDR_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(18),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_19_FFY_RST,
      O => macaddr(18)
    );
  macaddr_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_29_FFY_RST
    );
  mac_control_MACADDR_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(28),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_29_FFY_RST,
      O => macaddr(28)
    );
  macaddr_37_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_37_FFY_RST
    );
  mac_control_MACADDR_36 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(36),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_37_FFY_RST,
      O => macaddr(36)
    );
  macaddr_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_45_FFY_RST
    );
  mac_control_MACADDR_44 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(44),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_45_FFY_RST,
      O => macaddr(44)
    );
  macaddr_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_39_FFY_RST
    );
  mac_control_MACADDR_38 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(38),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_39_FFY_RST,
      O => macaddr(38)
    );
  macaddr_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_47_FFY_RST
    );
  mac_control_MACADDR_46 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(46),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_47_FFY_RST,
      O => macaddr(46)
    );
  mac_control_PHY_status_addrl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_addrl_1_FFY_RST
    );
  mac_control_PHY_status_addrl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(0),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_addrl_1_FFY_RST,
      O => mac_control_PHY_status_addrl(0)
    );
  mac_control_PHY_status_addrl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_addrl_4_FFY_RST
    );
  mac_control_PHY_status_addrl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(4),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_addrl_4_FFY_RST,
      O => mac_control_PHY_status_addrl(4)
    );
  rx_input_memio_crcl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_25_FFY_RST
    );
  rx_input_memio_crcl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_25_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_25_FFY_RST,
      O => rx_input_memio_crcl(25)
    );
  rx_input_memio_crccomb_Mxor_CO_25_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(17),
      ADR1 => rx_input_memio_crccomb_n0124(1),
      ADR2 => rx_input_memio_crcl(26),
      ADR3 => rx_input_memio_datal(5),
      O => rx_input_memio_crcl_25_FROM
    );
  rx_input_memio_n0048_25_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_25_Q,
      O => rx_input_memio_n0048_25_Q
    );
  rx_input_memio_crcl_25_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_25_FROM,
      O => rx_input_memio_crc_25_Q
    );
  tx_output_cs_Out12_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd10,
      ADR1 => tx_output_cs_FFd14,
      ADR2 => tx_output_cs_FFd11,
      ADR3 => tx_output_cs_FFd13,
      O => tx_output_outsell_1_FROM
    );
  tx_output_cs_Out12 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => tx_output_cs_FFd15,
      ADR2 => tx_output_cs_FFd12,
      ADR3 => tx_output_N72900,
      O => tx_output_outsel_1_Q
    );
  tx_output_outsell_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_outsell_1_CEMUXNOT
    );
  tx_output_outsell_1_XUSED : X_BUF
    port map (
      I => tx_output_outsell_1_FROM,
      O => tx_output_N72900
    );
  rx_input_memio_crccomb_Mxor_CO_17_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(9),
      ADR1 => rx_input_memio_crccomb_n0122(0),
      ADR2 => rx_input_memio_crccomb_n0118(0),
      ADR3 => rx_input_memio_crccomb_n0104(0),
      O => rx_input_memio_crcl_17_FROM
    );
  rx_input_memio_n0048_17_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_17_Q,
      O => rx_input_memio_n0048_17_Q
    );
  rx_input_memio_crcl_17_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_17_FROM,
      O => rx_input_memio_crc_17_Q
    );
  tx_output_cs_Out13_SW0 : X_LUT4
    generic map(
      INIT => X"EEEE"
    )
    port map (
      ADR0 => tx_output_cs_FFd6_1,
      ADR1 => tx_output_cs_FFd5_1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => tx_output_outsell_0_FROM
    );
  tx_output_cs_Out13 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => tx_output_cs_FFd8,
      ADR1 => tx_output_cs_FFd4_1,
      ADR2 => tx_output_cs_FFd17,
      ADR3 => tx_output_N70101,
      O => tx_output_outsel_0_Q
    );
  tx_output_outsell_0_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_outsell_0_CEMUXNOT
    );
  tx_output_outsell_0_XUSED : X_BUF
    port map (
      I => tx_output_outsell_0_FROM,
      O => tx_output_N70101
    );
  memcontroller_oel_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => memcontroller_oel_CEMUXNOT
    );
  memcontroller_oel_BYMUX : X_INV
    port map (
      I => memcontroller_oe,
      O => memcontroller_oel_BYMUXNOT
    );
  rx_output_cs_FFd18_In_SW0 : X_LUT4
    generic map(
      INIT => X"3000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_output_nfl,
      ADR2 => rx_output_nf,
      ADR3 => rx_output_cs_FFd19,
      O => rx_output_cs_FFd18_FROM
    );
  rx_output_cs_FFd18_In_1612 : X_LUT4
    generic map(
      INIT => X"FFA2"
    )
    port map (
      ADR0 => rx_output_cs_FFd18,
      ADR1 => clken3,
      ADR2 => rx_output_n0017,
      ADR3 => rx_output_N71130,
      O => rx_output_cs_FFd18_In
    );
  rx_output_cs_FFd18_XUSED : X_BUF
    port map (
      I => rx_output_cs_FFd18_FROM,
      O => rx_output_N71130
    );
  tx_input_Ker35859107 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_input_CNT(15),
      ADR1 => tx_input_CNT(13),
      ADR2 => tx_input_CNT(12),
      ADR3 => tx_input_CNT(14),
      O => tx_input_CHOICE2029_FROM
    );
  tx_input_Ker3585926 : X_LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      ADR0 => tx_input_CNT(13),
      ADR1 => tx_input_CNT(14),
      ADR2 => tx_input_CNT(12),
      ADR3 => tx_input_CNT(15),
      O => tx_input_CHOICE2029_GROM
    );
  tx_input_CHOICE2029_XUSED : X_BUF
    port map (
      I => tx_input_CHOICE2029_FROM,
      O => tx_input_CHOICE2029
    );
  tx_input_CHOICE2029_YUSED : X_BUF
    port map (
      I => tx_input_CHOICE2029_GROM,
      O => tx_input_CHOICE1998
    );
  tx_input_Ker3585994 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_input_CNT(11),
      ADR1 => tx_input_CNT(8),
      ADR2 => tx_input_CNT(10),
      ADR3 => tx_input_CNT(9),
      O => tx_input_CHOICE2022_GROM
    );
  tx_input_CHOICE2022_YUSED : X_BUF
    port map (
      I => tx_input_CHOICE2022_GROM,
      O => tx_input_CHOICE2022
    );
  rx_output_fifo_nearfull_1613 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_wrcount(1),
      CE => rx_output_fifo_nearfull_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_nearfull_FFY_RST,
      O => rx_output_fifo_nearfull
    );
  rx_output_fifo_nearfull_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifo_nearfull_FFY_RST
    );
  mac_control_PHY_status_cs_Out51 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd6,
      ADR1 => VCC,
      ADR2 => mac_control_PHY_status_cs_FFd3,
      ADR3 => mac_control_PHY_status_cs_FFd8,
      O => mac_control_PHY_status_MII_Interface_cs_FFd6_FROM
    );
  mac_control_PHY_status_MII_Interface_cs_FFd6_In1 : X_LUT4
    generic map(
      INIT => X"CCFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_PHY_status_done,
      ADR2 => mac_control_PHY_status_MII_Interface_cs_FFd6,
      ADR3 => mac_control_PHY_status_start,
      O => mac_control_PHY_status_MII_Interface_cs_FFd6_In
    );
  mac_control_PHY_status_MII_Interface_cs_FFd6_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd6_FROM,
      O => mac_control_PHY_status_start
    );
  rx_input_memio_addrchk_cs_FFd6_In25_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => rx_input_memio_addrchk_cs_FFd7,
      ADR1 => rx_input_memio_addrchk_CHOICE1789,
      ADR2 => rx_input_memio_addrchk_cs_FFd2,
      ADR3 => rx_input_memio_addrchk_cs_FFd1,
      O => rx_input_memio_addrchk_cs_FFd6_FROM
    );
  rx_input_memio_addrchk_cs_FFd6_In25 : X_LUT4
    generic map(
      INIT => X"F444"
    )
    port map (
      ADR0 => rx_input_memio_brdy,
      ADR1 => rx_input_memio_addrchk_cs_FFd6,
      ADR2 => rx_input_memio_cs_FFd16_1,
      ADR3 => rx_input_memio_addrchk_N80994,
      O => rx_input_memio_addrchk_cs_FFd6_In
    );
  rx_input_memio_addrchk_cs_FFd6_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_cs_FFd6_FROM,
      O => rx_input_memio_addrchk_N80994
    );
  rx_input_memio_crccomb_Mxor_CO_26_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_datal(3),
      ADR1 => rx_input_memio_crcl(24),
      ADR2 => rx_input_memio_datal(7),
      ADR3 => rx_input_memio_crcl(28),
      O => rx_input_memio_crccomb_Mxor_CO_26_Xo_1_GROM
    );
  rx_input_memio_crccomb_Mxor_CO_26_Xo_1_YUSED : X_BUF
    port map (
      I => rx_input_memio_crccomb_Mxor_CO_26_Xo_1_GROM,
      O => rx_input_memio_crccomb_Mxor_CO_26_Xo(1)
    );
  rx_input_memio_crccomb_Mxor_CO_18_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(10),
      ADR1 => rx_input_memio_datal(0),
      ADR2 => rx_input_memio_crccomb_Mxor_CO_18_Xo(0),
      ADR3 => rx_input_memio_crcl(31),
      O => rx_input_memio_crcl_18_FROM
    );
  rx_input_memio_n0048_18_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_18_Q,
      O => rx_input_memio_n0048_18_Q
    );
  rx_input_memio_crcl_18_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_18_FROM,
      O => rx_input_memio_crc_18_Q
    );
  rx_input_memio_crccomb_Mxor_CO_26_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_Mxor_CO_26_Xo(1),
      ADR1 => rx_input_memio_crccomb_n0124(1),
      ADR2 => rx_input_memio_crccomb_n0104(0),
      ADR3 => rx_input_memio_crcl(18),
      O => rx_input_memio_crcl_26_FROM
    );
  rx_input_memio_n0048_26_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_26_Q,
      O => rx_input_memio_n0048_26_Q
    );
  rx_input_memio_crcl_26_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_26_FROM,
      O => rx_input_memio_crc_26_Q
    );
  memcontroller_clknum_1_BYMUX : X_INV
    port map (
      I => memcontroller_clknum_0_1,
      O => memcontroller_clknum_1_BYMUXNOT
    );
  txfbbp_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => txfbbp_1_CEMUXNOT
    );
  txfbbp_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => txfbbp_3_CEMUXNOT
    );
  txfbbp_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => txfbbp_5_CEMUXNOT
    );
  txfbbp_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => txfbbp_7_CEMUXNOT
    );
  txfbbp_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => txfbbp_9_CEMUXNOT
    );
  mac_control_dout_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(5),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_5_FFY_RST,
      O => mac_control_dout(5)
    );
  mac_control_dout_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_5_FFY_RST
    );
  tx_input_MA_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_18,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_3_FFY_RST,
      O => addr4ext(2)
    );
  addr4ext_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_3_FFY_RST
    );
  rx_input_fifo_control_d0_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_3_FFY_RST
    );
  rx_input_fifo_control_d0_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(2),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_3_FFY_RST,
      O => rx_input_fifo_control_d0(2)
    );
  rx_input_fifo_control_d0_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_5_FFY_RST
    );
  rx_input_fifo_control_d0_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(4),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_5_FFY_RST,
      O => rx_input_fifo_control_d0(4)
    );
  rx_input_fifo_control_d1_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_1_FFY_RST
    );
  rx_input_fifo_control_d1_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(0),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_1_FFY_RST,
      O => rx_input_fifo_control_d1(0)
    );
  rx_input_fifo_control_d1_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_3_FFY_RST
    );
  rx_input_fifo_control_d1_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(2),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_3_FFY_RST,
      O => rx_input_fifo_control_d1(2)
    );
  tx_input_MA_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_16,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_1_FFY_RST,
      O => addr4ext(0)
    );
  addr4ext_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_1_FFY_RST
    );
  rx_input_fifo_control_d0_9_LOGIC_ZERO_1614 : X_ZERO
    port map (
      O => rx_input_fifo_control_d0_9_LOGIC_ZERO
    );
  rx_input_fifo_control_dinl_9_rt_1615 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_dinl(9),
      ADR3 => VCC,
      O => rx_input_fifo_control_dinl_9_rt
    );
  tx_input_MA_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_17,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_1_FFX_RST,
      O => addr4ext(1)
    );
  addr4ext_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_1_FFX_RST
    );
  rx_input_fifo_control_d1_9_LOGIC_ZERO_1616 : X_ZERO
    port map (
      O => rx_input_fifo_control_d1_9_LOGIC_ZERO
    );
  rx_input_fifo_control_d0_9_rt_1617 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rx_input_fifo_control_d0(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_fifo_control_d0_9_rt
    );
  rx_input_fifo_control_d2_9_LOGIC_ZERO_1618 : X_ZERO
    port map (
      O => rx_input_fifo_control_d2_9_LOGIC_ZERO
    );
  rx_input_fifo_control_d1_9_rt_1619 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_fifo_control_d1(9),
      O => rx_input_fifo_control_d1_9_rt
    );
  rx_input_fifo_control_d3_9_LOGIC_ZERO_1620 : X_ZERO
    port map (
      O => rx_input_fifo_control_d3_9_LOGIC_ZERO
    );
  rx_input_fifo_control_d2_9_rt_1621 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_fifo_control_d2(9),
      ADR3 => VCC,
      O => rx_input_fifo_control_d2_9_rt
    );
  tx_input_MA_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_19,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_3_FFX_RST,
      O => addr4ext(3)
    );
  addr4ext_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_3_FFX_RST
    );
  rx_input_memio_crccomb_Mxor_CO_27_Xo_3_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crcl(19),
      ADR1 => rx_input_memio_crccomb_n0118(0),
      ADR2 => rx_input_memio_crccomb_Mxor_CO_9_Xo(0),
      ADR3 => rx_input_memio_crccomb_n0124(0),
      O => rx_input_memio_crcl_27_FROM
    );
  rx_input_memio_n0048_27_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_27_Q,
      O => rx_input_memio_n0048_27_Q
    );
  rx_input_memio_crcl_27_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_27_FROM,
      O => rx_input_memio_crc_27_Q
    );
  mac_control_rxoferr_cntl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_11_CEMUXNOT
    );
  mac_control_rxoferr_cntl_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_21_CEMUXNOT
    );
  mac_control_rxoferr_cntl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_13_CEMUXNOT
    );
  mac_control_rxoferr_cntl_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_31_CEMUXNOT
    );
  mac_control_rxoferr_cntl_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_23_CEMUXNOT
    );
  mac_control_rxoferr_cntl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_15_CEMUXNOT
    );
  mac_control_rxoferr_cntl_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_25_CEMUXNOT
    );
  mac_control_rxoferr_cntl_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_17_CEMUXNOT
    );
  mac_control_rxoferr_cntl_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_27_CEMUXNOT
    );
  tx_input_MA_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_21,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_5_FFX_RST,
      O => addr4ext(5)
    );
  addr4ext_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_5_FFX_RST
    );
  mac_control_rxoferr_cntl_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_19_CEMUXNOT
    );
  mac_control_rxoferr_cntl_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxoferr_cntl_29_CEMUXNOT
    );
  mac_control_PHY_status_miirw1 : X_LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd5,
      ADR1 => mac_control_PHY_status_cs_FFd6,
      ADR2 => mac_control_PHY_status_N43105,
      ADR3 => mac_control_PHY_status_rwl,
      O => mac_control_PHY_status_miirw_FROM
    );
  mac_control_PHY_status_MII_Interface_sout273_SW2 : X_LUT4
    generic map(
      INIT => X"3120"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR2 => mac_control_PHY_status_din(12),
      ADR3 => mac_control_PHY_status_miirw,
      O => mac_control_PHY_status_miirw_GROM
    );
  mac_control_PHY_status_miirw_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miirw_FROM,
      O => mac_control_PHY_status_miirw
    );
  mac_control_PHY_status_miirw_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miirw_GROM,
      O => mac_control_PHY_status_MII_Interface_N81407
    );
  rx_input_fifo_control_cell_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_cell_CEMUXNOT
    );
  rx_input_memio_crccomb_Mxor_CO_28_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0104(0),
      ADR1 => rx_input_memio_crccomb_n0118(1),
      ADR2 => rx_input_memio_crcl(20),
      ADR3 => rx_input_memio_crccomb_n0118(0),
      O => rx_input_memio_crcl_28_FROM
    );
  rx_input_memio_n0048_28_1 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rx_input_memio_crcrst,
      ADR3 => rx_input_memio_crc_28_Q,
      O => rx_input_memio_n0048_28_Q
    );
  rx_input_memio_crcl_28_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_28_FROM,
      O => rx_input_memio_crc_28_Q
    );
  mac_control_PHY_status_Ker431031 : X_LUT4
    generic map(
      INIT => X"FEFE"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd4,
      ADR1 => mac_control_PHY_status_cs_FFd2,
      ADR2 => mac_control_PHY_status_cs_FFd3,
      ADR3 => VCC,
      O => mac_control_PHY_status_N43105_FROM
    );
  mac_control_PHY_status_miiaddr_3_1 : X_LUT4
    generic map(
      INIT => X"FEFA"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd5,
      ADR1 => mac_control_PHY_status_addrl(3),
      ADR2 => mac_control_PHY_status_cs_FFd6,
      ADR3 => mac_control_PHY_status_N43105,
      O => mac_control_PHY_status_N43105_GROM
    );
  mac_control_PHY_status_N43105_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_N43105_FROM,
      O => mac_control_PHY_status_N43105
    );
  mac_control_PHY_status_N43105_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_N43105_GROM,
      O => mac_control_PHY_status_miiaddr(3)
    );
  mac_control_PHY_status_miiaddr_0_1 : X_LUT4
    generic map(
      INIT => X"FFFB"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd6,
      ADR1 => mac_control_PHY_status_N43105,
      ADR2 => mac_control_PHY_status_addrl(0),
      ADR3 => mac_control_PHY_status_cs_FFd5,
      O => mac_control_PHY_status_miiaddr_0_GROM
    );
  mac_control_PHY_status_miiaddr_0_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_0_GROM,
      O => mac_control_PHY_status_miiaddr(0)
    );
  mac_control_PHY_status_miiaddr_2_1 : X_LUT4
    generic map(
      INIT => X"FEFA"
    )
    port map (
      ADR0 => mac_control_PHY_status_cs_FFd5,
      ADR1 => mac_control_PHY_status_addrl(2),
      ADR2 => mac_control_PHY_status_cs_FFd6,
      ADR3 => mac_control_PHY_status_N43105,
      O => mac_control_PHY_status_miiaddr_2_FROM
    );
  mac_control_PHY_status_MII_Interface_sout178 : X_LUT4
    generic map(
      INIT => X"A280"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR2 => mac_control_PHY_status_din(4),
      ADR3 => mac_control_PHY_status_miiaddr(2),
      O => mac_control_PHY_status_miiaddr_2_GROM
    );
  mac_control_PHY_status_miiaddr_2_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_2_FROM,
      O => mac_control_PHY_status_miiaddr(2)
    );
  mac_control_PHY_status_miiaddr_2_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_2_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE921
    );
  mac_control_PHY_status_miiaddr_4_1 : X_LUT4
    generic map(
      INIT => X"0031"
    )
    port map (
      ADR0 => mac_control_PHY_status_N43105,
      ADR1 => mac_control_PHY_status_cs_FFd6,
      ADR2 => mac_control_PHY_status_addrl(4),
      ADR3 => mac_control_PHY_status_cs_FFd5,
      O => mac_control_PHY_status_miiaddr_4_FROM
    );
  mac_control_PHY_status_MII_Interface_sout222 : X_LUT4
    generic map(
      INIT => X"D580"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR1 => mac_control_PHY_status_din(6),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR3 => mac_control_PHY_status_miiaddr(4),
      O => mac_control_PHY_status_miiaddr_4_GROM
    );
  mac_control_PHY_status_miiaddr_4_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_4_FROM,
      O => mac_control_PHY_status_miiaddr(4)
    );
  mac_control_PHY_status_miiaddr_4_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_miiaddr_4_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE935
    );
  tx_input_MA_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_23,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_7_FFX_RST,
      O => addr4ext(7)
    );
  addr4ext_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_7_FFX_RST
    );
  tx_fifocheck_n000212 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(1),
      ADR1 => tx_fifocheck_diff(0),
      ADR2 => tx_fifocheck_diff(2),
      ADR3 => tx_fifocheck_diff(3),
      O => tx_fifocheck_CHOICE1918_GROM
    );
  tx_fifocheck_CHOICE1918_YUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1918_GROM,
      O => tx_fifocheck_CHOICE1918
    );
  rx_input_memio_crccomb_Mxor_CO_29_Xo_2_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rx_input_memio_crccomb_n0124(0),
      ADR1 => rx_input_memio_crccomb_n0104(0),
      ADR2 => rx_input_memio_crccomb_n0124(1),
      ADR3 => rx_input_memio_crcl(21),
      O => rx_input_memio_crcl_29_FROM
    );
  rx_input_memio_n0048_29_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_crcrst,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_crc_29_Q,
      O => rx_input_memio_n0048_29_Q
    );
  rx_input_memio_crcl_29_XUSED : X_BUF
    port map (
      I => rx_input_memio_crcl_29_FROM,
      O => rx_input_memio_crc_29_Q
    );
  tx_fifocheck_n000225 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(5),
      ADR1 => tx_fifocheck_diff(7),
      ADR2 => tx_fifocheck_diff(6),
      ADR3 => tx_fifocheck_diff(4),
      O => tx_fifocheck_CHOICE1925_GROM
    );
  tx_fifocheck_CHOICE1925_YUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1925_GROM,
      O => tx_fifocheck_CHOICE1925
    );
  tx_fifocheck_n000262 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(15),
      ADR1 => tx_fifocheck_diff(12),
      ADR2 => tx_fifocheck_diff(13),
      ADR3 => tx_fifocheck_diff(14),
      O => tx_fifocheck_CHOICE1940_GROM
    );
  tx_fifocheck_CHOICE1940_YUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1940_GROM,
      O => tx_fifocheck_CHOICE1940
    );
  tx_fifocheck_n000263 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => tx_fifocheck_CHOICE1933,
      ADR2 => VCC,
      ADR3 => tx_fifocheck_CHOICE1940,
      O => tx_fifocheck_CHOICE1941_FROM
    );
  tx_fifocheck_n000292 : X_LUT4
    generic map(
      INIT => X"F8F0"
    )
    port map (
      ADR0 => tx_fifocheck_CHOICE1925,
      ADR1 => tx_fifocheck_CHOICE1918,
      ADR2 => tx_fifocheck_n0003,
      ADR3 => tx_fifocheck_CHOICE1941,
      O => tx_fifocheck_CHOICE1941_GROM
    );
  tx_fifocheck_CHOICE1941_XUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1941_FROM,
      O => tx_fifocheck_CHOICE1941
    );
  tx_fifocheck_CHOICE1941_YUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1941_GROM,
      O => tx_fifocheck_n0002
    );
  tx_fifocheck_n000249 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_fifocheck_diff(11),
      ADR1 => tx_fifocheck_diff(9),
      ADR2 => tx_fifocheck_diff(10),
      ADR3 => tx_fifocheck_diff(8),
      O => tx_fifocheck_CHOICE1933_GROM
    );
  tx_fifocheck_CHOICE1933_YUSED : X_BUF
    port map (
      I => tx_fifocheck_CHOICE1933_GROM,
      O => tx_fifocheck_CHOICE1933
    );
  rx_input_fifo_control_celll_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_celll_CEMUXNOT
    );
  tx_input_MD_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(0),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_1_FFY_RST,
      O => d4(0)
    );
  d4_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_1_FFY_RST
    );
  mac_control_rxcrcerr_cntl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_11_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_21_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_13_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_23_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_15_CEMUXNOT
    );
  tx_input_MA_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_25,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_9_FFX_RST,
      O => addr4ext(9)
    );
  addr4ext_9_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_9_FFX_RST
    );
  mac_control_rxcrcerr_cntl_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_31_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_17_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_25_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_19_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_27_CEMUXNOT
    );
  mac_control_rxcrcerr_cntl_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxcrcerr_cntl_29_CEMUXNOT
    );
  rx_input_memio_cs_FFd3_In_SW0 : X_LUT4
    generic map(
      INIT => X"7777"
    )
    port map (
      ADR0 => rx_input_memio_crcequal,
      ADR1 => rx_input_memio_destok,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rx_input_memio_cs_FFd3_FROM
    );
  rx_input_memio_cs_FFd3_In_1622 : X_LUT4
    generic map(
      INIT => X"CCC8"
    )
    port map (
      ADR0 => rx_input_memio_fifofulll,
      ADR1 => rx_input_memio_cs_FFd5,
      ADR2 => rx_input_memio_endbyte(2),
      ADR3 => rx_input_memio_N70157,
      O => rx_input_memio_cs_FFd3_In
    );
  rx_input_memio_cs_FFd3_XUSED : X_BUF
    port map (
      I => rx_input_memio_cs_FFd3_FROM,
      O => rx_input_memio_N70157
    );
  mac_control_ledrx_rst_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_ledrx_rst_CEMUXNOT
    );
  rx_input_memio_addrchk_validmcast_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_validmcast_CEMUXNOT
    );
  mac_control_ledtx_rst_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_ledtx_rst_CEMUXNOT
    );
  tx_input_MD_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(1),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_1_FFX_RST,
      O => d4(1)
    );
  d4_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_1_FFX_RST
    );
  rx_input_memio_cs_FFd4_In_SW0 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => rx_input_memio_endbyte(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rx_input_memio_fifofulll,
      O => rx_input_memio_cs_FFd4_FROM
    );
  rx_input_memio_cs_FFd4_In_1623 : X_LUT4
    generic map(
      INIT => X"0080"
    )
    port map (
      ADR0 => rx_input_memio_crcequal,
      ADR1 => rx_input_memio_cs_FFd5,
      ADR2 => rx_input_memio_destok,
      ADR3 => rx_input_memio_N70191,
      O => rx_input_memio_cs_FFd4_In
    );
  rx_input_memio_cs_FFd4_XUSED : X_BUF
    port map (
      I => rx_input_memio_cs_FFd4_FROM,
      O => rx_input_memio_N70191
    );
  rxallf_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxallf_FFY_RST
    );
  mac_control_RXALLF : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lrxallf,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxallf_FFY_RST,
      O => rxallf
    );
  d4_23_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_23_FFY_RST
    );
  tx_input_MD_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(6),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_23_FFY_RST,
      O => d4(22)
    );
  d4_31_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_31_FFY_RST
    );
  tx_input_MD_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(14),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_31_FFY_RST,
      O => d4(30)
    );
  tx_input_MD_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(3),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_3_FFX_RST,
      O => d4(3)
    );
  d4_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_3_FFX_RST
    );
  d4_17_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_17_FFY_RST
    );
  tx_input_MD_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(0),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_17_FFY_RST,
      O => d4(16)
    );
  d4_29_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_29_FFY_RST
    );
  tx_input_MD_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(12),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_29_FFY_RST,
      O => d4(28)
    );
  rx_fifocheck_FIFOFULL : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfifofull_LOGIC_ONE,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_fifocheck_n0002,
      O => rxfifofull
    );
  rxfifofull_LOGIC_ONE_1624 : X_ONE
    port map (
      O => rxfifofull_LOGIC_ONE
    );
  mac_control_rxf_cntl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_1_CEMUXNOT
    );
  mac_control_rxf_cntl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_3_CEMUXNOT
    );
  mac_control_rxf_cntl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_5_CEMUXNOT
    );
  mac_control_rxf_cntl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_7_CEMUXNOT
    );
  mac_control_rxf_cntl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxf_cntl_9_CEMUXNOT
    );
  tx_input_MD_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(5),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_5_FFX_RST,
      O => d4(5)
    );
  d4_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_5_FFX_RST
    );
  rx_input_memio_addrchk_rxbcastl_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_rxbcastl_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_11_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_21_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_21_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_13_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_31_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_31_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_23_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_23_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_15_CEMUXNOT
    );
  tx_input_MD_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(8),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_9_FFY_RST,
      O => d4(8)
    );
  d4_9_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_9_FFY_RST
    );
  mac_control_rxphyerr_cntl_25_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_25_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_17_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_17_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_27_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_27_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_19_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_19_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_29_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_rxphyerr_cntl_29_CEMUXNOT
    );
  mac_control_rxphyerr_cntl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(0),
      CE => mac_control_rxphyerr_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_1_FFY_RST,
      O => mac_control_rxphyerr_cntl(0)
    );
  mac_control_rxphyerr_cntl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_1_FFY_RST
    );
  mac_control_rxphyerr_cntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(1),
      CE => mac_control_rxphyerr_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_1_FFX_RST,
      O => mac_control_rxphyerr_cntl(1)
    );
  mac_control_rxphyerr_cntl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_1_FFX_RST
    );
  mac_control_rxphyerr_cntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(4),
      CE => mac_control_rxphyerr_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_5_FFY_RST,
      O => mac_control_rxphyerr_cntl(4)
    );
  mac_control_rxphyerr_cntl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_5_FFY_RST
    );
  mac_control_n0032102 : X_LUT4
    generic map(
      INIT => X"0F0E"
    )
    port map (
      ADR0 => mac_control_CHOICE1404,
      ADR1 => mac_control_CHOICE1388,
      ADR2 => mac_control_phyrstcnt_141,
      ADR3 => mac_control_CHOICE1381,
      O => mac_control_CHOICE1407_FROM
    );
  mac_control_n0032126 : X_LUT4
    generic map(
      INIT => X"5550"
    )
    port map (
      ADR0 => RESET_IBUF,
      ADR1 => VCC,
      ADR2 => mac_control_N53144,
      ADR3 => mac_control_CHOICE1407,
      O => mac_control_CHOICE1407_GROM
    );
  mac_control_CHOICE1407_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1407_FROM,
      O => mac_control_CHOICE1407
    );
  mac_control_CHOICE1407_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1407_GROM,
      O => mac_control_n0032
    );
  tx_input_MD_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(7),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_7_FFX_RST,
      O => d4(7)
    );
  d4_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_7_FFX_RST
    );
  mac_control_n0034111 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_127,
      ADR1 => mac_control_phyrstcnt_128,
      ADR2 => mac_control_phyrstcnt_111,
      ADR3 => mac_control_phyrstcnt_129,
      O => mac_control_CHOICE1356_GROM
    );
  mac_control_CHOICE1356_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1356_GROM,
      O => mac_control_CHOICE1356
    );
  mac_control_n0034135 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_130,
      ADR1 => mac_control_phyrstcnt_122,
      ADR2 => mac_control_phyrstcnt_121,
      ADR3 => mac_control_phyrstcnt_131,
      O => mac_control_CHOICE1364_GROM
    );
  mac_control_CHOICE1364_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1364_GROM,
      O => mac_control_CHOICE1364
    );
  mac_control_n0034161 : X_LUT4
    generic map(
      INIT => X"4000"
    )
    port map (
      ADR0 => mac_control_N80971,
      ADR1 => mac_control_CHOICE1356,
      ADR2 => mac_control_CHOICE1371,
      ADR3 => mac_control_CHOICE1364,
      O => mac_control_CHOICE1373_FROM
    );
  mac_control_n0034194 : X_LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_141,
      ADR1 => mac_control_CHOICE1341,
      ADR2 => mac_control_CHOICE1326,
      ADR3 => mac_control_CHOICE1373,
      O => mac_control_CHOICE1373_GROM
    );
  mac_control_CHOICE1373_XUSED : X_BUF
    port map (
      I => mac_control_CHOICE1373_FROM,
      O => mac_control_CHOICE1373
    );
  mac_control_CHOICE1373_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1373_GROM,
      O => mac_control_n0034
    );
  mac_control_n0034148 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_124,
      ADR1 => mac_control_phyrstcnt_110,
      ADR2 => mac_control_phyrstcnt_123,
      ADR3 => mac_control_phyrstcnt_119,
      O => mac_control_CHOICE1371_GROM
    );
  mac_control_CHOICE1371_YUSED : X_BUF
    port map (
      I => mac_control_CHOICE1371_GROM,
      O => mac_control_CHOICE1371
    );
  mac_control_n003277_SW0 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_phyrstcnt_132,
      ADR1 => mac_control_phyrstcnt_131,
      ADR2 => mac_control_phyrstcnt_133,
      ADR3 => mac_control_phyrstcnt_134,
      O => mac_control_N80967_FROM
    );
  mac_control_n003277 : X_LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      ADR0 => mac_control_CHOICE1395,
      ADR1 => mac_control_CHOICE1399,
      ADR2 => mac_control_CHOICE1402,
      ADR3 => mac_control_N80967,
      O => mac_control_N80967_GROM
    );
  mac_control_N80967_XUSED : X_BUF
    port map (
      I => mac_control_N80967_FROM,
      O => mac_control_N80967
    );
  mac_control_N80967_YUSED : X_BUF
    port map (
      I => mac_control_N80967_GROM,
      O => mac_control_CHOICE1404
    );
  mac_control_n0086_1625 : X_LUT4
    generic map(
      INIT => X"0002"
    )
    port map (
      ADR0 => mac_control_bitcnt_107,
      ADR1 => mac_control_N69675,
      ADR2 => mac_control_bitcnt_106,
      ADR3 => mac_control_bitcnt_104,
      O => mac_control_n0086_FROM
    );
  mac_control_n00441 : X_LUT4
    generic map(
      INIT => X"F000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => mac_control_sclkdeltall,
      ADR3 => mac_control_n0086,
      O => mac_control_n0086_GROM
    );
  mac_control_n0086_XUSED : X_BUF
    port map (
      I => mac_control_n0086_FROM,
      O => mac_control_n0086
    );
  mac_control_n0086_YUSED : X_BUF
    port map (
      I => mac_control_n0086_GROM,
      O => mac_control_n0044
    );
  tx_input_MD_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(9),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_9_FFX_RST,
      O => d4(9)
    );
  d4_9_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_9_FFX_RST
    );
  rx_input_memio_addrchk_rxmcastl_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_rxmcastl_CEMUXNOT
    );
  rx_input_fifo_control_dinl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_dinl_1_CEMUXNOT
    );
  rx_input_fifo_control_dinl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_dinl_3_CEMUXNOT
    );
  rx_input_fifo_control_dinl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_dinl_5_CEMUXNOT
    );
  rx_input_fifo_control_dinl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_dinl_7_CEMUXNOT
    );
  rx_input_fifo_control_dinl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_dinl_9_CEMUXNOT
    );
  mac_control_n00851_1_1626 : X_LUT4
    generic map(
      INIT => X"00C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => mac_control_N53132,
      ADR2 => mac_control_addr(3),
      ADR3 => mac_control_addr(0),
      O => mac_control_n00851_1_FROM
    );
  mac_control_Mmux_n0016_Result_4_22 : X_LUT4
    generic map(
      INIT => X"EAC0"
    )
    port map (
      ADR0 => mac_control_phyaddr(4),
      ADR1 => mac_control_rxphyerr_cntl(4),
      ADR2 => mac_control_n0065,
      ADR3 => mac_control_n00851_1,
      O => mac_control_n00851_1_GROM
    );
  mac_control_n00851_1_XUSED : X_BUF
    port map (
      I => mac_control_n00851_1_FROM,
      O => mac_control_n00851_1
    );
  mac_control_n00851_1_YUSED : X_BUF
    port map (
      I => mac_control_n00851_1_GROM,
      O => mac_control_CHOICE2415
    );
  tx_fifocheck_fbbpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_11_FFX_RST,
      O => tx_fifocheck_fbbpl(11)
    );
  tx_fifocheck_fbbpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_11_FFX_RST
    );
  rx_input_memio_addrchk_rxucastl_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_rxucastl_CEMUXNOT
    );
  rx_input_memio_Ker425461 : X_LUT4
    generic map(
      INIT => X"0505"
    )
    port map (
      ADR0 => rx_input_endf,
      ADR1 => VCC,
      ADR2 => rx_input_invalid,
      ADR3 => VCC,
      O => rx_input_memio_addrchk_cs_FFd1_FROM
    );
  rx_input_memio_addrchk_cs_FFd1_In1 : X_LUT4
    generic map(
      INIT => X"4450"
    )
    port map (
      ADR0 => rx_input_memio_cs_FFd16_1,
      ADR1 => rx_input_memio_addrchk_cs_FFd2,
      ADR2 => rx_input_memio_addrchk_cs_FFd1,
      ADR3 => rx_input_memio_brdy,
      O => rx_input_memio_addrchk_cs_FFd1_In
    );
  rx_input_memio_addrchk_cs_FFd1_XUSED : X_BUF
    port map (
      I => rx_input_memio_addrchk_cs_FFd1_FROM,
      O => rx_input_memio_brdy
    );
  tx_fifocheck_fbbpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_13_FFX_RST,
      O => tx_fifocheck_fbbpl(13)
    );
  tx_fifocheck_fbbpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_13_FFX_RST
    );
  tx_fifocheck_fbbpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_15_FFX_RST,
      O => tx_fifocheck_fbbpl(15)
    );
  tx_fifocheck_fbbpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_15_FFX_RST
    );
  rxbp_11_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxbp_11_CEMUXNOT
    );
  rxbp_13_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxbp_13_CEMUXNOT
    );
  rxbp_15_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxbp_15_CEMUXNOT
    );
  rx_output_cs_FFd12_1627 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd13,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd12_FFX_RST,
      O => rx_output_cs_FFd12
    );
  rx_output_cs_FFd12_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd12_FFX_RST
    );
  rx_output_ceinl_1628 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cein,
      CE => rx_output_ceinl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_ceinl_FFX_RST,
      O => rx_output_ceinl
    );
  rx_output_ceinl_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_ceinl_FFX_RST
    );
  tx_output_n000774_SW0 : X_LUT4
    generic map(
      INIT => X"FEFF"
    )
    port map (
      ADR0 => tx_output_bcnt_41,
      ADR1 => tx_output_bcnt_39,
      ADR2 => tx_output_bcnt_40,
      ADR3 => tx_output_bcnt_38,
      O => tx_output_N80951_GROM
    );
  tx_output_N80951_YUSED : X_BUF
    port map (
      I => tx_output_N80951_GROM,
      O => tx_output_N80951
    );
  tx_output_bpl_11_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bpl_11_CEMUXNOT
    );
  tx_output_bpl_13_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bpl_13_CEMUXNOT
    );
  tx_output_bpl_15_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_bpl_15_CEMUXNOT
    );
  rx_output_cs_FFd14_1629 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd15,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd14_FFX_RST,
      O => rx_output_cs_FFd14
    );
  rx_output_cs_FFd14_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd14_FFX_RST
    );
  tx_output_cs_Out1145 : X_LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      ADR0 => tx_output_cs_FFd15,
      ADR1 => tx_output_cs_FFd17,
      ADR2 => tx_output_cs_FFd12,
      ADR3 => tx_output_cs_FFd14,
      O => tx_output_outsell_2_FROM
    );
  tx_output_cs_Out1157 : X_LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      ADR0 => tx_output_N81401,
      ADR1 => tx_output_cs_FFd16_1,
      ADR2 => tx_output_CHOICE1760,
      ADR3 => tx_output_CHOICE1767,
      O => tx_output_outsel_3_Q
    );
  tx_output_outsell_2_CEMUX : X_INV
    port map (
      I => RESET_IBUF_2,
      O => tx_output_outsell_2_CEMUXNOT
    );
  tx_output_outsell_2_XUSED : X_BUF
    port map (
      I => tx_output_outsell_2_FROM,
      O => tx_output_CHOICE1767
    );
  rx_input_memio_fifofulll_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rx_input_memio_fifofulll_CEMUXNOT
    );
  rx_output_nfl_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => rx_output_nfl_CEMUXNOT
    );
  mac_control_txf_cntl_1_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_1_CEMUXNOT
    );
  mac_control_txf_cntl_3_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_3_CEMUXNOT
    );
  mac_control_txf_cntl_5_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_5_CEMUXNOT
    );
  mac_control_txf_cntl_7_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_7_CEMUXNOT
    );
  mac_control_txf_cntl_9_CEMUX : X_INV
    port map (
      I => RESET_IBUF,
      O => mac_control_txf_cntl_9_CEMUXNOT
    );
  rx_output_cs_FFd16_1630 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd17,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd16_FFX_RST,
      O => rx_output_cs_FFd16
    );
  rx_output_cs_FFd16_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd16_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_sout142_SW0 : X_LUT4
    generic map(
      INIT => X"D0DF"
    )
    port map (
      ADR0 => mac_control_PHY_status_miiaddr(0),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(1),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(0),
      ADR3 => mac_control_PHY_status_miiaddr(1),
      O => mac_control_PHY_status_MII_Interface_N81171_FROM
    );
  mac_control_PHY_status_MII_Interface_sout142 : X_LUT4
    generic map(
      INIT => X"0020"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(3),
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR3 => mac_control_PHY_status_MII_Interface_N81171,
      O => mac_control_PHY_status_MII_Interface_N81171_GROM
    );
  mac_control_PHY_status_MII_Interface_N81171_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81171_FROM,
      O => mac_control_PHY_status_MII_Interface_N81171
    );
  mac_control_PHY_status_MII_Interface_N81171_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81171_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE915
    );
  tx_output_crc_loigc_Mxor_CO_3_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_loigc_n0122(0),
      ADR1 => tx_output_crc_loigc_n0118(1),
      ADR2 => tx_output_crc_loigc_n0124(0),
      ADR3 => tx_output_crc_loigc_n0124(1),
      O => tx_output_crcl_3_FROM
    );
  tx_output_n0034_3_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_3_Q,
      O => tx_output_n0034_3_Q
    );
  tx_output_crcl_3_XUSED : X_BUF
    port map (
      I => tx_output_crcl_3_FROM,
      O => tx_output_crc_3_Q
    );
  mac_control_PHY_status_MII_Interface_sout273_SW1 : X_LUT4
    generic map(
      INIT => X"AAEF"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_CHOICE935,
      ADR1 => mac_control_PHY_status_din(14),
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(4),
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(3),
      O => mac_control_PHY_status_MII_Interface_N81405_FROM
    );
  mac_control_PHY_status_MII_Interface_sout273 : X_LUT4
    generic map(
      INIT => X"FDA8"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_statecnt(1),
      ADR1 => mac_control_PHY_status_MII_Interface_CHOICE921,
      ADR2 => mac_control_PHY_status_MII_Interface_N81407,
      ADR3 => mac_control_PHY_status_MII_Interface_N81405,
      O => mac_control_PHY_status_MII_Interface_N81405_GROM
    );
  mac_control_PHY_status_MII_Interface_N81405_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81405_FROM,
      O => mac_control_PHY_status_MII_Interface_N81405
    );
  mac_control_PHY_status_MII_Interface_N81405_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81405_GROM,
      O => mac_control_PHY_status_MII_Interface_CHOICE944
    );
  mac_control_dout_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(6),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_6_FFY_RST,
      O => mac_control_dout(6)
    );
  mac_control_dout_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_6_FFY_RST
    );
  rx_input_fifo_RESET_1_1631 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => RESET_IBUF_2,
      ADR3 => VCC,
      O => rx_input_fifo_RESET_1_GROM
    );
  rx_input_fifo_RESET_1_YUSED : X_BUF
    port map (
      I => rx_input_fifo_RESET_1_GROM,
      O => rx_input_fifo_RESET_1
    );
  rxf_CEMUX : X_INV
    port map (
      I => rx_input_memio_RESET_1,
      O => rxf_CEMUXNOT
    );
  tx_output_crc_loigc_Mxor_CO_4_Xo_1_1 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => tx_output_crc_0_Q,
      ADR1 => tx_output_crc_loigc_n0118(1),
      ADR2 => tx_output_crc_loigc_n0115(0),
      ADR3 => tx_output_crc_loigc_n0124(1),
      O => tx_output_crcl_4_FROM
    );
  tx_output_n0034_4_1 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => tx_output_cs_FFd16_1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => tx_output_crc_4_Q,
      O => tx_output_n0034_4_1_O
    );
  tx_output_crcl_4_XUSED : X_BUF
    port map (
      I => tx_output_crcl_4_FROM,
      O => tx_output_crc_4_Q
    );
  mac_control_PHY_status_MII_Interface_sout485_SW0 : X_LUT4
    generic map(
      INIT => X"F200"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_CHOICE944,
      ADR1 => mac_control_PHY_status_MII_Interface_statecnt(2),
      ADR2 => mac_control_PHY_status_MII_Interface_CHOICE951,
      ADR3 => mac_control_PHY_status_MII_Interface_statecnt(0),
      O => mac_control_PHY_status_MII_Interface_N81167_FROM
    );
  mac_control_PHY_status_MII_Interface_sout498 : X_LUT4
    generic map(
      INIT => X"FFEF"
    )
    port map (
      ADR0 => mac_control_PHY_status_MII_Interface_N81411,
      ADR1 => mac_control_PHY_status_MII_Interface_CHOICE915,
      ADR2 => mac_control_PHY_status_MII_Interface_statecnt(5),
      ADR3 => mac_control_PHY_status_MII_Interface_N81167,
      O => mac_control_PHY_status_MII_Interface_N81167_GROM
    );
  mac_control_PHY_status_MII_Interface_N81167_XUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81167_FROM,
      O => mac_control_PHY_status_MII_Interface_N81167
    );
  mac_control_PHY_status_MII_Interface_N81167_YUSED : X_BUF
    port map (
      I => mac_control_PHY_status_MII_Interface_N81167_GROM,
      O => mac_control_PHY_status_MII_Interface_sout
    );
  mac_control_dout_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(7),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_7_FFY_RST,
      O => mac_control_dout(7)
    );
  mac_control_dout_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_7_FFY_RST
    );
  mac_control_rxf_cross_1632 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxf,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_rxf_cross_FFY_RST,
      O => mac_control_rxf_cross
    );
  mac_control_rxf_cross_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cross_FFY_RST
    );
  mac_control_rxphyerr_cntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(5),
      CE => mac_control_rxphyerr_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_5_FFX_RST,
      O => mac_control_rxphyerr_cntl(5)
    );
  mac_control_rxphyerr_cntl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_5_FFX_RST
    );
  mac_control_rxphyerr_cntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(7),
      CE => mac_control_rxphyerr_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_7_FFX_RST,
      O => mac_control_rxphyerr_cntl(7)
    );
  mac_control_rxphyerr_cntl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_7_FFX_RST
    );
  mac_control_rxphyerr_cntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(9),
      CE => mac_control_rxphyerr_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_9_FFX_RST,
      O => mac_control_rxphyerr_cntl(9)
    );
  mac_control_rxphyerr_cntl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_9_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(0),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_2_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(1)
    );
  mac_control_PHY_status_MII_Interface_dreg_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_2_FFY_RST
    );
  tx_output_cs_FFd14_1633 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd15,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd14_FFX_RST,
      O => tx_output_cs_FFd14
    );
  tx_output_cs_FFd14_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd14_FFX_RST
    );
  tx_output_data_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(2),
      CE => tx_output_data_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_2_FFY_RST,
      O => tx_output_data(2)
    );
  tx_output_data_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_2_FFY_RST
    );
  tx_output_data_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(3),
      CE => tx_output_data_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_3_FFY_RST,
      O => tx_output_data(3)
    );
  tx_output_data_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_3_FFY_RST
    );
  rx_input_memio_addrchk_cs_FFd7_1634 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd7_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_memio_addrchk_cs_FFd7_FFX_SET,
      RST => GND,
      O => rx_input_memio_addrchk_cs_FFd7
    );
  rx_input_memio_addrchk_cs_FFd7_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_memio_RESET_1,
      O => rx_input_memio_addrchk_cs_FFd7_FFX_SET
    );
  tx_output_data_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(6),
      CE => tx_output_data_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_6_FFY_RST,
      O => tx_output_data(6)
    );
  tx_output_data_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_6_FFY_RST
    );
  tx_fifocheck_FIFOFULL : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfifofull_LOGIC_ONE,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => tx_fifocheck_n0002,
      O => txfifofull
    );
  tx_output_data_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(7),
      CE => tx_output_data_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_7_FFY_RST,
      O => tx_output_data(7)
    );
  tx_output_data_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_7_FFY_RST
    );
  tx_output_bcntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_39,
      CE => tx_output_bcntl_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_2_FFY_RST,
      O => tx_output_bcntl(1)
    );
  tx_output_bcntl_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_2_FFY_RST
    );
  tx_output_bcntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_40,
      CE => tx_output_bcntl_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_2_FFX_RST,
      O => tx_output_bcntl(2)
    );
  tx_output_bcntl_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_2_FFX_RST
    );
  tx_output_bcntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_42,
      CE => tx_output_bcntl_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_4_FFX_RST,
      O => tx_output_bcntl(4)
    );
  tx_output_bcntl_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_4_FFX_RST
    );
  tx_output_bcntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_44,
      CE => tx_output_bcntl_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_6_FFX_RST,
      O => tx_output_bcntl(6)
    );
  tx_output_bcntl_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_6_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(11),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_11_FFX_RST,
      O => mac_control_PHY_status_dout(11)
    );
  mac_control_PHY_status_dout_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_11_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(13),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_13_FFX_RST,
      O => mac_control_PHY_status_dout(13)
    );
  mac_control_PHY_status_dout_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_13_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(15),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_15_FFX_RST,
      O => mac_control_PHY_status_dout(15)
    );
  mac_control_PHY_status_dout_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_15_FFX_RST
    );
  tx_output_ncrcbytel_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(1),
      CE => tx_output_ncrcbytel_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_1_FFY_RST,
      O => tx_output_ncrcbytel(1)
    );
  tx_output_ncrcbytel_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_1_FFY_RST
    );
  tx_output_ncrcbytel_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(2),
      CE => tx_output_ncrcbytel_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_2_FFY_RST,
      O => tx_output_ncrcbytel(2)
    );
  tx_output_ncrcbytel_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_2_FFY_RST
    );
  tx_output_ncrcbytel_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(3),
      CE => tx_output_ncrcbytel_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_3_FFY_RST,
      O => tx_output_ncrcbytel(3)
    );
  tx_output_ncrcbytel_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_3_FFY_RST
    );
  mac_control_dout_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(8),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_8_FFY_RST,
      O => mac_control_dout(8)
    );
  mac_control_dout_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_8_FFY_RST
    );
  tx_input_dh_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(0),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_1_FFY_RST,
      O => tx_input_dh(0)
    );
  tx_input_dh_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_1_FFY_RST
    );
  tx_input_dh_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(1),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_1_FFX_RST,
      O => tx_input_dh(1)
    );
  tx_input_dh_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_1_FFX_RST
    );
  tx_input_dh_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(3),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_3_FFX_RST,
      O => tx_input_dh(3)
    );
  tx_input_dh_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_3_FFX_RST
    );
  tx_input_dh_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(5),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_5_FFX_RST,
      O => tx_input_dh(5)
    );
  tx_input_dh_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_5_FFX_RST
    );
  tx_input_dh_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(6),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_7_FFY_RST,
      O => tx_input_dh(6)
    );
  tx_input_dh_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_7_FFY_RST
    );
  tx_input_dh_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(7),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_7_FFX_RST,
      O => tx_input_dh(7)
    );
  tx_input_dh_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_7_FFX_RST
    );
  tx_input_dl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(0),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_1_FFY_RST,
      O => tx_input_dl(0)
    );
  tx_input_dl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_1_FFY_RST
    );
  tx_input_dh_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(9),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_9_FFX_RST,
      O => tx_input_dh(9)
    );
  tx_input_dh_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_9_FFX_RST
    );
  tx_input_dl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(9),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_9_FFX_RST,
      O => tx_input_dl(9)
    );
  tx_input_dl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_9_FFX_RST
    );
  tx_input_bp_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_24,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_9_FFY_RST,
      O => txbp(8)
    );
  txbp_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_9_FFY_RST
    );
  tx_input_bp_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_25,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_9_FFX_RST,
      O => txbp(9)
    );
  txbp_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_9_FFX_RST
    );
  mac_control_lmacaddr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_1_FFY_RST,
      O => mac_control_lmacaddr(0)
    );
  mac_control_lmacaddr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_1_FFY_RST
    );
  mac_control_lmacaddr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_1_FFX_RST,
      O => mac_control_lmacaddr(1)
    );
  mac_control_lmacaddr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_1_FFX_RST
    );
  mac_control_lmacaddr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_3_FFX_RST,
      O => mac_control_lmacaddr(3)
    );
  mac_control_lmacaddr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_3_FFX_RST
    );
  mac_control_lmacaddr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_5_FFX_RST,
      O => mac_control_lmacaddr(5)
    );
  mac_control_lmacaddr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_5_FFX_RST
    );
  mac_control_lmacaddr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_7_FFX_RST,
      O => mac_control_lmacaddr(7)
    );
  mac_control_lmacaddr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_7_FFX_RST
    );
  rx_input_memio_BPOUT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_0_69,
      CE => rxbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_1_FFY_RST,
      O => rxbp(0)
    );
  rxbp_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_1_FFY_RST
    );
  mac_control_lmacaddr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_9_FFX_RST,
      O => mac_control_lmacaddr(9)
    );
  mac_control_lmacaddr_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_9_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(15),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_15_FFX_RST,
      O => mac_control_phydo(15)
    );
  mac_control_phydo_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_15_FFX_RST
    );
  tx_output_ltxen2_1635 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ltxen,
      CE => tx_output_ltxen3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ltxen3_FFY_RST,
      O => tx_output_ltxen2
    );
  tx_output_ltxen3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ltxen3_FFY_RST
    );
  tx_output_ltxen3_1636 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ltxen2,
      CE => tx_output_ltxen3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ltxen3_FFX_RST,
      O => tx_output_ltxen3
    );
  tx_output_ltxen3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ltxen3_FFX_RST
    );
  tx_input_cs_FFd1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd2,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_DONE_FFY_RST,
      O => tx_input_DONE
    );
  tx_input_DONE_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_DONE_FFY_RST
    );
  memcontroller_dnout_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_13_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_13_OFF_RST,
      O => memcontroller_dnout(13)
    );
  MD_13_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_13_OFF_RST
    );
  memcontroller_qn_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(22),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_22_IFF_RST,
      O => memcontroller_qn(22)
    );
  MD_22_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_22_IFF_RST
    );
  memcontroller_dnout_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_22_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_22_OFF_RST,
      O => memcontroller_dnout(22)
    );
  MD_22_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_22_OFF_RST
    );
  memcontroller_qn_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_14_IFF_RST,
      O => memcontroller_qn(14)
    );
  MD_14_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_14_IFF_RST
    );
  memcontroller_dnout_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_14_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_14_OFF_RST,
      O => memcontroller_dnout(14)
    );
  MD_14_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_14_OFF_RST
    );
  memcontroller_qn_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(30),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_30_IFF_RST,
      O => memcontroller_qn(30)
    );
  MD_30_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_30_IFF_RST
    );
  memcontroller_qn_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(23),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_23_IFF_RST,
      O => memcontroller_qn(23)
    );
  MD_23_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_23_IFF_RST
    );
  memcontroller_dnout_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_30_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_30_OFF_RST,
      O => memcontroller_dnout(30)
    );
  MD_30_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_30_OFF_RST
    );
  tx_input_dl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(1),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_1_FFX_RST,
      O => tx_input_dl(1)
    );
  tx_input_dl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_1_FFX_RST
    );
  tx_input_bp_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_17,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_1_FFX_RST,
      O => txbp(1)
    );
  txbp_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_1_FFX_RST
    );
  tx_input_dl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(3),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_3_FFX_RST,
      O => tx_input_dl(3)
    );
  tx_input_dl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_3_FFX_RST
    );
  tx_input_bp_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_18,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_3_FFY_RST,
      O => txbp(2)
    );
  txbp_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_3_FFY_RST
    );
  tx_input_bp_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_19,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_3_FFX_RST,
      O => txbp(3)
    );
  txbp_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_3_FFX_RST
    );
  tx_input_dl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(5),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_5_FFX_RST,
      O => tx_input_dl(5)
    );
  tx_input_dl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_5_FFX_RST
    );
  tx_input_bp_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_20,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_5_FFY_RST,
      O => txbp(4)
    );
  txbp_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_5_FFY_RST
    );
  tx_input_bp_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_21,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_5_FFX_RST,
      O => txbp(5)
    );
  txbp_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_5_FFX_RST
    );
  tx_input_dl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(7),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_7_FFX_RST,
      O => tx_input_dl(7)
    );
  tx_input_dl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_7_FFX_RST
    );
  tx_input_bp_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_22,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_7_FFY_RST,
      O => txbp(6)
    );
  txbp_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_7_FFY_RST
    );
  tx_input_bp_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_23,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_7_FFX_RST,
      O => txbp(7)
    );
  txbp_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_7_FFX_RST
    );
  mac_control_dout_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(0),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_0_FFY_RST,
      O => mac_control_dout(0)
    );
  mac_control_dout_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_0_FFY_RST
    );
  mac_control_rxf_cntl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(25),
      CE => mac_control_rxf_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_25_FFX_RST,
      O => mac_control_rxf_cntl(25)
    );
  mac_control_rxf_cntl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_25_FFX_RST
    );
  mac_control_rxf_cntl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(17),
      CE => mac_control_rxf_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_17_FFX_RST,
      O => mac_control_rxf_cntl(17)
    );
  mac_control_rxf_cntl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_17_FFX_RST
    );
  mac_control_rxf_cntl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(27),
      CE => mac_control_rxf_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_27_FFX_RST,
      O => mac_control_rxf_cntl(27)
    );
  mac_control_rxf_cntl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_27_FFX_RST
    );
  mac_control_rxf_cntl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(19),
      CE => mac_control_rxf_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_19_FFX_RST,
      O => mac_control_rxf_cntl(19)
    );
  mac_control_rxf_cntl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_19_FFX_RST
    );
  mac_control_rxf_cntl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(29),
      CE => mac_control_rxf_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_29_FFX_RST,
      O => mac_control_rxf_cntl(29)
    );
  mac_control_rxf_cntl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_29_FFX_RST
    );
  mac_control_dout_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(10),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_10_FFY_RST,
      O => mac_control_dout(10)
    );
  mac_control_dout_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_10_FFY_RST
    );
  rx_output_DOUT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_3_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_3_OFF_RST,
      O => rx_output_DOUT_3_OBUF
    );
  DOUT_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_3_OFF_RST
    );
  rx_output_DOUT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_4_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_4_OFF_RST,
      O => rx_output_DOUT_4_OBUF
    );
  DOUT_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_4_OFF_RST
    );
  rx_output_DOUT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_5_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_5_OFF_RST,
      O => rx_output_DOUT_5_OBUF
    );
  DOUT_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_5_OFF_RST
    );
  rx_output_DOUT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_6_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_6_OFF_RST,
      O => rx_output_DOUT_6_OBUF
    );
  DOUT_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_6_OFF_RST
    );
  rx_output_DOUT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_7_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_7_OFF_RST,
      O => rx_output_DOUT_7_OBUF
    );
  DOUT_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_7_OFF_RST
    );
  tx_output_outselll_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_outsell(1),
      CE => tx_output_outselll_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outselll_1_FFX_RST,
      O => tx_output_outselll(1)
    );
  tx_output_outselll_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outselll_1_FFX_RST
    );
  tx_output_outselll_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => tx_output_outsell(0),
      CE => tx_output_outselll_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => tx_output_outselll_1_FFY_SET,
      RST => GND,
      O => tx_output_outselll(0)
    );
  tx_output_outselll_1_FFY_SETOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outselll_1_FFY_SET
    );
  tx_output_outselll_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_outsell(3),
      CE => tx_output_outselll_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outselll_3_FFX_RST,
      O => tx_output_outselll(3)
    );
  tx_output_outselll_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outselll_3_FFX_RST
    );
  mac_control_txf_cntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(10),
      CE => mac_control_txf_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_11_FFY_RST,
      O => mac_control_txf_cntl(10)
    );
  mac_control_txf_cntl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_11_FFY_RST
    );
  mac_control_txf_cntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(11),
      CE => mac_control_txf_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_11_FFX_RST,
      O => mac_control_txf_cntl(11)
    );
  mac_control_txf_cntl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_11_FFX_RST
    );
  mac_control_txf_cntl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(21),
      CE => mac_control_txf_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_21_FFX_RST,
      O => mac_control_txf_cntl(21)
    );
  mac_control_txf_cntl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_21_FFX_RST
    );
  mac_control_txf_cntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(13),
      CE => mac_control_txf_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_13_FFX_RST,
      O => mac_control_txf_cntl(13)
    );
  mac_control_txf_cntl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_13_FFX_RST
    );
  mac_control_rxf_cntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(11),
      CE => mac_control_rxf_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_11_FFX_RST,
      O => mac_control_rxf_cntl(11)
    );
  mac_control_rxf_cntl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_11_FFX_RST
    );
  mac_control_rxf_cntl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(21),
      CE => mac_control_rxf_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_21_FFX_RST,
      O => mac_control_rxf_cntl(21)
    );
  mac_control_rxf_cntl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_21_FFX_RST
    );
  mac_control_rxf_cntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(13),
      CE => mac_control_rxf_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_13_FFX_RST,
      O => mac_control_rxf_cntl(13)
    );
  mac_control_rxf_cntl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_13_FFX_RST
    );
  mac_control_rxf_cntl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(31),
      CE => mac_control_rxf_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_31_FFX_RST,
      O => mac_control_rxf_cntl(31)
    );
  mac_control_rxf_cntl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_31_FFX_RST
    );
  mac_control_rxf_cntl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(23),
      CE => mac_control_rxf_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_23_FFX_RST,
      O => mac_control_rxf_cntl(23)
    );
  mac_control_rxf_cntl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_23_FFX_RST
    );
  mac_control_rxf_cntl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(24),
      CE => mac_control_rxf_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_25_FFY_RST,
      O => mac_control_rxf_cntl(24)
    );
  mac_control_rxf_cntl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_25_FFY_RST
    );
  mac_control_rxf_cntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(15),
      CE => mac_control_rxf_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_15_FFX_RST,
      O => mac_control_rxf_cntl(15)
    );
  mac_control_rxf_cntl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_15_FFX_RST
    );
  rx_output_fifo_BU372 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1603_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1603
    );
  rx_output_fifo_N1603_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1603_FFX_SET
    );
  rx_output_fifo_BU364 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N7,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1607_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1607
    );
  rx_output_fifo_N1607_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1607_FFX_SET
    );
  mac_control_PHY_status_PHYSTAT_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(9),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_25_FFX_RST,
      O => mac_control_phystat(25)
    );
  mac_control_phystat_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_25_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(1),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_17_FFX_RST,
      O => mac_control_phystat(17)
    );
  mac_control_phystat_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_17_FFX_RST
    );
  memcontroller_Q3_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(31),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_31_FFX_RST,
      O => q3(31)
    );
  q3_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_31_FFX_RST
    );
  memcontroller_Q3_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(14),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_15_FFY_RST,
      O => q3(14)
    );
  q3_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_15_FFY_RST
    );
  memcontroller_Q3_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(15),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_15_FFX_RST,
      O => q3(15)
    );
  q3_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_15_FFX_RST
    );
  rx_output_denl_1637 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_CHOICE880,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => GSR,
      SSET => rx_output_CHOICE876,
      SRST => rx_output_denl_LOGIC_ZERO,
      O => rx_output_denl
    );
  rx_input_memio_addrchk_mcast_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmcast(0),
      CE => rx_input_memio_addrchk_mcast_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_mcast_0_FFY_RST,
      O => rx_input_memio_addrchk_mcast(0)
    );
  rx_input_memio_addrchk_mcast_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_mcast_0_FFY_RST
    );
  tx_output_ncrcbytel_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(0),
      CE => tx_output_ncrcbytel_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_0_FFY_RST,
      O => tx_output_ncrcbytel(0)
    );
  tx_output_ncrcbytel_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_0_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(10),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_11_FFY_RST,
      O => mac_control_PHY_status_dout(10)
    );
  mac_control_PHY_status_dout_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_11_FFY_RST
    );
  tx_output_addr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(4),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_4_FFX_RST,
      O => addr2ext(4)
    );
  addr2ext_4_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_4_FFX_RST
    );
  tx_output_addr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(6),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_6_FFX_RST,
      O => addr2ext(6)
    );
  addr2ext_6_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_6_FFX_RST
    );
  tx_output_addr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(9),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_8_FFY_RST,
      O => addr2ext(9)
    );
  addr2ext_8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_8_FFY_RST
    );
  tx_output_addr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(11),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_10_FFY_RST,
      O => addr2ext(11)
    );
  addr2ext_10_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_10_FFY_RST
    );
  tx_output_addr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(13),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_12_FFY_RST,
      O => addr2ext(13)
    );
  addr2ext_12_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_12_FFY_RST
    );
  tx_output_addr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(14),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_14_FFX_RST,
      O => addr2ext(14)
    );
  addr2ext_14_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_14_FFX_RST
    );
  rx_input_memio_bcnt_87_1638 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_236,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_87_FFX_RST,
      O => rx_input_memio_bcnt_87
    );
  rx_input_memio_bcnt_87_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_87_FFX_RST
    );
  rx_input_memio_bcnt_90_1639 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_239,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_89_FFY_RST,
      O => rx_input_memio_bcnt_90
    );
  rx_input_memio_bcnt_89_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_89_FFY_RST
    );
  rx_input_memio_bcnt_92_1640 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_241,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_91_FFY_RST,
      O => rx_input_memio_bcnt_92
    );
  rx_input_memio_bcnt_91_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_91_FFY_RST
    );
  tx_output_data_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(1),
      CE => tx_output_data_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_1_FFY_RST,
      O => tx_output_data(1)
    );
  tx_output_data_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_1_FFY_RST
    );
  rx_input_memio_addrchk_cs_FFd2_1641 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd2_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd2_FFX_RST,
      O => rx_input_memio_addrchk_cs_FFd2
    );
  rx_input_memio_addrchk_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd2_FFX_RST
    );
  tx_fifocheck_fbbpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_3_FFX_RST,
      O => tx_fifocheck_fbbpl(3)
    );
  tx_fifocheck_fbbpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_3_FFX_RST
    );
  tx_fifocheck_fbbpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_5_FFX_RST,
      O => tx_fifocheck_fbbpl(5)
    );
  tx_fifocheck_fbbpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_5_FFX_RST
    );
  tx_fifocheck_fbbpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_7_FFY_RST,
      O => tx_fifocheck_fbbpl(6)
    );
  tx_fifocheck_fbbpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_7_FFY_RST
    );
  tx_fifocheck_fbbpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_7_FFX_RST,
      O => tx_fifocheck_fbbpl(7)
    );
  tx_fifocheck_fbbpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_7_FFX_RST
    );
  tx_fifocheck_fbbpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_9_FFX_RST,
      O => tx_fifocheck_fbbpl(9)
    );
  tx_fifocheck_fbbpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_9_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(11),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_11_FFX_RST,
      O => mac_control_phydo(11)
    );
  mac_control_phydo_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_11_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(12),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_13_FFY_RST,
      O => mac_control_phydo(12)
    );
  mac_control_phydo_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_13_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(13),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_13_FFX_RST,
      O => mac_control_phydo(13)
    );
  mac_control_phydo_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_13_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(14),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_15_FFY_RST,
      O => mac_control_phydo(14)
    );
  mac_control_phydo_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_15_FFY_RST
    );
  mac_control_RXUCAST : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lrxucast,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxucast_FFY_RST,
      O => rxucast
    );
  rxucast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxucast_FFY_RST
    );
  mac_control_dout_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(11),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_11_FFY_RST,
      O => mac_control_dout(11)
    );
  mac_control_dout_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_11_FFY_RST
    );
  tx_output_crcl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_12_1_O,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_12_FFX_RST,
      O => tx_output_crcl(12)
    );
  tx_output_crcl_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_12_FFX_RST
    );
  tx_output_crcsell_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd2,
      CE => tx_output_crcsell_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcsell_0_FFY_RST,
      O => tx_output_crcsell(1)
    );
  tx_output_crcsell_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcsell_0_FFY_RST
    );
  mac_control_rxoferr_cntl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(0),
      CE => mac_control_rxoferr_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_1_FFY_RST,
      O => mac_control_rxoferr_cntl(0)
    );
  mac_control_rxoferr_cntl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_1_FFY_RST
    );
  tx_output_crcsell_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => tx_output_crcsel(0),
      CE => tx_output_crcsell_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => tx_output_crcsell_0_FFX_SET,
      RST => GND,
      O => tx_output_crcsell(0)
    );
  tx_output_crcsell_0_FFX_SETOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcsell_0_FFX_SET
    );
  rx_input_memio_addrchk_bcast_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(4),
      CE => rx_input_memio_addrchk_bcast_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_4_FFY_RST,
      O => rx_input_memio_addrchk_bcast(4)
    );
  rx_input_memio_addrchk_bcast_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_4_FFY_RST
    );
  rx_input_memio_addrchk_bcast_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(1),
      CE => rx_input_memio_addrchk_bcast_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_1_FFY_RST,
      O => rx_input_memio_addrchk_bcast(1)
    );
  rx_input_memio_addrchk_bcast_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_1_FFY_RST
    );
  rx_output_ldouten2_1642 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_denll,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_output_invalid,
      O => rx_output_ldouten2
    );
  tx_output_cs_FFd15_1643 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd16_1,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd15_FFY_RST,
      O => tx_output_cs_FFd15
    );
  tx_output_cs_FFd15_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd15_FFY_RST
    );
  tx_output_cs_FFd12_1644 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd13,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd12_FFX_RST,
      O => tx_output_cs_FFd12
    );
  tx_output_cs_FFd12_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd12_FFX_RST
    );
  tx_output_cs_FFd13_1645 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd14,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd14_FFY_RST,
      O => tx_output_cs_FFd13
    );
  tx_output_cs_FFd14_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd14_FFY_RST
    );
  tx_output_ncrcbytel_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(4),
      CE => tx_output_ncrcbytel_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_4_FFY_RST,
      O => tx_output_ncrcbytel(4)
    );
  tx_output_ncrcbytel_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_4_FFY_RST
    );
  tx_output_ncrcbytel_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(5),
      CE => tx_output_ncrcbytel_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_5_FFY_RST,
      O => tx_output_ncrcbytel(5)
    );
  tx_output_ncrcbytel_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_5_FFY_RST
    );
  tx_output_ncrcbytel_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(6),
      CE => tx_output_ncrcbytel_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_6_FFY_RST,
      O => tx_output_ncrcbytel(6)
    );
  tx_output_ncrcbytel_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_6_FFY_RST
    );
  tx_output_ncrcbytel_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ncrcbyte(7),
      CE => tx_output_ncrcbytel_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_ncrcbytel_7_FFY_RST,
      O => tx_output_ncrcbytel(7)
    );
  tx_output_ncrcbytel_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_ncrcbytel_7_FFY_RST
    );
  mac_control_RXMCAST : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lrxmcast,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxmcast_FFY_RST,
      O => rxmcast
    );
  rxmcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxmcast_FFY_RST
    );
  mac_control_txfifowerr_cntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(11),
      CE => mac_control_txfifowerr_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_11_FFX_RST,
      O => mac_control_txfifowerr_cntl(11)
    );
  mac_control_txfifowerr_cntl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_11_FFX_RST
    );
  mac_control_txfifowerr_cntl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(21),
      CE => mac_control_txfifowerr_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_21_FFX_RST,
      O => mac_control_txfifowerr_cntl(21)
    );
  mac_control_txfifowerr_cntl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_21_FFX_RST
    );
  mac_control_txfifowerr_cntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(13),
      CE => mac_control_txfifowerr_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_13_FFX_RST,
      O => mac_control_txfifowerr_cntl(13)
    );
  mac_control_txfifowerr_cntl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_13_FFX_RST
    );
  mac_control_txfifowerr_cntl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(31),
      CE => mac_control_txfifowerr_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_31_FFX_RST,
      O => mac_control_txfifowerr_cntl(31)
    );
  mac_control_txfifowerr_cntl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_31_FFX_RST
    );
  mac_control_txfifowerr_cntl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(23),
      CE => mac_control_txfifowerr_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_23_FFX_RST,
      O => mac_control_txfifowerr_cntl(23)
    );
  mac_control_txfifowerr_cntl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_23_FFX_RST
    );
  mac_control_txfifowerr_cntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(15),
      CE => mac_control_txfifowerr_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_15_FFX_RST,
      O => mac_control_txfifowerr_cntl(15)
    );
  mac_control_txfifowerr_cntl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_15_FFX_RST
    );
  mac_control_txfifowerr_cntl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(24),
      CE => mac_control_txfifowerr_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_25_FFY_RST,
      O => mac_control_txfifowerr_cntl(24)
    );
  mac_control_txfifowerr_cntl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_25_FFY_RST
    );
  mac_control_txfifowerr_cntl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(25),
      CE => mac_control_txfifowerr_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_25_FFX_RST,
      O => mac_control_txfifowerr_cntl(25)
    );
  mac_control_txfifowerr_cntl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_25_FFX_RST
    );
  mac_control_txfifowerr_cntl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(17),
      CE => mac_control_txfifowerr_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_17_FFX_RST,
      O => mac_control_txfifowerr_cntl(17)
    );
  mac_control_txfifowerr_cntl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_17_FFX_RST
    );
  mac_control_txfifowerr_cntl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(27),
      CE => mac_control_txfifowerr_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_27_FFX_RST,
      O => mac_control_txfifowerr_cntl(27)
    );
  mac_control_txfifowerr_cntl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_27_FFX_RST
    );
  mac_control_txfifowerr_cntl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(19),
      CE => mac_control_txfifowerr_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_19_FFX_RST,
      O => mac_control_txfifowerr_cntl(19)
    );
  mac_control_txfifowerr_cntl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_19_FFX_RST
    );
  mac_control_txfifowerr_cntl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(29),
      CE => mac_control_txfifowerr_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_29_FFX_RST,
      O => mac_control_txfifowerr_cntl(29)
    );
  mac_control_txfifowerr_cntl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_29_FFX_RST
    );
  tx_fifocheck_fbbpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_1_FFY_RST,
      O => tx_fifocheck_fbbpl(0)
    );
  tx_fifocheck_fbbpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_1_FFY_RST
    );
  tx_fifocheck_fbbpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txfbbp(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_fbbpl_1_FFX_RST,
      O => tx_fifocheck_fbbpl(1)
    );
  tx_fifocheck_fbbpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_fbbpl_1_FFX_RST
    );
  rx_input_memio_cs_FFd7_1646 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd13,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd8_FFY_RST,
      O => rx_input_memio_cs_FFd7
    );
  rx_input_memio_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd8_FFY_RST
    );
  rx_input_memio_cs_FFd8_1647 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd8_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd8_FFX_RST,
      O => rx_input_memio_cs_FFd8
    );
  rx_input_memio_cs_FFd8_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd8_FFX_RST
    );
  mac_control_bitcnt_109_1648 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_256,
      CE => mac_control_n0015,
      CLK => clksl,
      SET => GND,
      RST => mac_control_bitcnt_109_FFX_RST,
      O => mac_control_bitcnt_109
    );
  mac_control_bitcnt_109_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_109_FFX_RST
    );
  tx_output_data_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(4),
      CE => tx_output_data_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_4_FFY_RST,
      O => tx_output_data(4)
    );
  tx_output_data_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_4_FFY_RST
    );
  tx_output_bcntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_49,
      CE => tx_output_bcntl_12_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_12_FFY_RST,
      O => tx_output_bcntl(11)
    );
  tx_output_bcntl_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_12_FFY_RST
    );
  tx_output_bcntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_50,
      CE => tx_output_bcntl_12_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_12_FFX_RST,
      O => tx_output_bcntl(12)
    );
  tx_output_bcntl_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_12_FFX_RST
    );
  rx_input_memio_addrchk_cs_FFd5_1649 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd5_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd5_FFX_RST,
      O => rx_input_memio_addrchk_cs_FFd5
    );
  rx_input_memio_addrchk_cs_FFd5_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd5_FFX_RST
    );
  rx_input_memio_addrchk_bcast_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(3),
      CE => rx_input_memio_addrchk_bcast_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_3_FFY_RST,
      O => rx_input_memio_addrchk_bcast(3)
    );
  rx_input_memio_addrchk_bcast_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_3_FFY_RST
    );
  rx_input_memio_addrchk_bcast_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(0),
      CE => rx_input_memio_addrchk_bcast_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_0_FFY_RST,
      O => rx_input_memio_addrchk_bcast(0)
    );
  rx_input_memio_addrchk_bcast_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_0_FFY_RST
    );
  rx_input_memio_addrchk_bcast_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(5),
      CE => rx_input_memio_addrchk_bcast_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_5_FFY_RST,
      O => rx_input_memio_addrchk_bcast(5)
    );
  rx_input_memio_addrchk_bcast_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_5_FFY_RST
    );
  rx_input_memio_addrchk_bcast_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lbcast(2),
      CE => rx_input_memio_addrchk_bcast_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_bcast_2_FFY_RST,
      O => rx_input_memio_addrchk_bcast(2)
    );
  rx_input_memio_addrchk_bcast_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_bcast_2_FFY_RST
    );
  mac_control_dout_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(13),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_13_FFY_RST,
      O => mac_control_dout(13)
    );
  mac_control_dout_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_13_FFY_RST
    );
  mac_control_Mshreg_scslll_103_1650 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_Mshreg_scslll_net187,
      CE => mac_control_Mshreg_scslll_103_CEMUXNOT,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_Mshreg_scslll_103_FFY_RST,
      O => mac_control_Mshreg_scslll_103
    );
  mac_control_Mshreg_scslll_103_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_Mshreg_scslll_103_FFY_RST
    );
  mac_control_txfifowerr_cntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(10),
      CE => mac_control_txfifowerr_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_11_FFY_RST,
      O => mac_control_txfifowerr_cntl(10)
    );
  mac_control_txfifowerr_cntl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_11_FFY_RST
    );
  mac_control_rxoferr_cntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(1),
      CE => mac_control_rxoferr_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_1_FFX_RST,
      O => mac_control_rxoferr_cntl(1)
    );
  mac_control_rxoferr_cntl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_1_FFX_RST
    );
  mac_control_rxoferr_cntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(3),
      CE => mac_control_rxoferr_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_3_FFX_RST,
      O => mac_control_rxoferr_cntl(3)
    );
  mac_control_rxoferr_cntl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_3_FFX_RST
    );
  mac_control_rxoferr_cntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(5),
      CE => mac_control_rxoferr_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_5_FFX_RST,
      O => mac_control_rxoferr_cntl(5)
    );
  mac_control_rxoferr_cntl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_5_FFX_RST
    );
  mac_control_rxoferr_cntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(7),
      CE => mac_control_rxoferr_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_7_FFX_RST,
      O => mac_control_rxoferr_cntl(7)
    );
  mac_control_rxoferr_cntl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_7_FFX_RST
    );
  mac_control_rxoferr_cntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(9),
      CE => mac_control_rxoferr_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_9_FFX_RST,
      O => mac_control_rxoferr_cntl(9)
    );
  mac_control_rxoferr_cntl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_9_FFX_RST
    );
  mac_control_PHY_status_rwl_1651 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(5),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_rwl_FFY_RST,
      O => mac_control_PHY_status_rwl
    );
  mac_control_PHY_status_rwl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_rwl_FFY_RST
    );
  tx_output_crcl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_2_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_2_FFY_RST,
      O => tx_output_crcl(2)
    );
  tx_output_crcl_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_2_FFY_RST
    );
  tx_output_TXD_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_4_OD,
      CE => TXD_4_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_4_OFF_RST,
      O => tx_output_TXD_4_OBUF
    );
  TXD_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_4_OFF_RST
    );
  tx_output_TXD_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_5_OD,
      CE => TXD_5_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_5_OFF_RST,
      O => tx_output_TXD_5_OBUF
    );
  TXD_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_5_OFF_RST
    );
  tx_output_TXD_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_6_OD,
      CE => TXD_6_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_6_OFF_RST,
      O => tx_output_TXD_6_OBUF
    );
  TXD_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_6_OFF_RST
    );
  tx_output_TXD_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_7_OD,
      CE => TXD_7_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_7_OFF_RST,
      O => tx_output_TXD_7_OBUF
    );
  TXD_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_7_OFF_RST
    );
  mac_control_LEDDPX : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDDPX_OD,
      CE => LEDDPX_OCEMUXNOT,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => LEDDPX_OFF_RST,
      O => mac_control_LEDDPX_OBUF
    );
  LEDDPX_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDDPX_OFF_RST
    );
  rx_output_bpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(1),
      CE => rxfbbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_1_FFX_RST,
      O => rxfbbp(1)
    );
  rxfbbp_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_1_FFX_RST
    );
  tx_output_bcntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_46,
      CE => tx_output_bcntl_8_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_8_FFX_RST,
      O => tx_output_bcntl(8)
    );
  tx_output_bcntl_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_8_FFX_RST
    );
  rx_output_bpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(3),
      CE => rxfbbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_3_FFX_RST,
      O => rxfbbp(3)
    );
  rxfbbp_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_3_FFX_RST
    );
  tx_output_datal_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(1),
      CE => tx_output_datal_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_1_FFX_RST,
      O => tx_output_datal(1)
    );
  tx_output_datal_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_1_FFX_RST
    );
  tx_output_bcntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_48,
      CE => tx_output_bcntl_10_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcntl_10_FFX_RST,
      O => tx_output_bcntl(10)
    );
  tx_output_bcntl_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcntl_10_FFX_RST
    );
  rx_output_bpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(5),
      CE => rxfbbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_5_FFX_RST,
      O => rxfbbp(5)
    );
  rxfbbp_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_5_FFX_RST
    );
  tx_output_datal_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(3),
      CE => tx_output_datal_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_3_FFX_RST,
      O => tx_output_datal(3)
    );
  tx_output_datal_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_3_FFX_RST
    );
  rx_output_fifo_BU301 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N2,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1610_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1610
    );
  rx_output_fifo_N1610_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1610_FFX_SET
    );
  rx_output_fifo_BU318 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1547,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1563_FFX_RST,
      O => rx_output_fifo_N1563
    );
  rx_output_fifo_N1563_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1563_FFX_RST
    );
  rx_output_fifo_BU170 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1610,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1627_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1626
    );
  rx_output_fifo_N1627_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1627_FFY_SET
    );
  rx_output_fifo_BU310 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1551,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1567_FFX_RST,
      O => rx_output_fifo_N1567
    );
  rx_output_fifo_N1567_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1567_FFX_RST
    );
  memcontroller_Q2_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(10),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_11_FFY_RST,
      O => q2(10)
    );
  q2_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_11_FFY_RST
    );
  rx_output_fifo_BU167 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1611,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1627_FFX_RST,
      O => rx_output_fifo_N1627
    );
  rx_output_fifo_N1627_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1627_FFX_RST
    );
  memcontroller_Q2_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(11),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_11_FFX_RST,
      O => q2(11)
    );
  q2_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_11_FFX_RST
    );
  rx_output_fifo_BU308 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1552,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1569_FFY_RST,
      O => rx_output_fifo_N1568
    );
  rx_output_fifo_N1569_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1569_FFY_RST
    );
  rx_output_fifo_BU314 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1549,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1565_FFX_RST,
      O => rx_output_fifo_N1565
    );
  rx_output_fifo_N1565_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1565_FFX_RST
    );
  rx_output_fifo_BU368 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N5,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1605_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1605
    );
  rx_output_fifo_N1605_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1605_FFX_SET
    );
  rx_output_fifo_BU360 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N9,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1609_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1609
    );
  rx_output_fifo_N1609_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1609_FFX_SET
    );
  mac_control_PHY_status_PHYSTAT_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(5),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_21_FFX_RST,
      O => mac_control_phystat(21)
    );
  mac_control_phystat_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_21_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(13),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_13_FFX_RST,
      O => mac_control_phystat(13)
    );
  mac_control_phystat_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_13_FFX_RST
    );
  memcontroller_Q2_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(27),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_27_FFX_RST,
      O => q2(27)
    );
  q2_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_27_FFX_RST
    );
  memcontroller_Q2_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(19),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_19_FFX_RST,
      O => q2(19)
    );
  q2_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_19_FFX_RST
    );
  memcontroller_Q3_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(11),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_11_FFX_RST,
      O => q3(11)
    );
  q3_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_11_FFX_RST
    );
  rx_output_fifo_BU378 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1553,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1585_FFX_RST,
      O => rx_output_fifo_N1585
    );
  rx_output_fifo_N1585_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1585_FFX_RST
    );
  rx_input_memio_macnt_79_1652 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_228,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_79_FFX_RST,
      O => rx_input_memio_macnt_79
    );
  rx_input_memio_macnt_79_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_79_FFX_RST
    );
  rx_input_memio_macnt_81_1653 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_230,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_81_FFX_RST,
      O => rx_input_memio_macnt_81
    );
  rx_input_memio_macnt_81_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_81_FFX_RST
    );
  rx_input_memio_macnt_83_1654 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_232,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_83_FFX_RST,
      O => rx_input_memio_macnt_83
    );
  rx_input_memio_macnt_83_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_83_FFX_RST
    );
  rx_input_memio_macnt_85_1655 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_234,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_85_FFX_RST,
      O => rx_input_memio_macnt_85
    );
  rx_input_memio_macnt_85_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_85_FFX_RST
    );
  rx_output_fifo_BU392 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1546,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1579_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1578
    );
  rx_output_fifo_N1579_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1579_FFY_SET
    );
  rx_output_fifo_BU390 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1547,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1579_FFX_RST,
      O => rx_output_fifo_N1579
    );
  rx_output_fifo_N1579_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1579_FFX_RST
    );
  rx_output_fifo_BU384 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1550,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1583_FFY_RST,
      O => rx_output_fifo_N1582
    );
  rx_output_fifo_N1583_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1583_FFY_RST
    );
  rx_output_fifo_BU382 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1551,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1583_FFX_RST,
      O => rx_output_fifo_N1583
    );
  rx_output_fifo_N1583_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1583_FFX_RST
    );
  memcontroller_Q3_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(23),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_23_FFY_RST,
      O => q3(23)
    );
  q3_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_23_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(10),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_27_FFY_RST,
      O => mac_control_phystat(26)
    );
  mac_control_phystat_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_27_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(11),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_27_FFX_RST,
      O => mac_control_phystat(27)
    );
  mac_control_phystat_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_27_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(3),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_19_FFX_RST,
      O => mac_control_phystat(19)
    );
  mac_control_phystat_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_19_FFX_RST
    );
  memcontroller_Q3_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(25),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_25_FFX_RST,
      O => q3(25)
    );
  q3_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_25_FFX_RST
    );
  memcontroller_Q3_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(17),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_17_FFX_RST,
      O => q3(17)
    );
  q3_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_17_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(13),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_29_FFX_RST,
      O => mac_control_phystat(29)
    );
  mac_control_phystat_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_29_FFX_RST
    );
  rx_output_bpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(7),
      CE => rxfbbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_7_FFX_RST,
      O => rxfbbp(7)
    );
  rxfbbp_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_7_FFX_RST
    );
  tx_output_datal_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(5),
      CE => tx_output_datal_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_5_FFX_RST,
      O => tx_output_datal(5)
    );
  tx_output_datal_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_5_FFX_RST
    );
  rx_output_bpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(9),
      CE => rxfbbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_9_FFX_RST,
      O => rxfbbp(9)
    );
  rxfbbp_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_9_FFX_RST
    );
  rx_output_bpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_bp(8),
      CE => rxfbbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfbbp_9_FFY_RST,
      O => rxfbbp(8)
    );
  rxfbbp_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfbbp_9_FFY_RST
    );
  tx_output_datal_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_data(7),
      CE => tx_output_datal_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_datal_7_FFX_RST,
      O => tx_output_datal(7)
    );
  tx_output_datal_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_datal_7_FFX_RST
    );
  mac_control_rxfifowerr_cntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(1),
      CE => mac_control_rxfifowerr_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_1_FFX_RST,
      O => mac_control_rxfifowerr_cntl(1)
    );
  mac_control_rxfifowerr_cntl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_1_FFX_RST
    );
  mac_control_rxfifowerr_cntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(3),
      CE => mac_control_rxfifowerr_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_3_FFX_RST,
      O => mac_control_rxfifowerr_cntl(3)
    );
  mac_control_rxfifowerr_cntl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_3_FFX_RST
    );
  mac_control_rxfifowerr_cntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(4),
      CE => mac_control_rxfifowerr_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_5_FFY_RST,
      O => mac_control_rxfifowerr_cntl(4)
    );
  mac_control_rxfifowerr_cntl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_5_FFY_RST
    );
  memcontroller_Q3_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(27),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_27_FFX_RST,
      O => q3(27)
    );
  q3_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_27_FFX_RST
    );
  memcontroller_Q3_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(19),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_19_FFX_RST,
      O => q3(19)
    );
  q3_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_19_FFX_RST
    );
  rx_output_fifo_BU386 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1549,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1581_FFX_RST,
      O => rx_output_fifo_N1581
    );
  rx_output_fifo_N1581_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1581_FFX_RST
    );
  memcontroller_Q3_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(29),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_29_FFX_RST,
      O => q3(29)
    );
  q3_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_29_FFX_RST
    );
  rx_output_ceinll_1656 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_ceinl,
      CE => rx_output_ceinll_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_ceinll_FFY_RST,
      O => rx_output_ceinll
    );
  rx_output_ceinll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_ceinll_FFY_RST
    );
  tx_output_data_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_ldata(5),
      CE => tx_output_data_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_data_5_FFY_RST,
      O => tx_output_data(5)
    );
  tx_output_data_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_data_5_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd3_1657 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_cs_FFd3_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_cs_FFd3
    );
  mac_control_PHY_status_MII_Interface_cs_FFd3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_MII_Interface_cs_FFd3_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(7),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_23_FFX_RST,
      O => mac_control_phystat(23)
    );
  mac_control_phystat_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_23_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(15),
      CE => mac_control_PHY_status_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_31_FFX_RST,
      O => mac_control_phystat(31)
    );
  mac_control_phystat_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_31_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(15),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_15_FFX_RST,
      O => mac_control_phystat(15)
    );
  mac_control_phystat_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_15_FFX_RST
    );
  rx_output_fifo_BU346 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1563,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1571_FFX_RST,
      O => rx_output_fifo_N1571
    );
  rx_output_fifo_N1571_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1571_FFX_RST
    );
  memcontroller_Q2_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(29),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_29_FFX_RST,
      O => q2(29)
    );
  q2_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_29_FFX_RST
    );
  memcontroller_Q3_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(21),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_21_FFX_RST,
      O => q3(21)
    );
  q3_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_21_FFX_RST
    );
  memcontroller_Q3_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(13),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_13_FFX_RST,
      O => q3(13)
    );
  q3_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_13_FFX_RST
    );
  rx_output_fifo_BU470 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1578,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1586_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1586
    );
  rx_output_fifo_N1586_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1586_FFX_SET
    );
  mac_control_LEDACT : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDACT_OD,
      CE => LEDACT_OCEMUXNOT,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => LEDACT_OFF_RST,
      O => mac_control_LEDACT_OBUF
    );
  LEDACT_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDACT_OFF_RST
    );
  tx_output_TXD_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_0_OD,
      CE => TXD_0_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_0_OFF_RST,
      O => tx_output_TXD_0_OBUF
    );
  TXD_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_0_OFF_RST
    );
  tx_output_TXD_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_1_OD,
      CE => TXD_1_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_1_OFF_RST,
      O => tx_output_TXD_1_OBUF
    );
  TXD_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_1_OFF_RST
    );
  tx_output_TXD_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_2_OD,
      CE => TXD_2_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_2_OFF_RST,
      O => tx_output_TXD_2_OBUF
    );
  TXD_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_2_OFF_RST
    );
  tx_output_TXD_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TXD_3_OD,
      CE => TXD_3_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TXD_3_OFF_RST,
      O => tx_output_TXD_3_OBUF
    );
  TXD_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TXD_3_OFF_RST
    );
  mac_control_txf_cntl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(31),
      CE => mac_control_txf_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_31_FFX_RST,
      O => mac_control_txf_cntl(31)
    );
  mac_control_txf_cntl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_31_FFX_RST
    );
  mac_control_txf_cntl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(23),
      CE => mac_control_txf_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_23_FFX_RST,
      O => mac_control_txf_cntl(23)
    );
  mac_control_txf_cntl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_23_FFX_RST
    );
  mac_control_txf_cntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(15),
      CE => mac_control_txf_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_15_FFX_RST,
      O => mac_control_txf_cntl(15)
    );
  mac_control_txf_cntl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_15_FFX_RST
    );
  mac_control_txf_cntl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(25),
      CE => mac_control_txf_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_25_FFX_RST,
      O => mac_control_txf_cntl(25)
    );
  mac_control_txf_cntl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_25_FFX_RST
    );
  mac_control_txf_cntl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(26),
      CE => mac_control_txf_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_27_FFY_RST,
      O => mac_control_txf_cntl(26)
    );
  mac_control_txf_cntl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_27_FFY_RST
    );
  mac_control_txf_cntl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(17),
      CE => mac_control_txf_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_17_FFX_RST,
      O => mac_control_txf_cntl(17)
    );
  mac_control_txf_cntl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_17_FFX_RST
    );
  mac_control_txf_cntl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(18),
      CE => mac_control_txf_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_19_FFY_RST,
      O => mac_control_txf_cntl(18)
    );
  mac_control_txf_cntl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_19_FFY_RST
    );
  mac_control_txf_cntl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(27),
      CE => mac_control_txf_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_27_FFX_RST,
      O => mac_control_txf_cntl(27)
    );
  mac_control_txf_cntl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_27_FFX_RST
    );
  rx_output_mdl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(27),
      CE => rx_output_mdl_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_27_FFX_RST,
      O => rx_output_mdl(27)
    );
  rx_output_mdl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_27_FFX_RST
    );
  rx_output_mdl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(19),
      CE => rx_output_mdl_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_19_FFX_RST,
      O => rx_output_mdl(19)
    );
  rx_output_mdl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_19_FFX_RST
    );
  rx_output_mdl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(29),
      CE => rx_output_mdl_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_29_FFX_RST,
      O => rx_output_mdl(29)
    );
  rx_output_mdl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_29_FFX_RST
    );
  tx_output_cs_FFd1_1658 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd2,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd2_FFY_RST,
      O => tx_output_cs_FFd1
    );
  tx_output_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd2_FFY_RST
    );
  tx_output_cs_FFd9_1659 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd10,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd10_FFY_RST,
      O => tx_output_cs_FFd9
    );
  tx_output_cs_FFd10_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd10_FFY_RST
    );
  tx_output_cs_FFd2_1660 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd3,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd2_FFX_RST,
      O => tx_output_cs_FFd2
    );
  tx_output_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd2_FFX_RST
    );
  tx_output_cs_FFd3_1661 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd7,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd3_FFY_RST,
      O => tx_output_cs_FFd3
    );
  tx_output_cs_FFd3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd3_FFY_RST
    );
  tx_output_cs_FFd10_1662 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd11,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd10_FFX_RST,
      O => tx_output_cs_FFd10
    );
  tx_output_cs_FFd10_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd10_FFX_RST
    );
  tx_input_enable_1663 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_enable_LOGIC_ONE,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => tx_input_enable,
      O => tx_input_enable
    );
  rx_input_memio_crcl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_2_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_2_FFY_RST,
      O => rx_input_memio_crcl(2)
    );
  rx_input_memio_crcl_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_2_FFY_RST
    );
  rx_input_memio_crcl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_3_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_3_FFY_RST,
      O => rx_input_memio_crcl(3)
    );
  rx_input_memio_crcl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_3_FFY_RST
    );
  mac_control_txf_cntl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(19),
      CE => mac_control_txf_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_19_FFX_RST,
      O => mac_control_txf_cntl(19)
    );
  mac_control_txf_cntl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_19_FFX_RST
    );
  mac_control_txf_cntl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(29),
      CE => mac_control_txf_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_29_FFX_RST,
      O => mac_control_txf_cntl(29)
    );
  mac_control_txf_cntl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_29_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_sin,
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MDIO_IFF_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(0)
    );
  MDIO_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MDIO_IFF_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_37_1664 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_170,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_37_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_37
    );
  mac_control_PHY_status_MII_Interface_mdccnt_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_37_FFX_RST
    );
  tx_output_crcl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_10_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_10_FFY_RST,
      O => tx_output_crcl(10)
    );
  tx_output_crcl_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_10_FFY_RST
    );
  rx_output_len_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(10),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_11_FFY_RST,
      O => rx_output_len(10)
    );
  rx_output_len_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_11_FFY_RST
    );
  rx_output_len_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(11),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_11_FFX_RST,
      O => rx_output_len(11)
    );
  rx_output_len_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_11_FFX_RST
    );
  rx_output_mdl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(11),
      CE => rx_output_mdl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_11_FFX_RST,
      O => rx_output_mdl(11)
    );
  rx_output_mdl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_11_FFX_RST
    );
  rx_output_len_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(12),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_13_FFY_RST,
      O => rx_output_len(12)
    );
  rx_output_len_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_13_FFY_RST
    );
  rx_output_len_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(13),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_13_FFX_RST,
      O => rx_output_len(13)
    );
  rx_output_len_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_13_FFX_RST
    );
  rx_output_mdl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(21),
      CE => rx_output_mdl_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_21_FFX_RST,
      O => rx_output_mdl(21)
    );
  rx_output_mdl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_21_FFX_RST
    );
  mac_control_LED1000 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LED1000_OD,
      CE => LED1000_OCEMUXNOT,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => LED1000_OFF_RST,
      O => mac_control_LED1000_OBUF
    );
  LED1000_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LED1000_OFF_RST
    );
  tx_output_TXEN_1665 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => TX_EN_OD,
      CE => TX_EN_OCEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => TX_EN_OFF_RST,
      O => tx_output_TXEN
    );
  TX_EN_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => TX_EN_OFF_RST
    );
  rx_output_DOUTEN : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUTEN_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUTEN_OFF_RST,
      O => rx_output_DOUTEN_OBUF
    );
  DOUTEN_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUTEN_OFF_RST
    );
  memcontroller_we_1666 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => MWE_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => MWE_OFF_SET,
      RST => GND,
      O => memcontroller_we
    );
  MWE_OFF_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => MWE_OFF_SET
    );
  rx_output_nf_1667 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_NEXTFRAME_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => NEXTFRAME_IFF_RST,
      O => rx_output_nf
    );
  NEXTFRAME_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => NEXTFRAME_IFF_RST
    );
  rx_output_mdl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(13),
      CE => rx_output_mdl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_13_FFX_RST,
      O => rx_output_mdl(13)
    );
  rx_output_mdl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_13_FFX_RST
    );
  rx_output_len_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(14),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_15_FFY_RST,
      O => rx_output_len(14)
    );
  rx_output_len_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_15_FFY_RST
    );
  rx_output_len_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(15),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_15_FFX_RST,
      O => rx_output_len(15)
    );
  rx_output_len_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_15_FFX_RST
    );
  rx_output_mdl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(31),
      CE => rx_output_mdl_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_31_FFX_RST,
      O => rx_output_mdl(31)
    );
  rx_output_mdl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_31_FFX_RST
    );
  rx_output_mdl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(23),
      CE => rx_output_mdl_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_23_FFX_RST,
      O => rx_output_mdl(23)
    );
  rx_output_mdl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_23_FFX_RST
    );
  rx_output_mdl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(15),
      CE => rx_output_mdl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_15_FFX_RST,
      O => rx_output_mdl(15)
    );
  rx_output_mdl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_15_FFX_RST
    );
  rx_output_mdl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(24),
      CE => rx_output_mdl_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_25_FFY_RST,
      O => rx_output_mdl(24)
    );
  rx_output_mdl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_25_FFY_RST
    );
  rx_output_mdl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(25),
      CE => rx_output_mdl_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_25_FFX_RST,
      O => rx_output_mdl(25)
    );
  rx_output_mdl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_25_FFX_RST
    );
  rx_output_mdl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(17),
      CE => rx_output_mdl_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_17_FFX_RST,
      O => rx_output_mdl(17)
    );
  rx_output_mdl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_17_FFX_RST
    );
  memcontroller_dnl1_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(7),
      CE => memcontroller_dnl1_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_7_FFX_RST,
      O => memcontroller_dnl1(7)
    );
  memcontroller_dnl1_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_7_FFX_RST
    );
  memcontroller_dnl1_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(27),
      CE => memcontroller_dnl1_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_27_FFX_RST,
      O => memcontroller_dnl1(27)
    );
  memcontroller_dnl1_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_27_FFX_RST
    );
  memcontroller_dnl1_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(19),
      CE => memcontroller_dnl1_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_19_FFX_RST,
      O => memcontroller_dnl1(19)
    );
  memcontroller_dnl1_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_19_FFX_RST
    );
  memcontroller_dnl1_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(8),
      CE => memcontroller_dnl1_8_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_8_FFX_RST,
      O => memcontroller_dnl1(8)
    );
  memcontroller_dnl1_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_8_FFX_RST
    );
  memcontroller_dnl1_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(28),
      CE => memcontroller_dnl1_28_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_28_FFX_RST,
      O => memcontroller_dnl1(28)
    );
  memcontroller_dnl1_28_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_28_FFX_RST
    );
  rx_output_DOUT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_10_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_10_OFF_RST,
      O => rx_output_DOUT_10_OBUF
    );
  DOUT_10_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_10_OFF_RST
    );
  rx_output_DOUT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_11_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_11_OFF_RST,
      O => rx_output_DOUT_11_OBUF
    );
  DOUT_11_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_11_OFF_RST
    );
  rx_output_DOUT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_12_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_12_OFF_RST,
      O => rx_output_DOUT_12_OBUF
    );
  DOUT_12_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_12_OFF_RST
    );
  rx_output_DOUT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_13_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_13_OFF_RST,
      O => rx_output_DOUT_13_OBUF
    );
  DOUT_13_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_13_OFF_RST
    );
  rx_output_DOUT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_14_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_14_OFF_RST,
      O => rx_output_DOUT_14_OBUF
    );
  DOUT_14_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_14_OFF_RST
    );
  rx_output_len_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(5),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_5_FFX_RST,
      O => rx_output_len(5)
    );
  rx_output_len_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_5_FFX_RST
    );
  rx_output_mdl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(5),
      CE => rx_output_mdl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_5_FFX_RST,
      O => rx_output_mdl(5)
    );
  rx_output_mdl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_5_FFX_RST
    );
  rx_output_len_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(7),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_7_FFX_RST,
      O => rx_output_len(7)
    );
  rx_output_len_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_7_FFX_RST
    );
  rx_output_mdl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(7),
      CE => rx_output_mdl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_7_FFX_RST,
      O => rx_output_mdl(7)
    );
  rx_output_mdl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_7_FFX_RST
    );
  rx_output_len_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(9),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_9_FFX_RST,
      O => rx_output_len(9)
    );
  rx_output_len_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_9_FFX_RST
    );
  rx_output_mdl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(9),
      CE => rx_output_mdl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_9_FFX_RST,
      O => rx_output_mdl(9)
    );
  rx_output_mdl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_9_FFX_RST
    );
  rx_input_GMII_ro_1668 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_ro_LOGIC_ONE,
      CE => rx_input_GMII_dvdelta,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_endf,
      O => rx_input_GMII_ro
    );
  rx_input_memio_crcl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_4_1_O,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_4_FFY_RST,
      O => rx_input_memio_crcl(4)
    );
  rx_input_memio_crcl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_4_FFY_RST
    );
  mac_control_rxfifowerr_cntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(5),
      CE => mac_control_rxfifowerr_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_5_FFX_RST,
      O => mac_control_rxfifowerr_cntl(5)
    );
  mac_control_rxfifowerr_cntl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_5_FFX_RST
    );
  mac_control_rxfifowerr_cntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(7),
      CE => mac_control_rxfifowerr_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_7_FFX_RST,
      O => mac_control_rxfifowerr_cntl(7)
    );
  mac_control_rxfifowerr_cntl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_7_FFX_RST
    );
  mac_control_rxfifowerr_cntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt(9),
      CE => mac_control_rxfifowerr_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_cntl_9_FFX_RST,
      O => mac_control_rxfifowerr_cntl(9)
    );
  mac_control_rxfifowerr_cntl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_cntl_9_FFX_RST
    );
  rx_output_len_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(0),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_1_FFY_RST,
      O => rx_output_len(0)
    );
  rx_output_len_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_1_FFY_RST
    );
  rx_output_len_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(1),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_1_FFX_RST,
      O => rx_output_len(1)
    );
  rx_output_len_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_1_FFX_RST
    );
  rx_output_mdl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(1),
      CE => rx_output_mdl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_1_FFX_RST,
      O => rx_output_mdl(1)
    );
  rx_output_mdl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_1_FFX_RST
    );
  rx_output_len_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(3),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_3_FFX_RST,
      O => rx_output_len(3)
    );
  rx_output_len_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_3_FFX_RST
    );
  rx_output_len_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_mdl(4),
      CE => rx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_len_5_FFY_RST,
      O => rx_output_len(4)
    );
  rx_output_len_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_len_5_FFY_RST
    );
  rx_output_mdl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => q3(3),
      CE => rx_output_mdl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_mdl_3_FFX_RST,
      O => rx_output_mdl(3)
    );
  rx_output_mdl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_mdl_3_FFX_RST
    );
  rx_output_DOUT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_15_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_15_OFF_RST,
      O => rx_output_DOUT_15_OBUF
    );
  DOUT_15_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_15_OFF_RST
    );
  mac_control_LED100 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LED100_OD,
      CE => LED100_OCEMUXNOT,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => LED100_OFF_RST,
      O => mac_control_LED100_OBUF
    );
  LED100_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LED100_OFF_RST
    );
  tx_input_newframel_1669 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_NEWFRAME_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => NEWFRAME_IFF_RST,
      O => tx_input_newframel
    );
  NEWFRAME_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => NEWFRAME_IFF_RST
    );
  memcontroller_dnout_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_28_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_28_OFF_RST,
      O => memcontroller_dnout(28)
    );
  MD_28_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_28_OFF_RST
    );
  memcontroller_qn_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(29),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_29_IFF_RST,
      O => memcontroller_qn(29)
    );
  MD_29_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_29_IFF_RST
    );
  memcontroller_dnout_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_29_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_29_OFF_RST,
      O => memcontroller_dnout(29)
    );
  MD_29_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_29_OFF_RST
    );
  memcontroller_addr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_0_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_0_OFF_RST,
      O => memcontroller_addr(0)
    );
  MA_0_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_0_OFF_RST
    );
  memcontroller_addr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_1_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_1_OFF_RST,
      O => memcontroller_addr(1)
    );
  MA_1_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_1_OFF_RST
    );
  memcontroller_addr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_2_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_2_OFF_RST,
      O => memcontroller_addr(2)
    );
  MA_2_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_2_OFF_RST
    );
  memcontroller_dnout_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_23_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_23_OFF_RST,
      O => memcontroller_dnout(23)
    );
  MD_23_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_23_OFF_RST
    );
  memcontroller_qn_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_15_IFF_RST,
      O => memcontroller_qn(15)
    );
  MD_15_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_15_IFF_RST
    );
  memcontroller_dnout_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_15_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_15_OFF_RST,
      O => memcontroller_dnout(15)
    );
  MD_15_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_15_OFF_RST
    );
  memcontroller_qn_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(31),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_31_IFF_RST,
      O => memcontroller_qn(31)
    );
  MD_31_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_31_IFF_RST
    );
  memcontroller_dnout_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_31_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_31_OFF_RST,
      O => memcontroller_dnout(31)
    );
  MD_31_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_31_OFF_RST
    );
  memcontroller_qn_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(24),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_24_IFF_RST,
      O => memcontroller_qn(24)
    );
  MD_24_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_24_IFF_RST
    );
  memcontroller_addr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_3_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_3_OFF_RST,
      O => memcontroller_addr(3)
    );
  MA_3_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_3_OFF_RST
    );
  memcontroller_addr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_4_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_4_OFF_RST,
      O => memcontroller_addr(4)
    );
  MA_4_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_4_OFF_RST
    );
  memcontroller_addr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_5_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_5_OFF_RST,
      O => memcontroller_addr(5)
    );
  MA_5_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_5_OFF_RST
    );
  memcontroller_addr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_6_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_6_OFF_RST,
      O => memcontroller_addr(6)
    );
  MA_6_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_6_OFF_RST
    );
  memcontroller_addr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_7_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_7_OFF_RST,
      O => memcontroller_addr(7)
    );
  MA_7_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_7_OFF_RST
    );
  memcontroller_dnout_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_18_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_18_OFF_RST,
      O => memcontroller_dnout(18)
    );
  MD_18_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_18_OFF_RST
    );
  memcontroller_qn_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(26),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_26_IFF_RST,
      O => memcontroller_qn(26)
    );
  MD_26_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_26_IFF_RST
    );
  memcontroller_dnout_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_26_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_26_OFF_RST,
      O => memcontroller_dnout(26)
    );
  MD_26_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_26_OFF_RST
    );
  memcontroller_qn_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(19),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_19_IFF_RST,
      O => memcontroller_qn(19)
    );
  MD_19_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_19_IFF_RST
    );
  memcontroller_dnout_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_19_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_19_OFF_RST,
      O => memcontroller_dnout(19)
    );
  MD_19_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_19_OFF_RST
    );
  memcontroller_qn_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(27),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_27_IFF_RST,
      O => memcontroller_qn(27)
    );
  MD_27_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_27_IFF_RST
    );
  memcontroller_qn_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(28),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_28_IFF_RST,
      O => memcontroller_qn(28)
    );
  MD_28_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_28_IFF_RST
    );
  memcontroller_dnout_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_27_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_27_OFF_RST,
      O => memcontroller_dnout(27)
    );
  MD_27_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_27_OFF_RST
    );
  rx_input_GMII_rxdl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_0_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_0_IFF_RST,
      O => rx_input_GMII_rxdl(0)
    );
  RXD_0_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_0_IFF_RST
    );
  rx_input_GMII_rxdl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_1_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_1_IFF_RST,
      O => rx_input_GMII_rxdl(1)
    );
  RXD_1_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_1_IFF_RST
    );
  rx_input_GMII_rxdl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_2_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_2_IFF_RST,
      O => rx_input_GMII_rxdl(2)
    );
  RXD_2_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_2_IFF_RST
    );
  rx_input_GMII_rxdl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_3_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_3_IFF_RST,
      O => rx_input_GMII_rxdl(3)
    );
  RXD_3_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_3_IFF_RST
    );
  rx_input_GMII_rxdl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_4_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_4_IFF_RST,
      O => rx_input_GMII_rxdl(4)
    );
  RXD_4_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_4_IFF_RST
    );
  rx_input_GMII_rxdl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_5_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_5_IFF_RST,
      O => rx_input_GMII_rxdl(5)
    );
  RXD_5_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_5_IFF_RST
    );
  rx_input_GMII_rxdl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_6_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_6_IFF_RST,
      O => rx_input_GMII_rxdl(6)
    );
  RXD_6_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_6_IFF_RST
    );
  rx_input_GMII_rxdl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RXD_7_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RXD_7_IFF_RST,
      O => rx_input_GMII_rxdl(7)
    );
  RXD_7_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RXD_7_IFF_RST
    );
  tx_input_dinl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_10_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_10_IFF_RST,
      O => tx_input_dinl(10)
    );
  DIN_10_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_10_IFF_RST
    );
  tx_input_dinl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_11_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_11_IFF_RST,
      O => tx_input_dinl(11)
    );
  DIN_11_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_11_IFF_RST
    );
  tx_input_dinl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_12_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_12_IFF_RST,
      O => tx_input_dinl(12)
    );
  DIN_12_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_12_IFF_RST
    );
  tx_input_dinl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_13_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_13_IFF_RST,
      O => tx_input_dinl(13)
    );
  DIN_13_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_13_IFF_RST
    );
  tx_input_dinl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_14_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_14_IFF_RST,
      O => tx_input_dinl(14)
    );
  DIN_14_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_14_IFF_RST
    );
  tx_input_dinl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_15_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_15_IFF_RST,
      O => tx_input_dinl(15)
    );
  DIN_15_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_15_IFF_RST
    );
  rx_output_DOUT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_0_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_0_OFF_RST,
      O => rx_output_DOUT_0_OBUF
    );
  DOUT_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_0_OFF_RST
    );
  rx_output_DOUT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_1_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_1_OFF_RST,
      O => rx_output_DOUT_1_OBUF
    );
  DOUT_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_1_OFF_RST
    );
  rx_output_DOUT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_2_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_2_OFF_RST,
      O => rx_output_DOUT_2_OBUF
    );
  DOUT_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_2_OFF_RST
    );
  tx_input_dinl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_8_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_8_IFF_RST,
      O => tx_input_dinl(8)
    );
  DIN_8_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_8_IFF_RST
    );
  tx_input_dinl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_9_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_9_IFF_RST,
      O => tx_input_dinl(9)
    );
  DIN_9_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_9_IFF_RST
    );
  rx_input_GMII_rx_erl_1670 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RX_ER_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RX_ER_IFF_RST,
      O => rx_input_GMII_rx_erl
    );
  RX_ER_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RX_ER_IFF_RST
    );
  rx_input_GMII_rx_dvl_1671 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_RX_DV_IBUF,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => RX_DV_IFF_RST,
      O => rx_input_GMII_rx_dvl
    );
  RX_DV_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => RX_DV_IFF_RST
    );
  memcontroller_addr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_10_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_10_OFF_RST,
      O => memcontroller_addr(10)
    );
  MA_10_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_10_OFF_RST
    );
  memcontroller_addr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_11_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_11_OFF_RST,
      O => memcontroller_addr(11)
    );
  MA_11_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_11_OFF_RST
    );
  memcontroller_addr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_12_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_12_OFF_RST,
      O => memcontroller_addr(12)
    );
  MA_12_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_12_OFF_RST
    );
  memcontroller_addr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_13_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_13_OFF_RST,
      O => memcontroller_addr(13)
    );
  MA_13_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_13_OFF_RST
    );
  rx_output_DOUT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_8_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_8_OFF_RST,
      O => rx_output_DOUT_8_OBUF
    );
  DOUT_8_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_8_OFF_RST
    );
  rx_output_DOUT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => DOUT_9_OD,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DOUT_9_OFF_RST,
      O => rx_output_DOUT_9_OBUF
    );
  DOUT_9_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DOUT_9_OFF_RST
    );
  mac_control_SOUT : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => SOUT_OD,
      CE => SOUT_OCEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => SOUT_OFF_RST,
      O => mac_control_SOUT_OBUF
    );
  SOUT_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => SOUT_OFF_RST
    );
  mac_control_sclkl_1672 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => SCLK_IDELAY,
      CE => SCLK_ICEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => SCLK_IFF_RST,
      O => mac_control_sclkl
    );
  SCLK_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => SCLK_IFF_RST
    );
  mac_control_LEDRX : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDRX_OD,
      CE => LEDRX_OCEMUXNOT,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => LEDRX_OFF_RST,
      O => mac_control_LEDRX_OBUF
    );
  LEDRX_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDRX_OFF_RST
    );
  mac_control_txfifowerr_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(14),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(14)
    );
  mac_control_txfifowerr_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(16),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(16)
    );
  mac_control_txfifowerr_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(19),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(19)
    );
  mac_control_txfifowerr_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(23),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(23)
    );
  mac_control_txfifowerr_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(18),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(18)
    );
  mac_control_txfifowerr_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(21),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(21)
    );
  memcontroller_addr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_14_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_14_OFF_RST,
      O => memcontroller_addr(14)
    );
  MA_14_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_14_OFF_RST
    );
  memcontroller_addr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_15_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_15_OFF_RST,
      O => memcontroller_addr(15)
    );
  MA_15_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_15_OFF_RST
    );
  memcontroller_addr_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_16_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_16_OFF_RST,
      O => memcontroller_addr(16)
    );
  MA_16_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_16_OFF_RST
    );
  memcontroller_qn_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_10_IFF_RST,
      O => memcontroller_qn(10)
    );
  MD_10_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_10_IFF_RST
    );
  memcontroller_dnout_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_10_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_10_OFF_RST,
      O => memcontroller_dnout(10)
    );
  MD_10_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_10_OFF_RST
    );
  memcontroller_qn_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_11_IFF_RST,
      O => memcontroller_qn(11)
    );
  MD_11_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_11_IFF_RST
    );
  mac_control_LEDTX : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => LEDTX_OD,
      CE => LEDTX_OCEMUXNOT,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => LEDTX_OFF_RST,
      O => mac_control_LEDTX_OBUF
    );
  LEDTX_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => LEDTX_OFF_RST
    );
  tx_input_dinl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_0_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_0_IFF_RST,
      O => tx_input_dinl(0)
    );
  DIN_0_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_0_IFF_RST
    );
  tx_input_dinl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_1_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_1_IFF_RST,
      O => tx_input_dinl(1)
    );
  DIN_1_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_1_IFF_RST
    );
  tx_input_dinl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_2_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_2_IFF_RST,
      O => tx_input_dinl(2)
    );
  DIN_2_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_2_IFF_RST
    );
  tx_input_dinl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_3_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_3_IFF_RST,
      O => tx_input_dinl(3)
    );
  DIN_3_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_3_IFF_RST
    );
  tx_input_dinl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_4_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_4_IFF_RST,
      O => tx_input_dinl(4)
    );
  DIN_4_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_4_IFF_RST
    );
  tx_input_dinl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_5_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_5_IFF_RST,
      O => tx_input_dinl(5)
    );
  DIN_5_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_5_IFF_RST
    );
  tx_input_dinl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_6_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_6_IFF_RST,
      O => tx_input_dinl(6)
    );
  DIN_6_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_6_IFF_RST
    );
  tx_input_dinl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_DIN_7_IBUF,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => DIN_7_IFF_RST,
      O => tx_input_dinl(7)
    );
  DIN_7_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => DIN_7_IFF_RST
    );
  memcontroller_dnout_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_9_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_9_OFF_RST,
      O => memcontroller_dnout(9)
    );
  MD_9_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_9_OFF_RST
    );
  mac_control_dout_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(30),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_30_FFX_RST,
      O => mac_control_dout(30)
    );
  mac_control_dout_30_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_30_FFX_RST
    );
  memcontroller_dnout_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_1_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_1_OFF_RST,
      O => memcontroller_dnout(1)
    );
  MD_1_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_1_OFF_RST
    );
  memcontroller_qn_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_2_IFF_RST,
      O => memcontroller_qn(2)
    );
  MD_2_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_2_IFF_RST
    );
  memcontroller_dnout_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_2_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_2_OFF_RST,
      O => memcontroller_dnout(2)
    );
  MD_2_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_2_OFF_RST
    );
  memcontroller_qn_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_3_IFF_RST,
      O => memcontroller_qn(3)
    );
  MD_3_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_3_IFF_RST
    );
  memcontroller_dnout_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_3_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_3_OFF_RST,
      O => memcontroller_dnout(3)
    );
  MD_3_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_3_OFF_RST
    );
  memcontroller_qn_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_4_IFF_RST,
      O => memcontroller_qn(4)
    );
  MD_4_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_4_IFF_RST
    );
  memcontroller_qn_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_5_IFF_RST,
      O => memcontroller_qn(5)
    );
  MD_5_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_5_IFF_RST
    );
  memcontroller_dnout_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_4_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_4_OFF_RST,
      O => memcontroller_dnout(4)
    );
  MD_4_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_4_OFF_RST
    );
  memcontroller_addr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_8_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_8_OFF_RST,
      O => memcontroller_addr(8)
    );
  MA_8_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_8_OFF_RST
    );
  memcontroller_addr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MA_9_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MA_9_OFF_RST,
      O => memcontroller_addr(9)
    );
  MA_9_OFF_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => MA_9_OFF_RST
    );
  mac_control_PHYRESET : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => PHYRESET_OD,
      CE => mac_control_n0033,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => PHYRESET_OFF_RST,
      O => mac_control_PHYRESET_OBUF
    );
  PHYRESET_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => PHYRESET_OFF_RST
    );
  memcontroller_qn_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_0_IFF_RST,
      O => memcontroller_qn(0)
    );
  MD_0_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_0_IFF_RST
    );
  memcontroller_dnout_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_0_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_0_OFF_RST,
      O => memcontroller_dnout(0)
    );
  MD_0_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_0_OFF_RST
    );
  memcontroller_qn_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_1_IFF_RST,
      O => memcontroller_qn(1)
    );
  MD_1_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_1_IFF_RST
    );
  memcontroller_qn_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(16),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_16_IFF_RST,
      O => memcontroller_qn(16)
    );
  MD_16_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_16_IFF_RST
    );
  memcontroller_dnout_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_24_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_24_OFF_RST,
      O => memcontroller_dnout(24)
    );
  MD_24_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_24_OFF_RST
    );
  memcontroller_dnout_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_16_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_16_OFF_RST,
      O => memcontroller_dnout(16)
    );
  MD_16_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_16_OFF_RST
    );
  memcontroller_qn_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(17),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_17_IFF_RST,
      O => memcontroller_qn(17)
    );
  MD_17_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_17_IFF_RST
    );
  memcontroller_dnout_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_17_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_17_OFF_RST,
      O => memcontroller_dnout(17)
    );
  MD_17_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_17_OFF_RST
    );
  memcontroller_qn_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(25),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_25_IFF_RST,
      O => memcontroller_qn(25)
    );
  MD_25_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_25_IFF_RST
    );
  memcontroller_dnout_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_25_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_25_OFF_RST,
      O => memcontroller_dnout(25)
    );
  MD_25_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_25_OFF_RST
    );
  memcontroller_qn_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(18),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_18_IFF_RST,
      O => memcontroller_qn(18)
    );
  MD_18_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_18_IFF_RST
    );
  memcontroller_dnout_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_11_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_11_OFF_RST,
      O => memcontroller_dnout(11)
    );
  MD_11_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_11_OFF_RST
    );
  memcontroller_qn_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(20),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_20_IFF_RST,
      O => memcontroller_qn(20)
    );
  MD_20_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_20_IFF_RST
    );
  memcontroller_dnout_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_20_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_20_OFF_RST,
      O => memcontroller_dnout(20)
    );
  MD_20_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_20_OFF_RST
    );
  memcontroller_qn_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_12_IFF_RST,
      O => memcontroller_qn(12)
    );
  MD_12_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_12_IFF_RST
    );
  memcontroller_dnout_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_12_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_12_OFF_RST,
      O => memcontroller_dnout(12)
    );
  MD_12_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_12_OFF_RST
    );
  memcontroller_qn_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(21),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_21_IFF_RST,
      O => memcontroller_qn(21)
    );
  MD_21_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_21_IFF_RST
    );
  memcontroller_qn_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_13_IFF_RST,
      O => memcontroller_qn(13)
    );
  MD_13_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_13_IFF_RST
    );
  memcontroller_dnout_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_21_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_21_OFF_RST,
      O => memcontroller_dnout(21)
    );
  MD_21_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_21_OFF_RST
    );
  tx_output_addr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(8),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_8_FFX_RST,
      O => addr2ext(8)
    );
  addr2ext_8_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_8_FFX_RST
    );
  tx_output_addr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(10),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_10_FFX_RST,
      O => addr2ext(10)
    );
  addr2ext_10_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_10_FFX_RST
    );
  tx_output_addr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(12),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_12_FFX_RST,
      O => addr2ext(12)
    );
  addr2ext_12_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_12_FFX_RST
    );
  tx_output_addr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(15),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_14_FFY_RST,
      O => addr2ext(15)
    );
  addr2ext_14_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_14_FFY_RST
    );
  rx_input_memio_bcnt_86_1673 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_235,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_86_FFY_RST,
      O => rx_input_memio_bcnt_86
    );
  rx_input_memio_bcnt_86_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_86_FFY_RST
    );
  mac_control_dout_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(21),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_21_FFX_RST,
      O => mac_control_dout(21)
    );
  mac_control_dout_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_21_FFX_RST
    );
  mac_control_dout_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(22),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_22_FFX_RST,
      O => mac_control_dout(22)
    );
  mac_control_dout_22_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_22_FFX_RST
    );
  mac_control_dout_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(23),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_23_FFX_RST,
      O => mac_control_dout(23)
    );
  mac_control_dout_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_23_FFX_RST
    );
  mac_control_dout_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(20),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_20_FFX_RST,
      O => mac_control_dout(20)
    );
  mac_control_dout_20_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_20_FFX_RST
    );
  memcontroller_dnout_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_5_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_5_OFF_RST,
      O => memcontroller_dnout(5)
    );
  MD_5_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_5_OFF_RST
    );
  memcontroller_qn_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_6_IFF_RST,
      O => memcontroller_qn(6)
    );
  MD_6_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_6_IFF_RST
    );
  memcontroller_dnout_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_6_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_6_OFF_RST,
      O => memcontroller_dnout(6)
    );
  MD_6_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_6_OFF_RST
    );
  memcontroller_qn_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_7_IFF_RST,
      O => memcontroller_qn(7)
    );
  MD_7_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_7_IFF_RST
    );
  memcontroller_dnout_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_7_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_7_OFF_RST,
      O => memcontroller_dnout(7)
    );
  MD_7_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_7_OFF_RST
    );
  memcontroller_qn_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_8_IFF_RST,
      O => memcontroller_qn(8)
    );
  MD_8_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_8_IFF_RST
    );
  memcontroller_qn_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_q(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_9_IFF_RST,
      O => memcontroller_qn(9)
    );
  MD_9_IFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_9_IFF_RST
    );
  memcontroller_dnout_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => MD_8_OD,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => MD_8_OFF_RST,
      O => memcontroller_dnout(8)
    );
  MD_8_OFF_RSTOR : X_BUF
    port map (
      I => GSR,
      O => MD_8_OFF_RST
    );
  memcontroller_dnl1_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(20),
      CE => memcontroller_dnl1_20_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_20_FFX_RST,
      O => memcontroller_dnl1(20)
    );
  memcontroller_dnl1_20_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_20_FFX_RST
    );
  memcontroller_dnl1_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(2),
      CE => memcontroller_dnl1_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_2_FFX_RST,
      O => memcontroller_dnl1(2)
    );
  memcontroller_dnl1_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_2_FFX_RST
    );
  memcontroller_dnl1_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(21),
      CE => memcontroller_dnl1_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_21_FFX_RST,
      O => memcontroller_dnl1(21)
    );
  memcontroller_dnl1_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_21_FFX_RST
    );
  memcontroller_dnl1_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(13),
      CE => memcontroller_dnl1_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_13_FFX_RST,
      O => memcontroller_dnl1(13)
    );
  memcontroller_dnl1_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_13_FFX_RST
    );
  memcontroller_dnl1_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(30),
      CE => memcontroller_dnl1_30_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_30_FFX_RST,
      O => memcontroller_dnl1(30)
    );
  memcontroller_dnl1_30_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_30_FFX_RST
    );
  mac_control_dout_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(16),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_16_FFX_RST,
      O => mac_control_dout(16)
    );
  mac_control_dout_16_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_16_FFX_RST
    );
  mac_control_dout_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(24),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_24_FFX_RST,
      O => mac_control_dout(24)
    );
  mac_control_dout_24_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_24_FFX_RST
    );
  mac_control_dout_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(25),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_25_FFX_RST,
      O => mac_control_dout(25)
    );
  mac_control_dout_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_25_FFX_RST
    );
  mac_control_dout_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(17),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_17_FFX_RST,
      O => mac_control_dout(17)
    );
  mac_control_dout_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_17_FFX_RST
    );
  memcontroller_dnl1_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(10),
      CE => memcontroller_dnl1_10_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_10_FFX_RST,
      O => memcontroller_dnl1(10)
    );
  memcontroller_dnl1_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_10_FFX_RST
    );
  memcontroller_dnl1_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(1),
      CE => memcontroller_dnl1_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_1_FFX_RST,
      O => memcontroller_dnl1(1)
    );
  memcontroller_dnl1_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_1_FFX_RST
    );
  memcontroller_dnl1_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(11),
      CE => memcontroller_dnl1_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_11_FFX_RST,
      O => memcontroller_dnl1(11)
    );
  memcontroller_dnl1_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_11_FFX_RST
    );
  memcontroller_dnl1_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(0),
      CE => memcontroller_dnl1_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_0_FFX_RST,
      O => memcontroller_dnl1(0)
    );
  memcontroller_dnl1_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_0_FFX_RST
    );
  memcontroller_dnl1_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(12),
      CE => memcontroller_dnl1_12_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_12_FFX_RST,
      O => memcontroller_dnl1(12)
    );
  memcontroller_dnl1_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_12_FFX_RST
    );
  memcontroller_dnl1_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(25),
      CE => memcontroller_dnl1_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_25_FFX_RST,
      O => memcontroller_dnl1(25)
    );
  memcontroller_dnl1_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_25_FFX_RST
    );
  memcontroller_dnl1_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(17),
      CE => memcontroller_dnl1_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_17_FFX_RST,
      O => memcontroller_dnl1(17)
    );
  memcontroller_dnl1_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_17_FFX_RST
    );
  memcontroller_dnl1_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(6),
      CE => memcontroller_dnl1_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_6_FFX_RST,
      O => memcontroller_dnl1(6)
    );
  memcontroller_dnl1_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_6_FFX_RST
    );
  memcontroller_dnl1_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(26),
      CE => memcontroller_dnl1_26_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_26_FFX_RST,
      O => memcontroller_dnl1(26)
    );
  memcontroller_dnl1_26_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_26_FFX_RST
    );
  memcontroller_dnl1_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(18),
      CE => memcontroller_dnl1_18_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_18_FFX_RST,
      O => memcontroller_dnl1(18)
    );
  memcontroller_dnl1_18_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_18_FFX_RST
    );
  memcontroller_dnl1_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(22),
      CE => memcontroller_dnl1_22_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_22_FFX_RST,
      O => memcontroller_dnl1(22)
    );
  memcontroller_dnl1_22_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_22_FFX_RST
    );
  memcontroller_dnl1_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(14),
      CE => memcontroller_dnl1_14_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_14_FFX_RST,
      O => memcontroller_dnl1(14)
    );
  memcontroller_dnl1_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_14_FFX_RST
    );
  memcontroller_dnl1_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(31),
      CE => memcontroller_dnl1_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_31_FFX_RST,
      O => memcontroller_dnl1(31)
    );
  memcontroller_dnl1_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_31_FFX_RST
    );
  memcontroller_dnl1_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(15),
      CE => memcontroller_dnl1_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_15_FFX_RST,
      O => memcontroller_dnl1(15)
    );
  memcontroller_dnl1_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_15_FFX_RST
    );
  memcontroller_dnl1_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(23),
      CE => memcontroller_dnl1_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_23_FFX_RST,
      O => memcontroller_dnl1(23)
    );
  memcontroller_dnl1_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_23_FFX_RST
    );
  mac_control_dout_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(18),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_18_FFX_RST,
      O => mac_control_dout(18)
    );
  mac_control_dout_18_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_18_FFX_RST
    );
  mac_control_dout_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(26),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_26_FFX_RST,
      O => mac_control_dout(26)
    );
  mac_control_dout_26_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_26_FFX_RST
    );
  mac_control_dout_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(19),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_19_FFX_RST,
      O => mac_control_dout(19)
    );
  mac_control_dout_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_19_FFX_RST
    );
  mac_control_dout_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(27),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_27_FFX_RST,
      O => mac_control_dout(27)
    );
  mac_control_dout_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_27_FFX_RST
    );
  mac_control_dout_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(28),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_28_FFX_RST,
      O => mac_control_dout(28)
    );
  mac_control_dout_28_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_28_FFX_RST
    );
  mac_control_dout_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(29),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_29_FFX_RST,
      O => mac_control_dout(29)
    );
  mac_control_dout_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_29_FFX_RST
    );
  memcontroller_dnl1_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(3),
      CE => memcontroller_dnl1_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_3_FFX_RST,
      O => memcontroller_dnl1(3)
    );
  memcontroller_dnl1_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_3_FFX_RST
    );
  memcontroller_dnl1_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(4),
      CE => memcontroller_dnl1_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_4_FFX_RST,
      O => memcontroller_dnl1(4)
    );
  memcontroller_dnl1_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_4_FFX_RST
    );
  memcontroller_dnl1_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(24),
      CE => memcontroller_dnl1_24_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_24_FFX_RST,
      O => memcontroller_dnl1(24)
    );
  memcontroller_dnl1_24_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_24_FFX_RST
    );
  memcontroller_dnl1_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(16),
      CE => memcontroller_dnl1_16_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_16_FFX_RST,
      O => memcontroller_dnl1(16)
    );
  memcontroller_dnl1_16_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_16_FFX_RST
    );
  memcontroller_dnl1_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(5),
      CE => memcontroller_dnl1_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_5_FFX_RST,
      O => memcontroller_dnl1(5)
    );
  memcontroller_dnl1_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_5_FFX_RST
    );
  rx_input_memio_addrchk_datal_47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_47_FFX_RST,
      O => rx_input_memio_addrchk_datal(47)
    );
  rx_input_memio_addrchk_datal_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_47_FFX_RST
    );
  rx_input_memio_crcll_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(0),
      CE => rx_input_memio_crcll_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_1_FFY_RST,
      O => rx_input_memio_crcll(0)
    );
  rx_input_memio_crcll_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_1_FFY_RST
    );
  rx_input_memio_crcll_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(1),
      CE => rx_input_memio_crcll_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_1_FFX_RST,
      O => rx_input_memio_crcll(1)
    );
  rx_input_memio_crcll_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_1_FFX_RST
    );
  rx_input_memio_crcll_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(2),
      CE => rx_input_memio_crcll_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_3_FFY_RST,
      O => rx_input_memio_crcll(2)
    );
  rx_input_memio_crcll_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_3_FFY_RST
    );
  rx_input_memio_crcll_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(3),
      CE => rx_input_memio_crcll_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_3_FFX_RST,
      O => rx_input_memio_crcll(3)
    );
  rx_input_memio_crcll_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_3_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(0),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_1_FFY_RST,
      O => mac_control_phystat(0)
    );
  mac_control_phystat_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_1_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(1),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_1_FFX_RST,
      O => mac_control_phystat(1)
    );
  mac_control_phystat_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_1_FFX_RST
    );
  rx_input_memio_crcll_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(4),
      CE => rx_input_memio_crcll_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_5_FFY_RST,
      O => rx_input_memio_crcll(4)
    );
  rx_input_memio_crcll_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_5_FFY_RST
    );
  rx_input_memio_crcll_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(5),
      CE => rx_input_memio_crcll_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_5_FFX_RST,
      O => rx_input_memio_crcll(5)
    );
  rx_input_memio_crcll_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_5_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(2),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_3_FFY_RST,
      O => mac_control_phystat(2)
    );
  mac_control_phystat_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_3_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(3),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_3_FFX_RST,
      O => mac_control_phystat(3)
    );
  mac_control_phystat_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_3_FFX_RST
    );
  rx_input_memio_crcll_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(6),
      CE => rx_input_memio_crcll_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_7_FFY_RST,
      O => rx_input_memio_crcll(6)
    );
  rx_input_memio_crcll_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_7_FFY_RST
    );
  rx_input_memio_crcll_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(7),
      CE => rx_input_memio_crcll_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_7_FFX_RST,
      O => rx_input_memio_crcll(7)
    );
  rx_input_memio_crcll_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_7_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(4),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_5_FFY_RST,
      O => mac_control_phystat(4)
    );
  mac_control_phystat_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_5_FFY_RST
    );
  rx_input_memio_crcll_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(8),
      CE => rx_input_memio_crcll_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_9_FFY_RST,
      O => rx_input_memio_crcll(8)
    );
  rx_input_memio_crcll_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_9_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(5),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_5_FFX_RST,
      O => mac_control_phystat(5)
    );
  mac_control_phystat_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_5_FFX_RST
    );
  rx_input_memio_crcll_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(9),
      CE => rx_input_memio_crcll_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_9_FFX_RST,
      O => rx_input_memio_crcll(9)
    );
  rx_input_memio_crcll_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_9_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(6),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_7_FFY_RST,
      O => mac_control_phystat(6)
    );
  mac_control_phystat_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_7_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(7),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_7_FFX_RST,
      O => mac_control_phystat(7)
    );
  mac_control_phystat_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_7_FFX_RST
    );
  mac_control_PHY_status_PHYSTAT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(8),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_9_FFY_RST,
      O => mac_control_phystat(8)
    );
  mac_control_phystat_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_9_FFY_RST
    );
  mac_control_PHY_status_PHYSTAT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(9),
      CE => mac_control_PHY_status_n0019,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phystat_9_FFX_RST,
      O => mac_control_phystat(9)
    );
  mac_control_phystat_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phystat_9_FFX_RST
    );
  tx_output_crcl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_25_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_25_FFY_RST,
      O => tx_output_crcl(25)
    );
  tx_output_crcl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_25_FFY_RST
    );
  tx_output_crcl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_17_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_17_FFY_RST,
      O => tx_output_crcl(17)
    );
  tx_output_crcl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_17_FFY_RST
    );
  memcontroller_clknum_0_1_1674 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_0_1_BYMUXNOT,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_clknum_0_1_FFY_RST,
      O => memcontroller_clknum_0_1
    );
  memcontroller_clknum_0_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_0_1_FFY_RST
    );
  memcontroller_clknum_1_3_1675 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_n0149,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_clknum_1_3_FFY_RST,
      O => memcontroller_clknum_1_3
    );
  memcontroller_clknum_1_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_1_3_FFY_RST
    );
  rx_fifocheck_fbbpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_11_FFY_RST,
      O => rx_fifocheck_fbbpl(10)
    );
  rx_fifocheck_fbbpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_11_FFY_RST
    );
  rx_input_memio_doutl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(29),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_29_FFX_RST,
      O => rx_input_memio_doutl(29)
    );
  rx_input_memio_doutl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_29_FFX_RST
    );
  rx_input_fifo_control_d0_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(0),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_1_FFY_RST,
      O => rx_input_fifo_control_d0(0)
    );
  rx_input_fifo_control_d0_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_1_FFY_RST
    );
  rx_input_fifo_control_d0_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(1),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_1_FFX_RST,
      O => rx_input_fifo_control_d0(1)
    );
  rx_input_fifo_control_d0_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_1_FFX_RST
    );
  rx_input_fifo_control_d0_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(3),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_3_FFX_RST,
      O => rx_input_fifo_control_d0(3)
    );
  rx_input_fifo_control_d0_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_3_FFX_RST
    );
  rx_input_fifo_control_d0_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(5),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_5_FFX_RST,
      O => rx_input_fifo_control_d0(5)
    );
  rx_input_fifo_control_d0_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_5_FFX_RST
    );
  rx_input_fifo_control_d1_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(1),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_1_FFX_RST,
      O => rx_input_fifo_control_d1(1)
    );
  rx_input_fifo_control_d1_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_1_FFX_RST
    );
  rx_input_fifo_control_d0_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(6),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_7_FFY_RST,
      O => rx_input_fifo_control_d0(6)
    );
  rx_input_fifo_control_d0_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_7_FFY_RST
    );
  rx_input_fifo_control_d0_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(7),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_7_FFX_RST,
      O => rx_input_fifo_control_d0(7)
    );
  rx_input_fifo_control_d0_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_7_FFX_RST
    );
  rx_input_fifo_control_d1_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(4),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_5_FFY_RST,
      O => rx_input_fifo_control_d1(4)
    );
  rx_input_fifo_control_d1_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_5_FFY_RST
    );
  rx_input_fifo_control_d1_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(3),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_3_FFX_RST,
      O => rx_input_fifo_control_d1(3)
    );
  rx_input_fifo_control_d1_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_3_FFX_RST
    );
  rx_input_fifo_control_d0_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl(8),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d0_8_FFY_RST,
      O => rx_input_fifo_control_d0(8)
    );
  rx_input_fifo_control_d0_8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d0_8_FFY_RST
    );
  rx_input_fifo_control_d2_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(0),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_1_FFY_RST,
      O => rx_input_fifo_control_d2(0)
    );
  rx_input_fifo_control_d2_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_1_FFY_RST
    );
  rx_input_fifo_control_d0_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_dinl_9_rt,
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_control_d0_9_FFY_SET,
      RST => rx_input_fifo_control_d0_9_FFY_RST,
      O => rx_input_fifo_control_d0(9)
    );
  rx_input_fifo_control_d0_9_FFY_SETOR : X_BUF
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_d0_9_FFY_SET
    );
  rx_input_fifo_control_d0_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_control_d0_9_LOGIC_ZERO,
      I1 => GSR,
      O => rx_input_fifo_control_d0_9_FFY_RST
    );
  rx_input_fifo_control_d1_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(5),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_5_FFX_RST,
      O => rx_input_fifo_control_d1(5)
    );
  rx_input_fifo_control_d1_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_5_FFX_RST
    );
  tx_fifocheck_bpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_1_FFY_RST,
      O => tx_fifocheck_bpl(0)
    );
  tx_fifocheck_bpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_1_FFY_RST
    );
  tx_fifocheck_bpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_1_FFX_RST,
      O => tx_fifocheck_bpl(1)
    );
  tx_fifocheck_bpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_1_FFX_RST
    );
  tx_fifocheck_bpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_3_FFY_RST,
      O => tx_fifocheck_bpl(2)
    );
  tx_fifocheck_bpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_3_FFY_RST
    );
  tx_fifocheck_bpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_3_FFX_RST,
      O => tx_fifocheck_bpl(3)
    );
  tx_fifocheck_bpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_3_FFX_RST
    );
  tx_fifocheck_bpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_5_FFY_RST,
      O => tx_fifocheck_bpl(4)
    );
  tx_fifocheck_bpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_5_FFY_RST
    );
  tx_fifocheck_bpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_5_FFX_RST,
      O => tx_fifocheck_bpl(5)
    );
  tx_fifocheck_bpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_5_FFX_RST
    );
  tx_fifocheck_bpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_7_FFY_RST,
      O => tx_fifocheck_bpl(6)
    );
  tx_fifocheck_bpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_7_FFY_RST
    );
  tx_fifocheck_bpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_7_FFX_RST,
      O => tx_fifocheck_bpl(7)
    );
  tx_fifocheck_bpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_7_FFX_RST
    );
  tx_fifocheck_bpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_9_FFY_RST,
      O => tx_fifocheck_bpl(8)
    );
  tx_fifocheck_bpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_9_FFY_RST
    );
  tx_fifocheck_bpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_9_FFX_RST,
      O => tx_fifocheck_bpl(9)
    );
  tx_fifocheck_bpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_9_FFX_RST
    );
  tx_output_crcl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_29_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_29_FFY_RST,
      O => tx_output_crcl(29)
    );
  tx_output_crcl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_29_FFY_RST
    );
  rx_input_memio_crcll_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(11),
      CE => rx_input_memio_crcll_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_11_FFX_RST,
      O => rx_input_memio_crcll(11)
    );
  rx_input_memio_crcll_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_11_FFX_RST
    );
  rx_input_memio_crcll_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(10),
      CE => rx_input_memio_crcll_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_11_FFY_RST,
      O => rx_input_memio_crcll(10)
    );
  rx_input_memio_crcll_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_11_FFY_RST
    );
  rx_input_memio_crcll_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(12),
      CE => rx_input_memio_crcll_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_13_FFY_RST,
      O => rx_input_memio_crcll(12)
    );
  rx_input_memio_crcll_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_13_FFY_RST
    );
  tx_output_addr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(1),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_0_FFY_RST,
      O => addr2ext(1)
    );
  addr2ext_0_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_0_FFY_RST
    );
  tx_output_addr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(3),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_2_FFY_RST,
      O => addr2ext(3)
    );
  addr2ext_2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_2_FFY_RST
    );
  tx_output_addr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(7),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_6_FFY_RST,
      O => addr2ext(7)
    );
  addr2ext_6_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_6_FFY_RST
    );
  tx_output_addr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_Madd_n0000_inst_lut2_0,
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_0_FFX_RST,
      O => addr2ext(0)
    );
  addr2ext_0_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_0_FFX_RST
    );
  tx_output_addr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(2),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_2_FFX_RST,
      O => addr2ext(2)
    );
  addr2ext_2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_2_FFX_RST
    );
  tx_output_addr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_addr_n0000(5),
      CE => tx_output_addrinc,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr2ext_4_FFY_RST,
      O => addr2ext(5)
    );
  addr2ext_4_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => addr2ext_4_FFY_RST
    );
  rx_input_memio_bcnt_89_1676 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_238,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_89_FFX_RST,
      O => rx_input_memio_bcnt_89
    );
  rx_input_memio_bcnt_89_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_89_FFX_RST
    );
  rx_input_memio_bcnt_91_1677 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_240,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_91_FFX_RST,
      O => rx_input_memio_bcnt_91
    );
  rx_input_memio_bcnt_91_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_91_FFX_RST
    );
  rx_input_memio_bcnt_94_1678 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_243,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_93_FFY_RST,
      O => rx_input_memio_bcnt_94
    );
  rx_input_memio_bcnt_93_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_93_FFY_RST
    );
  rx_input_memio_bcnt_93_1679 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_242,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_93_FFX_RST,
      O => rx_input_memio_bcnt_93
    );
  rx_input_memio_bcnt_93_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_93_FFX_RST
    );
  rx_input_memio_bcnt_96_1680 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_245,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_95_FFY_RST,
      O => rx_input_memio_bcnt_96
    );
  rx_input_memio_bcnt_95_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_95_FFY_RST
    );
  rx_input_memio_bcnt_98_1681 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_247,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_97_FFY_RST,
      O => rx_input_memio_bcnt_98
    );
  rx_input_memio_bcnt_97_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_97_FFY_RST
    );
  mac_control_rxoferr_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(8),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(8)
    );
  mac_control_rxoferr_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(10),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(10)
    );
  mac_control_rxoferr_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(13),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(13)
    );
  mac_control_rxoferr_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(17),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(17)
    );
  mac_control_rxoferr_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(12),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(12)
    );
  mac_control_rxoferr_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(15),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(15)
    );
  memcontroller_dnl1_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(9),
      CE => memcontroller_dnl1_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_9_FFX_RST,
      O => memcontroller_dnl1(9)
    );
  memcontroller_dnl1_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_9_FFX_RST
    );
  memcontroller_dnl1_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dn(29),
      CE => memcontroller_dnl1_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl1_29_FFX_RST,
      O => memcontroller_dnl1(29)
    );
  memcontroller_dnl1_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl1_29_FFX_RST
    );
  rx_input_memio_bp_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(6),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_6_FFX_RST,
      O => rx_input_memio_bp(6)
    );
  rx_input_memio_bp_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_6_FFX_RST
    );
  rx_input_memio_bp_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(8),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_8_FFX_RST,
      O => rx_input_memio_bp(8)
    );
  rx_input_memio_bp_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_8_FFX_RST
    );
  rx_input_memio_bp_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(10),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_10_FFX_RST,
      O => rx_input_memio_bp(10)
    );
  rx_input_memio_bp_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_10_FFX_RST
    );
  mac_control_rxcrcerr_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(20),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(20)
    );
  mac_control_rxcrcerr_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(22),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(22)
    );
  mac_control_rxcrcerr_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(25),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(25)
    );
  mac_control_rxcrcerr_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(29),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(29)
    );
  mac_control_rxcrcerr_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(24),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(24)
    );
  mac_control_rxcrcerr_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(27),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(27)
    );
  mac_control_rxcrcerr_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(14),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(14)
    );
  mac_control_rxcrcerr_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(16),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(16)
    );
  mac_control_rxcrcerr_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(19),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(19)
    );
  mac_control_rxcrcerr_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(23),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(23)
    );
  mac_control_rxcrcerr_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(18),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(18)
    );
  mac_control_rxcrcerr_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(21),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(21)
    );
  mac_control_rxcrcerr_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(2),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(2)
    );
  mac_control_rxcrcerr_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(4),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(4)
    );
  mac_control_rxcrcerr_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(7),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(7)
    );
  mac_control_rxcrcerr_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(11),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(11)
    );
  mac_control_rxcrcerr_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(6),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(6)
    );
  mac_control_rxcrcerr_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(9),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(9)
    );
  mac_control_rxcrcerr_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(26),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(26)
    );
  mac_control_rxcrcerr_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(28),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(28)
    );
  mac_control_rxcrcerr_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(31),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(31)
    );
  mac_control_rxcrcerr_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(30),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(30)
    );
  rx_input_memio_bp_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(1),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_0_FFY_RST,
      O => rx_input_memio_bp(1)
    );
  rx_input_memio_bp_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_0_FFY_RST
    );
  mac_control_rxcrcerr_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(8),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(8)
    );
  mac_control_rxcrcerr_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(10),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(10)
    );
  mac_control_rxcrcerr_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(13),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(13)
    );
  mac_control_rxcrcerr_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(17),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(17)
    );
  mac_control_rxcrcerr_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(12),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(12)
    );
  mac_control_rxcrcerr_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(15),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(15)
    );
  mac_control_txfifowerr_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(8),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(8)
    );
  mac_control_txfifowerr_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(10),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(10)
    );
  mac_control_txfifowerr_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(13),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(13)
    );
  mac_control_txfifowerr_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(17),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(17)
    );
  mac_control_txfifowerr_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(12),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(12)
    );
  mac_control_txfifowerr_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(15),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(15)
    );
  rx_input_memio_bcnt_95_1682 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_244,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_95_FFX_RST,
      O => rx_input_memio_bcnt_95
    );
  rx_input_memio_bcnt_95_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_95_FFX_RST
    );
  rx_input_memio_bcnt_97_1683 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_246,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_97_FFX_RST,
      O => rx_input_memio_bcnt_97
    );
  rx_input_memio_bcnt_97_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_97_FFX_RST
    );
  rx_input_memio_bcnt_100_1684 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_249,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_99_FFY_RST,
      O => rx_input_memio_bcnt_100
    );
  rx_input_memio_bcnt_99_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_99_FFY_RST
    );
  rx_input_memio_bcnt_101_1685 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_250,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_101_FFX_RST,
      O => rx_input_memio_bcnt_101
    );
  rx_input_memio_bcnt_101_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_101_FFX_RST
    );
  rx_input_memio_bcnt_99_1686 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_248,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_99_FFX_RST,
      O => rx_input_memio_bcnt_99
    );
  rx_input_memio_bcnt_99_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_99_FFX_RST
    );
  rx_input_memio_bp_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(0),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_0_FFX_RST,
      O => rx_input_memio_bp(0)
    );
  rx_input_memio_bp_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_0_FFX_RST
    );
  rx_input_memio_bp_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(2),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_2_FFX_RST,
      O => rx_input_memio_bp(2)
    );
  rx_input_memio_bp_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_2_FFX_RST
    );
  rx_input_memio_bp_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0043(4),
      CE => rx_input_memio_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bp_4_FFX_RST,
      O => rx_input_memio_bp(4)
    );
  rx_input_memio_bp_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bp_4_FFX_RST
    );
  mac_control_rxcrcerr_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(1),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(1)
    );
  mac_control_rxcrcerr_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_Madd_n0000_inst_lut2_16,
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(0)
    );
  mac_control_rxcrcerr_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt_n0000(3),
      CE => rxcrcerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxcrcerr_rst,
      O => mac_control_rxcrcerr_cnt(3)
    );
  mac_control_rxoferr_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(14),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(14)
    );
  mac_control_rxoferr_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(16),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(16)
    );
  mac_control_rxoferr_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(19),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(19)
    );
  mac_control_rxoferr_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(23),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(23)
    );
  mac_control_rxoferr_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(18),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(18)
    );
  mac_control_rxoferr_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt_n0000(21),
      CE => rxoferr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxoferr_rst,
      O => mac_control_rxoferr_cnt(21)
    );
  mac_control_rxphyerr_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(4),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(4)
    );
  mac_control_rxphyerr_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(6),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(6)
    );
  mac_control_rxphyerr_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(13),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(13)
    );
  mac_control_rxphyerr_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(8),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(8)
    );
  mac_control_rxphyerr_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(11),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(11)
    );
  mac_control_rxphyerr_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(15),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(15)
    );
  mac_control_ledrx_cnt_165_1687 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_312,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_165_FFX_RST,
      O => mac_control_ledrx_cnt_165
    );
  mac_control_ledrx_cnt_165_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_165_FFX_RST
    );
  mac_control_ledrx_cnt_159_1688 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_306,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_159_FFX_RST,
      O => mac_control_ledrx_cnt_159
    );
  mac_control_ledrx_cnt_159_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_159_FFX_RST
    );
  mac_control_ledrx_cnt_161_1689 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_308,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_161_FFX_RST,
      O => mac_control_ledrx_cnt_161
    );
  mac_control_ledrx_cnt_161_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_161_FFX_RST
    );
  mac_control_ledrx_cnt_164_1690 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_311,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_163_FFY_RST,
      O => mac_control_ledrx_cnt_164
    );
  mac_control_ledrx_cnt_163_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_163_FFY_RST
    );
  mac_control_ledrx_cnt_163_1691 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledrx_cnt_inst_sum_310,
      CE => mac_control_n0039,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_cnt_163_FFX_RST,
      O => mac_control_ledrx_cnt_163
    );
  mac_control_ledrx_cnt_163_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_cnt_163_FFX_RST
    );
  mac_control_rxfifowerr_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(22),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(22)
    );
  mac_control_rxfifowerr_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(29),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(29)
    );
  mac_control_rxfifowerr_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(24),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(24)
    );
  mac_control_rxfifowerr_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(27),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(27)
    );
  mac_control_rxfifowerr_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(31),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(31)
    );
  mac_control_rxfifowerr_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(26),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(26)
    );
  mac_control_ledtx_cnt_147_1692 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_294,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_147_FFX_RST,
      O => mac_control_ledtx_cnt_147
    );
  mac_control_ledtx_cnt_147_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_147_FFX_RST
    );
  rx_output_fifo_BU47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1905,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N17_FFY_RST,
      O => rx_output_fifo_N16
    );
  rx_output_fifo_N17_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N17_FFY_RST
    );
  mac_control_ledtx_cnt_149_1693 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_296,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_149_FFX_RST,
      O => mac_control_ledtx_cnt_149
    );
  mac_control_ledtx_cnt_149_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_149_FFX_RST
    );
  mac_control_ledtx_cnt_152_1694 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_299,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_151_FFY_RST,
      O => mac_control_ledtx_cnt_152
    );
  mac_control_ledtx_cnt_151_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_151_FFY_RST
    );
  mac_control_ledtx_cnt_151_1695 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_298,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_151_FFX_RST,
      O => mac_control_ledtx_cnt_151
    );
  mac_control_ledtx_cnt_151_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_151_FFX_RST
    );
  mac_control_ledtx_cnt_153_1696 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_300,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_153_FFX_RST,
      O => mac_control_ledtx_cnt_153
    );
  mac_control_ledtx_cnt_153_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_153_FFX_RST
    );
  tx_fifocheck_diff_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_10_FFX_RST,
      O => tx_fifocheck_diff(10)
    );
  tx_fifocheck_diff_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_10_FFX_RST
    );
  tx_fifocheck_diff_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_12_FFX_RST,
      O => tx_fifocheck_diff(12)
    );
  tx_fifocheck_diff_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_12_FFX_RST
    );
  mac_control_ledtx_cnt_144_1697 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_291,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_143_FFY_RST,
      O => mac_control_ledtx_cnt_144
    );
  mac_control_ledtx_cnt_143_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_143_FFY_RST
    );
  tx_fifocheck_diff_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_14_FFX_RST,
      O => tx_fifocheck_diff(14)
    );
  tx_fifocheck_diff_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_14_FFX_RST
    );
  mac_control_rxfifowerr_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(10),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(10)
    );
  mac_control_rxfifowerr_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(17),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(17)
    );
  mac_control_rxfifowerr_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(12),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(12)
    );
  mac_control_rxfifowerr_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(15),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(15)
    );
  mac_control_rxfifowerr_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(19),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(19)
    );
  mac_control_rxfifowerr_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(14),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(14)
    );
  mac_control_rxphyerr_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(16),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(16)
    );
  mac_control_rxphyerr_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(18),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(18)
    );
  mac_control_rxphyerr_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(25),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(25)
    );
  mac_control_rxphyerr_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(20),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(20)
    );
  mac_control_rxphyerr_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(23),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(23)
    );
  mac_control_rxphyerr_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(27),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(27)
    );
  tx_fifocheck_diff_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_4_FFX_RST,
      O => tx_fifocheck_diff(4)
    );
  tx_fifocheck_diff_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_4_FFX_RST
    );
  tx_fifocheck_diff_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_6_FFX_RST,
      O => tx_fifocheck_diff(6)
    );
  tx_fifocheck_diff_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_6_FFX_RST
    );
  tx_fifocheck_diff_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_8_FFX_RST,
      O => tx_fifocheck_diff(8)
    );
  tx_fifocheck_diff_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_8_FFX_RST
    );
  mac_control_rxfifowerr_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(16),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(16)
    );
  mac_control_rxfifowerr_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(23),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(23)
    );
  mac_control_rxfifowerr_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(18),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(18)
    );
  mac_control_rxfifowerr_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(21),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(21)
    );
  mac_control_rxfifowerr_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(25),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(25)
    );
  mac_control_rxfifowerr_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(20),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(20)
    );
  tx_output_bcnt_40_1698 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_173,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_39_FFY_RST,
      O => tx_output_bcnt_40
    );
  tx_output_bcnt_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_39_FFY_RST
    );
  tx_output_bcnt_39_1699 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_172,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_39_FFX_RST,
      O => tx_output_bcnt_39
    );
  tx_output_bcnt_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_39_FFX_RST
    );
  tx_output_bcnt_42_1700 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_175,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_41_FFY_RST,
      O => tx_output_bcnt_42
    );
  tx_output_bcnt_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_41_FFY_RST
    );
  tx_output_bcnt_46_1701 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_179,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_45_FFY_RST,
      O => tx_output_bcnt_46
    );
  tx_output_bcnt_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_45_FFY_RST
    );
  tx_output_bcnt_41_1702 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_174,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_41_FFX_RST,
      O => tx_output_bcnt_41
    );
  tx_output_bcnt_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_41_FFX_RST
    );
  tx_output_bcnt_44_1703 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_177,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_43_FFY_RST,
      O => tx_output_bcnt_44
    );
  tx_output_bcnt_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_43_FFY_RST
    );
  mac_control_rxphyerr_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(28),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(28)
    );
  mac_control_rxphyerr_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt_n0000(30),
      CE => rxphyerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxphyerr_rst,
      O => mac_control_rxphyerr_cnt(30)
    );
  mac_control_rxfifowerr_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_Madd_n0000_inst_lut2_16,
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(0)
    );
  mac_control_rxfifowerr_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(5),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(5)
    );
  mac_control_rxfifowerr_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(7),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(7)
    );
  mac_control_rxfifowerr_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(2),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(2)
    );
  mac_control_rxfifowerr_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(28),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(28)
    );
  mac_control_rxfifowerr_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxfifowerr_cnt_n0000(30),
      CE => rxfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxfifowerr_rst,
      O => mac_control_rxfifowerr_cnt(30)
    );
  mac_control_txfifowerr_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(1),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(1)
    );
  mac_control_txfifowerr_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(5),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(5)
    );
  mac_control_txfifowerr_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_Madd_n0000_inst_lut2_16,
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(0)
    );
  mac_control_txfifowerr_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(3),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(3)
    );
  mac_control_txfifowerr_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(20),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(20)
    );
  mac_control_txfifowerr_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(22),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(22)
    );
  mac_control_txfifowerr_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(25),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(25)
    );
  mac_control_txfifowerr_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(29),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(29)
    );
  mac_control_txfifowerr_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(24),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(24)
    );
  mac_control_txfifowerr_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(27),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(27)
    );
  rx_fifocheck_diff_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_8_FFX_RST,
      O => rx_fifocheck_diff(8)
    );
  rx_fifocheck_diff_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_8_FFX_RST
    );
  rx_fifocheck_diff_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_10_FFX_RST,
      O => rx_fifocheck_diff(10)
    );
  rx_fifocheck_diff_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_10_FFX_RST
    );
  rx_fifocheck_diff_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_12_FFY_RST,
      O => rx_fifocheck_diff(13)
    );
  rx_fifocheck_diff_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_12_FFY_RST
    );
  tx_fifocheck_diff_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_0_FFY_RST,
      O => tx_fifocheck_diff(1)
    );
  tx_fifocheck_diff_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_0_FFY_RST
    );
  rx_fifocheck_diff_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_12_FFX_RST,
      O => rx_fifocheck_diff(12)
    );
  rx_fifocheck_diff_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_12_FFX_RST
    );
  rx_fifocheck_diff_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_14_FFY_RST,
      O => rx_fifocheck_diff(15)
    );
  rx_fifocheck_diff_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_14_FFY_RST
    );
  mac_control_txf_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(26),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(26)
    );
  mac_control_txf_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(28),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(28)
    );
  rx_output_macnt_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_97,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_1_FFY_RST,
      O => addr3ext(2)
    );
  addr3ext_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_1_FFY_RST
    );
  mac_control_txf_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(30),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(30)
    );
  rx_output_macnt_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_95,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_0_FFY_RST,
      O => addr3ext(0)
    );
  addr3ext_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_0_FFY_RST
    );
  mac_control_txfifowerr_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(26),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(26)
    );
  mac_control_txfifowerr_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(28),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(28)
    );
  mac_control_txfifowerr_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(31),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(31)
    );
  mac_control_txfifowerr_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt_n0000(30),
      CE => txfifowerr,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txfifowerr_rst,
      O => mac_control_txfifowerr_cnt(30)
    );
  mac_control_phyrstcnt_117_1704 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_264,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_117_FFX_RST,
      O => mac_control_phyrstcnt_117
    );
  mac_control_phyrstcnt_117_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_117_FFX_RST
    );
  mac_control_phyrstcnt_119_1705 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_266,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_119_FFX_RST,
      O => mac_control_phyrstcnt_119
    );
  mac_control_phyrstcnt_119_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_119_FFX_RST
    );
  mac_control_phyrstcnt_122_1706 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_269,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_121_FFY_RST,
      O => mac_control_phyrstcnt_122
    );
  mac_control_phyrstcnt_121_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_121_FFY_RST
    );
  mac_control_phyrstcnt_126_1707 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_273,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_125_FFY_RST,
      O => mac_control_phyrstcnt_126
    );
  mac_control_phyrstcnt_125_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_125_FFY_RST
    );
  mac_control_phyrstcnt_121_1708 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_268,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_121_FFX_RST,
      O => mac_control_phyrstcnt_121
    );
  mac_control_phyrstcnt_121_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_121_FFX_RST
    );
  mac_control_phyrstcnt_124_1709 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_271,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_123_FFY_RST,
      O => mac_control_phyrstcnt_124
    );
  mac_control_phyrstcnt_123_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_123_FFY_RST
    );
  rx_output_bp_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(10),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_10_FFX_RST,
      O => rx_output_bp(10)
    );
  rx_output_bp_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_10_FFX_RST
    );
  rx_output_bp_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(12),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_12_FFX_RST,
      O => rx_output_bp(12)
    );
  rx_output_bp_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_12_FFX_RST
    );
  rx_output_bp_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(15),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_14_FFY_RST,
      O => rx_output_bp(15)
    );
  rx_output_bp_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_14_FFY_RST
    );
  rx_output_bp_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(14),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_14_FFX_RST,
      O => rx_output_bp(14)
    );
  rx_output_bp_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_14_FFX_RST
    );
  tx_output_bcnt_38_1710 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_171,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_38_FFY_RST,
      O => tx_output_bcnt_38
    );
  tx_output_bcnt_38_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_38_FFY_RST
    );
  tx_output_bcnt_43_1711 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_176,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_43_FFX_RST,
      O => tx_output_bcnt_43
    );
  tx_output_bcnt_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_43_FFX_RST
    );
  tx_output_bcnt_45_1712 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_178,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_45_FFX_RST,
      O => tx_output_bcnt_45
    );
  tx_output_bcnt_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_45_FFX_RST
    );
  tx_output_bcnt_48_1713 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_181,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_47_FFY_RST,
      O => tx_output_bcnt_48
    );
  tx_output_bcnt_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_47_FFY_RST
    );
  tx_output_bcnt_52_1714 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_185,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_51_FFY_RST,
      O => tx_output_bcnt_52
    );
  tx_output_bcnt_51_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_51_FFY_RST
    );
  tx_output_bcnt_47_1715 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_180,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_47_FFX_RST,
      O => tx_output_bcnt_47
    );
  tx_output_bcnt_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_47_FFX_RST
    );
  tx_output_bcnt_50_1716 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_183,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_49_FFY_RST,
      O => tx_output_bcnt_50
    );
  tx_output_bcnt_49_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_49_FFY_RST
    );
  rx_output_bp_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(4),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_4_FFX_RST,
      O => rx_output_bp(4)
    );
  rx_output_bp_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_4_FFX_RST
    );
  rx_output_bp_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(6),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_6_FFX_RST,
      O => rx_output_bp(6)
    );
  rx_output_bp_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_6_FFX_RST
    );
  rx_output_bp_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(9),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_8_FFY_RST,
      O => rx_output_bp(9)
    );
  rx_output_bp_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_8_FFY_RST
    );
  rx_output_bp_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(13),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_12_FFY_RST,
      O => rx_output_bp(13)
    );
  rx_output_bp_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_12_FFY_RST
    );
  rx_output_bp_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(8),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_8_FFX_RST,
      O => rx_output_bp(8)
    );
  rx_output_bp_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_8_FFX_RST
    );
  rx_output_bp_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lbp(11),
      CE => rx_output_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_bp_10_FFY_RST,
      O => rx_output_bp(11)
    );
  rx_output_bp_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_bp_10_FFY_RST
    );
  tx_output_bcnt_49_1717 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_182,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_49_FFX_RST,
      O => tx_output_bcnt_49
    );
  tx_output_bcnt_49_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_49_FFX_RST
    );
  tx_output_bcnt_51_1718 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_bcnt_inst_sum_184,
      CE => tx_output_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bcnt_51_FFX_RST,
      O => tx_output_bcnt_51
    );
  tx_output_bcnt_51_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bcnt_51_FFX_RST
    );
  rx_output_macnt_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_102,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_7_FFX_RST,
      O => addr3ext(7)
    );
  addr3ext_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_7_FFX_RST
    );
  rx_output_macnt_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_105,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_9_FFY_RST,
      O => addr3ext(10)
    );
  addr3ext_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_9_FFY_RST
    );
  rx_output_macnt_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_104,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_9_FFX_RST,
      O => addr3ext(9)
    );
  addr3ext_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_9_FFX_RST
    );
  rx_output_macnt_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_107,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_11_FFY_RST,
      O => addr3ext(12)
    );
  addr3ext_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_11_FFY_RST
    );
  rx_output_macnt_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_109,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_13_FFY_RST,
      O => addr3ext(14)
    );
  addr3ext_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_13_FFY_RST
    );
  rx_output_macnt_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_106,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_11_FFX_RST,
      O => addr3ext(11)
    );
  addr3ext_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_11_FFX_RST
    );
  rx_fifocheck_diff_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_2_FFX_RST,
      O => rx_fifocheck_diff(2)
    );
  rx_fifocheck_diff_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_2_FFX_RST
    );
  rx_fifocheck_diff_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_4_FFX_RST,
      O => rx_fifocheck_diff(4)
    );
  rx_fifocheck_diff_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_4_FFX_RST
    );
  rx_fifocheck_diff_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_6_FFY_RST,
      O => rx_fifocheck_diff(7)
    );
  rx_fifocheck_diff_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_6_FFY_RST
    );
  rx_fifocheck_diff_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_10_FFY_RST,
      O => rx_fifocheck_diff(11)
    );
  rx_fifocheck_diff_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_10_FFY_RST
    );
  rx_fifocheck_diff_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_6_FFX_RST,
      O => rx_fifocheck_diff(6)
    );
  rx_fifocheck_diff_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_6_FFX_RST
    );
  rx_fifocheck_diff_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_8_FFY_RST,
      O => rx_fifocheck_diff(9)
    );
  rx_fifocheck_diff_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_8_FFY_RST
    );
  rx_output_fifo_BU65 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1908,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N13_FFX_RST,
      O => rx_output_fifo_N13
    );
  rx_output_fifo_N13_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N13_FFX_RST
    );
  rx_output_fifo_BU77 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1910,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N11_FFX_RST,
      O => rx_output_fifo_N11
    );
  rx_output_fifo_N11_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N11_FFX_RST
    );
  rx_fifocheck_diff_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_fifocheck_n0001(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_diff_14_FFX_RST,
      O => rx_fifocheck_diff(14)
    );
  rx_fifocheck_diff_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_diff_14_FFX_RST
    );
  tx_fifocheck_diff_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_0_FFX_RST,
      O => tx_fifocheck_diff(0)
    );
  tx_fifocheck_diff_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_0_FFX_RST
    );
  tx_fifocheck_diff_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_fifocheck_n0001(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_diff_2_FFX_RST,
      O => tx_fifocheck_diff(2)
    );
  tx_fifocheck_diff_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_diff_2_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_34_1719 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_167,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_33_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_34
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_33_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_32_1720 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_165,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_32_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_32
    );
  mac_control_PHY_status_MII_Interface_mdccnt_32_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_32_FFY_RST
    );
  mac_control_phyrstcnt_129_1721 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_276,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_129_FFX_RST,
      O => mac_control_phyrstcnt_129
    );
  mac_control_phyrstcnt_129_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_129_FFX_RST
    );
  mac_control_phyrstcnt_131_1722 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_278,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_131_FFX_RST,
      O => mac_control_phyrstcnt_131
    );
  mac_control_phyrstcnt_131_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_131_FFX_RST
    );
  mac_control_phyrstcnt_134_1723 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_281,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_133_FFY_RST,
      O => mac_control_phyrstcnt_134
    );
  mac_control_phyrstcnt_133_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_133_FFY_RST
    );
  mac_control_phyrstcnt_133_1724 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_280,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_133_FFX_RST,
      O => mac_control_phyrstcnt_133
    );
  mac_control_phyrstcnt_133_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_133_FFX_RST
    );
  mac_control_phyrstcnt_136_1725 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_283,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_135_FFY_RST,
      O => mac_control_phyrstcnt_136
    );
  mac_control_phyrstcnt_135_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_135_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_1726 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_166,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_33_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_33
    );
  mac_control_PHY_status_MII_Interface_mdccnt_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_33_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_36_1727 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_169,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_35_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_36
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_35_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_1728 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_mdccnt_inst_sum_168,
      CE => mac_control_PHY_status_MII_Interface_n0013,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_mdccnt_35_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_mdccnt_35
    );
  mac_control_PHY_status_MII_Interface_mdccnt_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_mdccnt_35_FFX_RST
    );
  mac_control_ledtx_cnt_143_1729 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_290,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_143_FFX_RST,
      O => mac_control_ledtx_cnt_143
    );
  mac_control_ledtx_cnt_143_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_143_FFX_RST
    );
  mac_control_ledtx_cnt_146_1730 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_293,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_145_FFY_RST,
      O => mac_control_ledtx_cnt_146
    );
  mac_control_ledtx_cnt_145_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_145_FFY_RST
    );
  mac_control_ledtx_cnt_150_1731 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_297,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_149_FFY_RST,
      O => mac_control_ledtx_cnt_150
    );
  mac_control_ledtx_cnt_149_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_149_FFY_RST
    );
  mac_control_ledtx_cnt_145_1732 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_292,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_145_FFX_RST,
      O => mac_control_ledtx_cnt_145
    );
  mac_control_ledtx_cnt_145_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_145_FFX_RST
    );
  mac_control_ledtx_cnt_148_1733 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_ledtx_cnt_inst_sum_295,
      CE => mac_control_n0037,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_cnt_147_FFY_RST,
      O => mac_control_ledtx_cnt_148
    );
  mac_control_ledtx_cnt_147_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_cnt_147_FFY_RST
    );
  rx_output_fifo_BU41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1904,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N17_FFX_RST,
      O => rx_output_fifo_N17
    );
  rx_output_fifo_N17_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N17_FFX_RST
    );
  rx_output_fifo_BU59 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1907,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N15_FFY_RST,
      O => rx_output_fifo_N14
    );
  rx_output_fifo_N15_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N15_FFY_RST
    );
  rx_output_fifo_BU53 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1906,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N15_FFX_RST,
      O => rx_output_fifo_N15
    );
  rx_output_fifo_N15_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N15_FFX_RST
    );
  rx_output_fifo_BU71 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1909,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N13_FFY_RST,
      O => rx_output_fifo_N12
    );
  rx_output_fifo_N13_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N13_FFY_RST
    );
  rx_output_fifo_BU82 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1911,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N11_FFY_RST,
      O => rx_output_fifo_N10
    );
  rx_output_fifo_N11_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N11_FFY_RST
    );
  mac_control_txf_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(8),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(8)
    );
  mac_control_txf_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(10),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(10)
    );
  mac_control_txf_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(17),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(17)
    );
  mac_control_txf_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(12),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(12)
    );
  mac_control_txf_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(15),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(15)
    );
  mac_control_txf_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(19),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(19)
    );
  mac_control_txf_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(1),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(1)
    );
  mac_control_txf_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(7),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(7)
    );
  mac_control_txf_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_Madd_n0000_inst_lut2_16,
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(0)
    );
  mac_control_txf_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(5),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(5)
    );
  mac_control_phyrstcnt_139_1734 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_286,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_139_FFX_RST,
      O => mac_control_phyrstcnt_139
    );
  mac_control_phyrstcnt_139_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_139_FFX_RST
    );
  rx_input_memio_macnt_70_1735 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_219,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_70_FFY_RST,
      O => rx_input_memio_macnt_70
    );
  rx_input_memio_macnt_70_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_70_FFY_RST
    );
  rx_input_memio_macnt_78_1736 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_227,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_77_FFY_RST,
      O => rx_input_memio_macnt_78
    );
  rx_input_memio_macnt_77_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_77_FFY_RST
    );
  rx_input_memio_macnt_71_1737 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_220,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_71_FFX_RST,
      O => rx_input_memio_macnt_71
    );
  rx_input_memio_macnt_71_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_71_FFX_RST
    );
  rx_input_memio_macnt_74_1738 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_223,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_73_FFY_RST,
      O => rx_input_memio_macnt_74
    );
  rx_input_memio_macnt_73_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_73_FFY_RST
    );
  rx_input_memio_macnt_76_1739 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_225,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_75_FFY_RST,
      O => rx_input_memio_macnt_76
    );
  rx_input_memio_macnt_75_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_75_FFY_RST
    );
  mac_control_txf_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(20),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(20)
    );
  mac_control_txf_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(22),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(22)
    );
  mac_control_txf_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(29),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(29)
    );
  mac_control_txf_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(24),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(24)
    );
  mac_control_txf_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(27),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(27)
    );
  mac_control_txf_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(31),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(31)
    );
  tx_input_addr_17_1740 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_128,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_17_FFX_RST,
      O => tx_input_addr_17
    );
  tx_input_addr_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_17_FFX_RST
    );
  tx_input_addr_20_1741 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_131,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_19_FFY_RST,
      O => tx_input_addr_20
    );
  tx_input_addr_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_19_FFY_RST
    );
  tx_input_addr_19_1742 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_130,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_19_FFX_RST,
      O => tx_input_addr_19
    );
  tx_input_addr_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_19_FFX_RST
    );
  tx_input_addr_22_1743 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_133,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_21_FFY_RST,
      O => tx_input_addr_22
    );
  tx_input_addr_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_21_FFY_RST
    );
  tx_input_addr_24_1744 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_135,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_23_FFY_RST,
      O => tx_input_addr_24
    );
  tx_input_addr_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_23_FFY_RST
    );
  mac_control_txf_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(14),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(14)
    );
  mac_control_txf_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(16),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(16)
    );
  mac_control_txf_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(23),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(23)
    );
  mac_control_txf_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(18),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(18)
    );
  mac_control_txf_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(21),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(21)
    );
  mac_control_txf_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(25),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(25)
    );
  mac_control_txf_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(2),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(2)
    );
  mac_control_txf_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(4),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(4)
    );
  mac_control_txf_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(11),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(11)
    );
  mac_control_txf_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(6),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(6)
    );
  mac_control_txf_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(9),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(9)
    );
  mac_control_txf_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt_n0000(13),
      CE => txf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_txf_rst,
      O => mac_control_txf_cnt(13)
    );
  mac_control_phyrstcnt_112_1745 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_259,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_111_FFY_RST,
      O => mac_control_phyrstcnt_112
    );
  mac_control_phyrstcnt_111_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_111_FFY_RST
    );
  mac_control_phyrstcnt_110_1746 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_257,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_110_FFY_RST,
      O => mac_control_phyrstcnt_110
    );
  mac_control_phyrstcnt_110_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_110_FFY_RST
    );
  mac_control_phyrstcnt_114_1747 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_261,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_113_FFY_RST,
      O => mac_control_phyrstcnt_114
    );
  mac_control_phyrstcnt_113_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_113_FFY_RST
    );
  rx_output_macnt_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_96,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_1_FFX_RST,
      O => addr3ext(1)
    );
  addr3ext_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_1_FFX_RST
    );
  rx_output_macnt_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_99,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_3_FFY_RST,
      O => addr3ext(4)
    );
  addr3ext_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_3_FFY_RST
    );
  rx_output_macnt_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_98,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_3_FFX_RST,
      O => addr3ext(3)
    );
  addr3ext_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_3_FFX_RST
    );
  rx_output_macnt_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_101,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_5_FFY_RST,
      O => addr3ext(6)
    );
  addr3ext_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_5_FFY_RST
    );
  rx_output_macnt_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_103,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_7_FFY_RST,
      O => addr3ext(8)
    );
  addr3ext_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_7_FFY_RST
    );
  rx_output_macnt_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_100,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_5_FFX_RST,
      O => addr3ext(5)
    );
  addr3ext_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_5_FFX_RST
    );
  mac_control_phyrstcnt_123_1748 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_270,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_123_FFX_RST,
      O => mac_control_phyrstcnt_123
    );
  mac_control_phyrstcnt_123_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_123_FFX_RST
    );
  mac_control_phyrstcnt_125_1749 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_272,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_125_FFX_RST,
      O => mac_control_phyrstcnt_125
    );
  mac_control_phyrstcnt_125_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_125_FFX_RST
    );
  mac_control_phyrstcnt_128_1750 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_275,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_127_FFY_RST,
      O => mac_control_phyrstcnt_128
    );
  mac_control_phyrstcnt_127_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_127_FFY_RST
    );
  mac_control_phyrstcnt_132_1751 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_279,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_131_FFY_RST,
      O => mac_control_phyrstcnt_132
    );
  mac_control_phyrstcnt_131_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_131_FFY_RST
    );
  mac_control_phyrstcnt_127_1752 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_274,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_127_FFX_RST,
      O => mac_control_phyrstcnt_127
    );
  mac_control_phyrstcnt_127_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_127_FFX_RST
    );
  mac_control_phyrstcnt_130_1753 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_277,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_129_FFY_RST,
      O => mac_control_phyrstcnt_130
    );
  mac_control_phyrstcnt_129_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_129_FFY_RST
    );
  rx_input_memio_bcntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(1),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_0_FFY_RST,
      O => rx_input_memio_bcntl(1)
    );
  rx_input_memio_bcntl_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_0_FFY_RST
    );
  rx_output_macnt_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_108,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_13_FFX_RST,
      O => addr3ext(13)
    );
  addr3ext_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_13_FFX_RST
    );
  rx_output_macnt_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_macnt_inst_sum_110,
      CE => rx_output_n0043,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr3ext_15_FFX_RST,
      O => addr3ext(15)
    );
  addr3ext_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => addr3ext_15_FFX_RST
    );
  mac_control_phyrstcnt_135_1754 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_282,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_135_FFX_RST,
      O => mac_control_phyrstcnt_135
    );
  mac_control_phyrstcnt_135_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_135_FFX_RST
    );
  mac_control_phyrstcnt_138_1755 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_285,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_137_FFY_RST,
      O => mac_control_phyrstcnt_138
    );
  mac_control_phyrstcnt_137_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_137_FFY_RST
    );
  mac_control_phyrstcnt_137_1756 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_284,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_137_FFX_RST,
      O => mac_control_phyrstcnt_137
    );
  mac_control_phyrstcnt_137_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_137_FFX_RST
    );
  mac_control_phyrstcnt_140_1757 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_287,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_139_FFY_RST,
      O => mac_control_phyrstcnt_140
    );
  mac_control_phyrstcnt_139_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_139_FFY_RST
    );
  mac_control_phyrstcnt_141_1758 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_288,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_phyrstcnt_141_FFX_RST,
      O => mac_control_phyrstcnt_141
    );
  mac_control_phyrstcnt_141_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_141_FFX_RST
    );
  mac_control_phyrstcnt_111_1759 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_258,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_111_FFX_RST,
      O => mac_control_phyrstcnt_111
    );
  mac_control_phyrstcnt_111_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_111_FFX_RST
    );
  mac_control_phyrstcnt_113_1760 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_260,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_113_FFX_RST,
      O => mac_control_phyrstcnt_113
    );
  mac_control_phyrstcnt_113_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_113_FFX_RST
    );
  mac_control_phyrstcnt_116_1761 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_263,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_115_FFY_RST,
      O => mac_control_phyrstcnt_116
    );
  mac_control_phyrstcnt_115_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_115_FFY_RST
    );
  mac_control_phyrstcnt_120_1762 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_267,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_119_FFY_RST,
      O => mac_control_phyrstcnt_120
    );
  mac_control_phyrstcnt_119_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_119_FFY_RST
    );
  mac_control_phyrstcnt_115_1763 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_262,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_115_FFX_RST,
      O => mac_control_phyrstcnt_115
    );
  mac_control_phyrstcnt_115_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_115_FFX_RST
    );
  mac_control_phyrstcnt_118_1764 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyrstcnt_inst_sum_265,
      CE => mac_control_n0032,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyrstcnt_117_FFY_RST,
      O => mac_control_phyrstcnt_118
    );
  mac_control_phyrstcnt_117_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyrstcnt_117_FFY_RST
    );
  rx_input_memio_macnt_73_1765 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_222,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_73_FFX_RST,
      O => rx_input_memio_macnt_73
    );
  rx_input_memio_macnt_73_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_73_FFX_RST
    );
  rx_input_memio_macnt_84_1766 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_233,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_83_FFY_RST,
      O => rx_input_memio_macnt_84
    );
  rx_input_memio_macnt_83_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_83_FFY_RST
    );
  rx_input_memio_macnt_75_1767 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_224,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_75_FFX_RST,
      O => rx_input_memio_macnt_75
    );
  rx_input_memio_macnt_75_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_75_FFX_RST
    );
  rx_input_memio_macnt_77_1768 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_226,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_77_FFX_RST,
      O => rx_input_memio_macnt_77
    );
  rx_input_memio_macnt_77_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_77_FFX_RST
    );
  rx_input_memio_macnt_80_1769 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_229,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_79_FFY_RST,
      O => rx_input_memio_macnt_80
    );
  rx_input_memio_macnt_79_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_79_FFY_RST
    );
  rx_input_memio_macnt_82_1770 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_231,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_81_FFY_RST,
      O => rx_input_memio_macnt_82
    );
  rx_input_memio_macnt_81_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_81_FFY_RST
    );
  mac_control_rxf_cnt_14 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(14),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(14)
    );
  mac_control_rxf_cnt_16 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(16),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(16)
    );
  mac_control_rxf_cnt_23 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(23),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(23)
    );
  mac_control_rxf_cnt_18 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(18),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(18)
    );
  mac_control_rxf_cnt_21 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(21),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(21)
    );
  mac_control_rxf_cnt_25 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(25),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(25)
    );
  rx_input_memio_bcntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(6),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_6_FFX_RST,
      O => rx_input_memio_bcntl(6)
    );
  rx_input_memio_bcntl_6_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_6_FFX_RST
    );
  rx_input_memio_bcntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(8),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_8_FFX_RST,
      O => rx_input_memio_bcntl(8)
    );
  rx_input_memio_bcntl_8_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_8_FFX_RST
    );
  tx_input_addr_21_1771 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_132,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_21_FFX_RST,
      O => tx_input_addr_21
    );
  tx_input_addr_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_21_FFX_RST
    );
  tx_input_addr_23_1772 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_134,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_23_FFX_RST,
      O => tx_input_addr_23
    );
  tx_input_addr_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_23_FFX_RST
    );
  tx_input_addr_26_1773 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_137,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_25_FFY_RST,
      O => tx_input_addr_26
    );
  tx_input_addr_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_25_FFY_RST
    );
  tx_input_addr_25_1774 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_136,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_25_FFX_RST,
      O => tx_input_addr_25
    );
  tx_input_addr_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_25_FFX_RST
    );
  tx_input_addr_28_1775 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_139,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_27_FFY_RST,
      O => tx_input_addr_28
    );
  tx_input_addr_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_27_FFY_RST
    );
  tx_input_addr_30_1776 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_141,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_29_FFY_RST,
      O => tx_input_addr_30
    );
  tx_input_addr_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_29_FFY_RST
    );
  mac_control_txf_rst_1777 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0046,
      CE => mac_control_txf_rst_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_rst_FFX_RST,
      O => mac_control_txf_rst
    );
  mac_control_txf_rst_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_rst_FFX_RST
    );
  rx_input_memio_addrchk_cs_FFd4_1778 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd4_FFX_RST,
      O => rx_input_memio_addrchk_cs_FFd4
    );
  rx_input_memio_addrchk_cs_FFd4_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd4_FFX_RST
    );
  rx_input_memio_cs_FFd9_1779 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd9_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd10_FFY_RST,
      O => rx_input_memio_cs_FFd9
    );
  rx_input_memio_cs_FFd10_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd10_FFY_RST
    );
  rx_input_memio_cs_FFd10_1780 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd10_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd10_FFX_RST,
      O => rx_input_memio_cs_FFd10
    );
  rx_input_memio_cs_FFd10_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd10_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(0),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_1_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(0)
    );
  mac_control_PHY_status_MII_Interface_statecnt_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_1_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(2),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_3_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(2)
    );
  mac_control_PHY_status_MII_Interface_statecnt_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_3_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(1),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_1_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(1)
    );
  mac_control_PHY_status_MII_Interface_statecnt_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_1_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(3),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_3_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(3)
    );
  mac_control_PHY_status_MII_Interface_statecnt_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_3_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(4),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_5_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(4)
    );
  mac_control_PHY_status_MII_Interface_statecnt_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_5_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_statecnt_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_n0014(5),
      CE => mac_control_PHY_status_MII_Interface_n0010,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_statecnt_5_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_statecnt(5)
    );
  mac_control_PHY_status_MII_Interface_statecnt_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_statecnt_5_FFX_RST
    );
  rx_input_memio_MA_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_1_FFY_RST,
      O => addr1ext(0)
    );
  addr1ext_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_1_FFY_RST
    );
  rx_input_memio_bcntl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(0),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_0_FFX_RST,
      O => rx_input_memio_bcntl(0)
    );
  rx_input_memio_bcntl_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_0_FFX_RST
    );
  rx_input_memio_bcntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(2),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_2_FFX_RST,
      O => rx_input_memio_bcntl(2)
    );
  rx_input_memio_bcntl_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_2_FFX_RST
    );
  rx_input_memio_bcntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(4),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_4_FFX_RST,
      O => rx_input_memio_bcntl(4)
    );
  rx_input_memio_bcntl_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_4_FFX_RST
    );
  mac_control_rxf_cnt_20 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(20),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(20)
    );
  mac_control_rxf_cnt_22 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(22),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(22)
    );
  mac_control_rxf_cnt_29 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(29),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(29)
    );
  mac_control_rxf_cnt_24 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(24),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(24)
    );
  mac_control_rxf_cnt_27 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(27),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(27)
    );
  mac_control_rxf_cnt_31 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(31),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(31)
    );
  tx_input_addr_27_1781 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_138,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_27_FFX_RST,
      O => tx_input_addr_27
    );
  tx_input_addr_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_27_FFX_RST
    );
  mac_control_rxf_cnt_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(1),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(1)
    );
  tx_input_addr_29_1782 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_140,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_29_FFX_RST,
      O => tx_input_addr_29
    );
  tx_input_addr_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_29_FFX_RST
    );
  tx_input_addr_31_1783 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_142,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_31_FFX_RST,
      O => tx_input_addr_31
    );
  tx_input_addr_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_31_FFX_RST
    );
  mac_control_rxf_cnt_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(3),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(3)
    );
  mac_control_rxf_cnt_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(7),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(7)
    );
  mac_control_rxf_cnt_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_Madd_n0000_inst_lut2_16,
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(0)
    );
  mac_control_rxf_cnt_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(5),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(5)
    );
  rx_input_memio_bcntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(10),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_10_FFX_RST,
      O => rx_input_memio_bcntl(10)
    );
  rx_input_memio_bcntl_10_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_10_FFX_RST
    );
  rx_input_memio_bcntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(12),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_12_FFX_RST,
      O => rx_input_memio_bcntl(12)
    );
  rx_input_memio_bcntl_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_12_FFX_RST
    );
  tx_input_addr_18_1784 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_inst_sum_129,
      CE => tx_input_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_addr_17_FFY_RST,
      O => tx_input_addr_18
    );
  tx_input_addr_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_addr_17_FFY_RST
    );
  rx_input_memio_bcntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0042(14),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcntl_14_FFX_RST,
      O => rx_input_memio_bcntl(14)
    );
  rx_input_memio_bcntl_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bcntl_14_FFX_RST
    );
  mac_control_rxf_cnt_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(2),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(2)
    );
  mac_control_rxf_cnt_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(4),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(4)
    );
  mac_control_rxf_cnt_11 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(11),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(11)
    );
  mac_control_rxf_cnt_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(6),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(6)
    );
  mac_control_rxf_cnt_9 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(9),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(9)
    );
  mac_control_rxf_cnt_13 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(13),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(13)
    );
  rx_output_fifo_BU226 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2836,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N5_FFX_RST,
      O => rx_output_fifo_N5
    );
  rx_output_fifo_N5_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N5_FFX_RST
    );
  rx_output_fifo_BU238 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2838,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N3_FFX_RST,
      O => rx_output_fifo_N3
    );
  rx_output_fifo_N3_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N3_FFX_RST
    );
  rx_output_fifo_BU176 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N2580,
      CE => rx_output_fifo_N2579,
      CLK => clkio,
      SET => rx_output_fifo_empty_FFX_SET,
      RST => GND,
      O => rx_output_fifo_empty
    );
  rx_output_fifo_empty_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_empty_FFX_SET
    );
  rx_input_fifo_control_INVALID : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(9),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_endf_FFY_RST,
      O => rx_input_invalid
    );
  rx_input_endf_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_endf_FFY_RST
    );
  tx_output_crcl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_15_1_O,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_15_FFX_RST,
      O => tx_output_crcl(15)
    );
  tx_output_crcl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_15_FFX_RST
    );
  tx_output_crcl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_5_1_O,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_15_FFY_RST,
      O => tx_output_crcl(5)
    );
  tx_output_crcl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_15_FFY_RST
    );
  rx_input_fifo_control_ENDF : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_ldata(8),
      CE => rx_input_fifo_control_n0008,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_endf_FFX_RST,
      O => rx_input_endf
    );
  rx_input_endf_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_endf_FFX_RST
    );
  rx_input_memio_crcl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_5_1_O,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_22_FFY_RST,
      O => rx_input_memio_crcl(5)
    );
  rx_input_memio_crcl_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_22_FFY_RST
    );
  rx_input_memio_crcl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_22_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_22_FFX_RST,
      O => rx_input_memio_crcl(22)
    );
  rx_input_memio_crcl_22_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_22_FFX_RST
    );
  rx_output_lenr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_10_O,
      CE => rx_output_lenr_10_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_10_FFY_RST,
      O => rx_output_lenr(10)
    );
  rx_output_lenr_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_10_FFY_RST
    );
  mac_control_rxf_cnt_8 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(8),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(8)
    );
  mac_control_rxf_cnt_10 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(10),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(10)
    );
  mac_control_rxf_cnt_17 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(17),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(17)
    );
  mac_control_rxf_cnt_12 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(12),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(12)
    );
  mac_control_rxf_cnt_15 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(15),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(15)
    );
  mac_control_rxf_cnt_19 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(19),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(19)
    );
  rx_input_memio_crcl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_15_1_O,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_15_FFX_RST,
      O => rx_input_memio_crcl(15)
    );
  rx_input_memio_crcl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_15_FFX_RST
    );
  rx_input_memio_crcl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_31_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_31_FFX_RST,
      O => rx_input_memio_crcl(31)
    );
  rx_input_memio_crcl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_31_FFX_RST
    );
  rx_input_memio_cs_FFd15_1785 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd15_In7_O,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd15_FFY_RST,
      O => rx_input_memio_cs_FFd15
    );
  rx_input_memio_cs_FFd15_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd15_FFY_RST
    );
  rx_input_memio_menl_1786 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_menl_GROM,
      CE => rx_input_memio_menl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_menl_FFY_RST,
      O => rx_input_memio_menl
    );
  rx_input_memio_menl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_menl_FFY_RST
    );
  mac_control_rxf_cnt_26 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(26),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(26)
    );
  mac_control_rxf_cnt_28 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(28),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(28)
    );
  mac_control_rxf_cnt_30 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt_n0000(30),
      CE => rxf,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => mac_control_rxf_rst,
      O => mac_control_rxf_cnt(30)
    );
  rx_output_lenr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_2_O,
      CE => rx_output_lenr_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_2_FFY_RST,
      O => rx_output_lenr(2)
    );
  rx_output_lenr_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_2_FFY_RST
    );
  rx_output_lenr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_3_O,
      CE => rx_output_lenr_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_3_FFY_RST,
      O => rx_output_lenr(3)
    );
  rx_output_lenr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_3_FFY_RST
    );
  rx_output_lenr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_4_O,
      CE => rx_output_lenr_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_4_FFY_RST,
      O => rx_output_lenr(4)
    );
  rx_output_lenr_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_4_FFY_RST
    );
  rx_output_lenr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_5_O,
      CE => rx_output_lenr_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_5_FFY_RST,
      O => rx_output_lenr(5)
    );
  rx_output_lenr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_5_FFY_RST
    );
  rx_output_lenr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_6_O,
      CE => rx_output_lenr_6_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_6_FFY_RST,
      O => rx_output_lenr(6)
    );
  rx_output_lenr_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_6_FFY_RST
    );
  tx_output_crcenl_1787 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_crcenl_FROM,
      CE => tx_output_crcenl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcenl_FFX_RST,
      O => tx_output_crcenl
    );
  tx_output_crcenl_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcenl_FFX_RST
    );
  mac_control_bitcnt_106_1788 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_253,
      CE => mac_control_n0015,
      CLK => clksl,
      SET => GND,
      RST => mac_control_bitcnt_105_FFY_RST,
      O => mac_control_bitcnt_106
    );
  mac_control_bitcnt_105_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_105_FFY_RST
    );
  mac_control_bitcnt_105_1789 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_252,
      CE => mac_control_n0015,
      CLK => clksl,
      SET => GND,
      RST => mac_control_bitcnt_105_FFX_RST,
      O => mac_control_bitcnt_105
    );
  mac_control_bitcnt_105_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_105_FFX_RST
    );
  mac_control_bitcnt_108_1790 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_255,
      CE => mac_control_n0015,
      CLK => clksl,
      SET => GND,
      RST => mac_control_bitcnt_107_FFY_RST,
      O => mac_control_bitcnt_108
    );
  mac_control_bitcnt_107_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_107_FFY_RST
    );
  rx_input_memio_crcl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_12_1_O,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_15_FFY_RST,
      O => rx_input_memio_crcl(12)
    );
  rx_input_memio_crcl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_15_FFY_RST
    );
  mac_control_bitcnt_107_1791 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_254,
      CE => mac_control_n0015,
      CLK => clksl,
      SET => GND,
      RST => mac_control_bitcnt_107_FFX_RST,
      O => mac_control_bitcnt_107
    );
  mac_control_bitcnt_107_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_107_FFX_RST
    );
  rx_input_memio_MD_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_11_FFX_RST,
      O => d1(11)
    );
  d1_11_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_11_FFX_RST
    );
  rx_input_memio_MD_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(21),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_21_FFX_RST,
      O => d1(21)
    );
  d1_21_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_21_FFX_RST
    );
  rx_input_memio_MD_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(20),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_21_FFY_RST,
      O => d1(20)
    );
  d1_21_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_21_FFY_RST
    );
  rx_input_memio_MD_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_13_FFY_RST,
      O => d1(12)
    );
  d1_13_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_13_FFY_RST
    );
  rx_input_memio_MD_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_13_FFX_RST,
      O => d1(13)
    );
  d1_13_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_13_FFX_RST
    );
  rx_input_memio_MD_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(31),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_31_FFX_RST,
      O => d1(31)
    );
  d1_31_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_31_FFX_RST
    );
  rx_input_memio_MD_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(30),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_31_FFY_RST,
      O => d1(30)
    );
  d1_31_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_31_FFY_RST
    );
  rx_input_memio_MD_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(22),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_23_FFY_RST,
      O => d1(22)
    );
  d1_23_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_23_FFY_RST
    );
  rx_input_memio_MD_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(23),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_23_FFX_RST,
      O => d1(23)
    );
  d1_23_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_23_FFX_RST
    );
  rx_input_memio_MD_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(24),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_25_FFY_RST,
      O => d1(24)
    );
  d1_25_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_25_FFY_RST
    );
  rx_output_fifo_BU208 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2833,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N9_FFY_RST,
      O => rx_output_fifo_N8
    );
  rx_output_fifo_N9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N9_FFY_RST
    );
  rx_output_fifo_BU202 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2832,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N9_FFX_RST,
      O => rx_output_fifo_N9
    );
  rx_output_fifo_N9_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N9_FFX_RST
    );
  rx_output_fifo_BU220 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2835,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N7_FFY_RST,
      O => rx_output_fifo_N6
    );
  rx_output_fifo_N7_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N7_FFY_RST
    );
  rx_output_fifo_BU214 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2834,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N7_FFX_RST,
      O => rx_output_fifo_N7
    );
  rx_output_fifo_N7_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N7_FFX_RST
    );
  rx_output_fifo_BU232 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2837,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N5_FFY_RST,
      O => rx_output_fifo_N4
    );
  rx_output_fifo_N5_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N5_FFY_RST
    );
  rx_output_fifo_BU243 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2839,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N3_FFY_RST,
      O => rx_output_fifo_N2
    );
  rx_output_fifo_N3_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N3_FFY_RST
    );
  rx_output_fifo_BU355 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3618,
      CE => rx_output_fifo_N3617,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_full_FFX_SET,
      RST => GND,
      O => rx_output_fifo_full_0
    );
  rx_output_fifo_full_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_full_FFX_SET
    );
  rx_output_fifo_BU504 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N4755,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_wrcount_0_FFY_RST,
      O => rx_output_fifo_wrcount(1)
    );
  rx_output_fifo_wrcount_0_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_wrcount_0_FFY_RST
    );
  mac_control_bitcnt_104_1792 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_bitcnt_inst_sum_251,
      CE => mac_control_n0015,
      CLK => clksl,
      SET => GND,
      RST => mac_control_bitcnt_104_FFY_RST,
      O => mac_control_bitcnt_104
    );
  mac_control_bitcnt_104_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_bitcnt_104_FFY_RST
    );
  rx_output_fifo_BU498 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N4754,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_wrcount_0_FFX_RST,
      O => rx_output_fifo_wrcount(0)
    );
  rx_output_fifo_wrcount_0_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_wrcount_0_FFX_RST
    );
  rx_output_lenr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_11_O,
      CE => rx_output_lenr_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_11_FFY_RST,
      O => rx_output_lenr(11)
    );
  rx_output_lenr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_11_FFY_RST
    );
  rx_output_lenr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_12_O,
      CE => rx_output_lenr_12_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_12_FFY_RST,
      O => rx_output_lenr(12)
    );
  rx_output_lenr_12_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_12_FFY_RST
    );
  rx_output_lenr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_13_O,
      CE => rx_output_lenr_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_13_FFY_RST,
      O => rx_output_lenr(13)
    );
  rx_output_lenr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_13_FFY_RST
    );
  rx_output_lenr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_14_O,
      CE => rx_output_lenr_14_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_14_FFY_RST,
      O => rx_output_lenr(14)
    );
  rx_output_lenr_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_14_FFY_RST
    );
  rx_output_lenr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_15_O,
      CE => rx_output_lenr_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_15_FFY_RST,
      O => rx_output_lenr(15)
    );
  rx_output_lenr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_15_FFY_RST
    );
  tx_input_cs_FFd6_1793 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd6_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd6_FFX_RST,
      O => tx_input_cs_FFd6
    );
  tx_input_cs_FFd6_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd6_FFX_RST
    );
  tx_input_cs_FFd8_1794 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd8_In1_O,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd8_FFX_RST,
      O => tx_input_cs_FFd8
    );
  tx_input_cs_FFd8_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd8_FFX_RST
    );
  rx_input_fifo_control_cel : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_rd_en_FROM,
      CE => rx_input_fifo_rd_en_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_rd_en_FFX_RST,
      O => rx_input_fifo_rd_en
    );
  rx_input_fifo_rd_en_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_rd_en_FFX_RST
    );
  mac_control_PHY_status_PHYADDRSTATUS : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_n00181_O,
      CE => mac_control_PHY_status_n00171_O,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phyaddr_31_FFY_RST,
      O => mac_control_phyaddr(31)
    );
  mac_control_phyaddr_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_31_FFY_RST
    );
  mac_control_txfifowerr_rst_1795 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0048,
      CE => mac_control_txf_rst_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_rst_FFY_RST,
      O => mac_control_txfifowerr_rst
    );
  mac_control_txf_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_rst_FFY_RST
    );
  rx_input_memio_addrchk_cs_FFd3_1796 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd4_FFY_RST,
      O => rx_input_memio_addrchk_cs_FFd3
    );
  rx_input_memio_addrchk_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd4_FFY_RST
    );
  rx_input_memio_MA_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_3_FFX_RST,
      O => addr1ext(3)
    );
  addr1ext_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_3_FFX_RST
    );
  rx_input_memio_MA_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_1_FFX_RST,
      O => addr1ext(1)
    );
  addr1ext_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_1_FFX_RST
    );
  rx_input_memio_MA_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_3_FFY_RST,
      O => addr1ext(2)
    );
  addr1ext_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => addr1ext_3_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd5_1797 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd5_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_cs_FFd5_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_cs_FFd5
    );
  mac_control_PHY_status_MII_Interface_cs_FFd5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_MII_Interface_cs_FFd5_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd4_1798 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_cs_FFd5_FFY_RST,
      O => mac_control_PHY_status_MII_Interface_cs_FFd4
    );
  mac_control_PHY_status_MII_Interface_cs_FFd5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_MII_Interface_cs_FFd5_FFY_RST
    );
  rx_input_memio_MA_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_5_FFY_RST,
      O => addr1ext(4)
    );
  addr1ext_5_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_5_FFY_RST
    );
  rx_input_memio_MA_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_7_FFX_RST,
      O => addr1ext(7)
    );
  addr1ext_7_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_7_FFX_RST
    );
  rx_input_memio_MA_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_5_FFX_RST,
      O => addr1ext(5)
    );
  addr1ext_5_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_5_FFX_RST
    );
  rx_input_memio_MA_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_7_FFY_RST,
      O => addr1ext(6)
    );
  addr1ext_7_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_7_FFY_RST
    );
  rx_input_memio_MA_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_9_FFY_RST,
      O => addr1ext(8)
    );
  addr1ext_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_9_FFY_RST
    );
  rx_input_memio_MD_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_15_FFY_RST,
      O => d1(0)
    );
  d1_15_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_15_FFY_RST
    );
  tx_input_CNT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(1),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_1_FFX_RST,
      O => tx_input_CNT(1)
    );
  tx_input_CNT_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_1_FFX_RST
    );
  tx_input_CNT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(3),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_3_FFX_RST,
      O => tx_input_CNT(3)
    );
  tx_input_CNT_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_3_FFX_RST
    );
  tx_input_CNT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(5),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_5_FFX_RST,
      O => tx_input_CNT(5)
    );
  tx_input_CNT_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_5_FFX_RST
    );
  tx_input_CNT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(4),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_5_FFY_RST,
      O => tx_input_CNT(4)
    );
  tx_input_CNT_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_5_FFY_RST
    );
  tx_input_CNT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(7),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_7_FFX_RST,
      O => tx_input_CNT(7)
    );
  tx_input_CNT_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_7_FFX_RST
    );
  tx_input_CNT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(6),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_7_FFY_RST,
      O => tx_input_CNT(6)
    );
  tx_input_CNT_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_7_FFY_RST
    );
  tx_input_CNT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(9),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_9_FFX_RST,
      O => tx_input_CNT(9)
    );
  tx_input_CNT_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_9_FFX_RST
    );
  tx_input_CNT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(8),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_9_FFY_RST,
      O => tx_input_CNT(8)
    );
  tx_input_CNT_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_9_FFY_RST
    );
  rx_input_GMII_ENDFIN : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_endfin_GROM,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_endfin_FFY_RST,
      O => rx_input_endfin
    );
  rx_input_endfin_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_endfin_FFY_RST
    );
  rx_output_fifo_BU30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N1835,
      CE => VCC,
      CLK => clkio,
      SET => GND,
      RST => rx_output_invalid_FFY_RST,
      O => rx_output_invalid
    );
  rx_output_invalid_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_invalid_FFY_RST
    );
  rx_input_memio_MA_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_9_FFX_RST,
      O => addr1ext(9)
    );
  addr1ext_9_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_9_FFX_RST
    );
  rx_input_memio_MD_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_15_FFX_RST,
      O => d1(15)
    );
  d1_15_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_15_FFX_RST
    );
  rx_input_memio_MD_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_14_FFX_RST,
      O => d1(14)
    );
  d1_14_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_14_FFX_RST
    );
  rx_input_memio_MD_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_14_FFY_RST,
      O => d1(1)
    );
  d1_14_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_14_FFY_RST
    );
  rx_input_memio_MD_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_3_FFX_RST,
      O => d1(3)
    );
  d1_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_3_FFX_RST
    );
  rx_input_memio_MD_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_3_FFY_RST,
      O => d1(2)
    );
  d1_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_3_FFY_RST
    );
  rx_input_memio_MD_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_5_FFX_RST,
      O => d1(5)
    );
  d1_5_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_5_FFX_RST
    );
  rx_input_memio_MD_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_5_FFY_RST,
      O => d1(4)
    );
  d1_5_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_5_FFY_RST
    );
  rx_input_memio_MD_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_7_FFX_RST,
      O => d1(7)
    );
  d1_7_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_7_FFX_RST
    );
  rx_input_memio_MD_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_7_FFY_RST,
      O => d1(6)
    );
  d1_7_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_7_FFY_RST
    );
  rx_input_memio_MD_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_9_FFY_RST,
      O => d1(8)
    );
  d1_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_9_FFY_RST
    );
  mac_control_rxfifowerr_rst_1799 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0049,
      CE => mac_control_rxfifowerr_rst_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_rst_FFX_RST,
      O => mac_control_rxfifowerr_rst
    );
  mac_control_rxfifowerr_rst_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_rst_FFX_RST
    );
  rx_input_memio_cs_FFd16_1_1800 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_memio_cs_FFd16_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_memio_cs_FFd16_1_FFX_SET,
      RST => GND,
      O => rx_input_memio_cs_FFd16_1
    );
  rx_input_memio_cs_FFd16_1_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_RESET_1,
      O => rx_input_memio_cs_FFd16_1_FFX_SET
    );
  rx_input_memio_MA_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_11_FFY_RST,
      O => addr1ext(10)
    );
  addr1ext_11_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_11_FFY_RST
    );
  mac_control_rxf_rst_1801 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0047,
      CE => mac_control_rxf_rst_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_rst_FFY_RST,
      O => mac_control_rxf_rst
    );
  mac_control_rxf_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_rst_FFY_RST
    );
  rx_input_memio_MA_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_11_FFX_RST,
      O => addr1ext(11)
    );
  addr1ext_11_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_11_FFX_RST
    );
  rx_input_memio_MA_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_13_FFX_RST,
      O => addr1ext(13)
    );
  addr1ext_13_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_13_FFX_RST
    );
  rx_input_memio_MA_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_13_FFY_RST,
      O => addr1ext(12)
    );
  addr1ext_13_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_13_FFY_RST
    );
  rx_input_memio_MA_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_15_FFX_RST,
      O => addr1ext(15)
    );
  addr1ext_15_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_15_FFX_RST
    );
  rx_input_memio_MA_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lma(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr1ext_15_FFY_RST,
      O => addr1ext(14)
    );
  addr1ext_15_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => addr1ext_15_FFY_RST
    );
  rx_input_memio_MD_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_11_FFY_RST,
      O => d1(10)
    );
  d1_11_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_11_FFY_RST
    );
  rx_output_fifo_BU98 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2299,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1553_FFY_RST,
      O => rx_output_fifo_N1552
    );
  rx_output_fifo_N1553_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1553_FFY_RST
    );
  rx_input_memio_crcl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_0_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_1_FFY_RST,
      O => rx_input_memio_crcl(0)
    );
  rx_input_memio_crcl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_1_FFY_RST
    );
  rx_output_fifo_BU91 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2259,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1553_FFX_RST,
      O => rx_output_fifo_N1553
    );
  rx_output_fifo_N1553_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1553_FFX_RST
    );
  tx_output_crcl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_0_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_1_FFY_RST,
      O => tx_output_crcl(0)
    );
  tx_output_crcl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_1_FFY_RST
    );
  tx_output_crcl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_1_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_1_FFX_RST,
      O => tx_output_crcl(1)
    );
  tx_output_crcl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_1_FFX_RST
    );
  mac_control_sclkdelta_1802 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lsclkdelta,
      CE => mac_control_sclkdelta_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_sclkdelta_FFY_RST,
      O => mac_control_sclkdelta
    );
  mac_control_sclkdelta_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_sclkdelta_FFY_RST
    );
  mac_control_rxphyerr_rst_1803 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0050,
      CE => mac_control_rxphyerr_rst_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_rst_FFY_RST,
      O => mac_control_rxphyerr_rst
    );
  mac_control_rxphyerr_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_rst_FFY_RST
    );
  rx_input_memio_crcl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_1_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_1_FFX_RST,
      O => rx_input_memio_crcl(1)
    );
  rx_input_memio_crcl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_1_FFX_RST
    );
  rx_output_lenr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_7_O,
      CE => rx_output_lenr_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_7_FFY_RST,
      O => rx_output_lenr(7)
    );
  rx_output_lenr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_7_FFY_RST
    );
  rx_output_lenr_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_8_O,
      CE => rx_output_lenr_8_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_8_FFY_RST,
      O => rx_output_lenr(8)
    );
  rx_output_lenr_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_8_FFY_RST
    );
  rx_output_lenr_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0046_9_O,
      CE => rx_output_lenr_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_lenr_9_FFY_RST,
      O => rx_output_lenr(9)
    );
  rx_output_lenr_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_lenr_9_FFY_RST
    );
  tx_input_cs_FFd5_1804 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd5_In1_O,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd6_FFY_RST,
      O => tx_input_cs_FFd5
    );
  tx_input_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd6_FFY_RST
    );
  tx_input_cs_FFd7_1805 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd7_In1_O,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd8_FFY_RST,
      O => tx_input_cs_FFd7
    );
  tx_input_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd8_FFY_RST
    );
  rx_output_fifodin_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(9),
      CE => rx_output_fifodin_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_9_FFX_RST,
      O => rx_output_fifodin(9)
    );
  rx_output_fifodin_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_9_FFX_RST
    );
  rx_output_fifo_full_1806 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_n0051,
      CE => rx_output_fifo_full_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_full_FFY_RST,
      O => rx_output_fifo_full
    );
  rx_output_fifo_full_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifo_full_FFY_RST
    );
  rx_input_GMII_FIFOIN_0 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_GMII_N79913,
      CE => VCC,
      CLK => clkrx,
      SET => GSR,
      RST => GND,
      SSET => rx_input_GMII_rx_erl,
      SRST => GND,
      O => rx_input_fifoin(0)
    );
  rx_input_GMII_FIFOIN_1 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_GMII_N79916,
      CE => VCC,
      CLK => clkrx,
      SET => GSR,
      RST => GND,
      SSET => rx_input_GMII_rx_of,
      SRST => GND,
      O => rx_input_fifoin(1)
    );
  rx_input_GMII_FIFOIN_2 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_GMII_N79919,
      CE => VCC,
      CLK => clkrx,
      SET => GSR,
      RST => GND,
      SSET => rx_input_GMII_rx_of,
      SRST => GND,
      O => rx_input_fifoin(2)
    );
  rx_input_GMII_FIFOIN_3 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_N79922,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_rx_of,
      O => rx_input_fifoin(3)
    );
  rx_input_GMII_FIFOIN_4 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_N79910,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_rx_of,
      O => rx_input_fifoin(4)
    );
  rx_input_GMII_FIFOIN_5 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_N79901,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_rx_of,
      O => rx_input_fifoin(5)
    );
  tx_input_dinint_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(10),
      CE => tx_input_dinint_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_11_FFY_RST,
      O => tx_input_dinint(10)
    );
  tx_input_dinint_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_11_FFY_RST
    );
  rx_input_GMII_FIFOIN_6 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_N79904,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_rx_of,
      O => rx_input_fifoin(6)
    );
  rx_input_GMII_FIFOIN_7 : X_SFF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_N79907,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => GSR,
      SSET => GND,
      SRST => rx_input_GMII_rx_of,
      O => rx_input_fifoin(7)
    );
  rx_input_memio_MD_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_9_FFX_RST,
      O => d1(9)
    );
  d1_9_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => d1_9_FFX_RST
    );
  rx_input_memio_crcl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_21_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_21_FFX_RST,
      O => rx_input_memio_crcl(21)
    );
  rx_input_memio_crcl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_21_FFX_RST
    );
  rx_input_memio_crcl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_20_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_21_FFY_RST,
      O => rx_input_memio_crcl(20)
    );
  rx_input_memio_crcl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_21_FFY_RST
    );
  rx_input_memio_cs_FFd11_1807 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd11_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd12_FFY_RST,
      O => rx_input_memio_cs_FFd11
    );
  rx_input_memio_cs_FFd12_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd12_FFY_RST
    );
  memcontroller_clknum_1_2_1808 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_n0149,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_clknum_1_2_FFX_RST,
      O => memcontroller_clknum_1_2
    );
  memcontroller_clknum_1_2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_1_2_FFX_RST
    );
  rx_input_memio_cs_FFd12_1809 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd12_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd12_FFX_RST,
      O => rx_input_memio_cs_FFd12
    );
  rx_input_memio_cs_FFd12_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd12_FFX_RST
    );
  rx_input_memio_cs_FFd13_1810 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd13_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd14_FFY_RST,
      O => rx_input_memio_cs_FFd13
    );
  rx_input_memio_cs_FFd14_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd14_FFY_RST
    );
  rx_input_memio_cs_FFd14_1811 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd14_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd14_FFX_RST,
      O => rx_input_memio_cs_FFd14
    );
  rx_input_memio_cs_FFd14_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd14_FFX_RST
    );
  rx_input_memio_cs_FFd16_1812 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_memio_cs_FFd16_1_GROM,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_memio_cs_FFd16_1_FFY_SET,
      RST => GND,
      O => rx_input_memio_cs_FFd16
    );
  rx_input_memio_cs_FFd16_1_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_RESET_1,
      O => rx_input_memio_cs_FFd16_1_FFY_SET
    );
  mac_control_rxoferr_rst_1813 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0051,
      CE => mac_control_rxfifowerr_rst_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxfifowerr_rst_FFY_RST,
      O => mac_control_rxoferr_rst
    );
  mac_control_rxfifowerr_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxfifowerr_rst_FFY_RST
    );
  tx_input_dinint_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(11),
      CE => tx_input_dinint_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_11_FFX_RST,
      O => tx_input_dinint(11)
    );
  tx_input_dinint_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_11_FFX_RST
    );
  tx_input_dinint_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(13),
      CE => tx_input_dinint_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_13_FFX_RST,
      O => tx_input_dinint(13)
    );
  tx_input_dinint_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_13_FFX_RST
    );
  tx_input_dinint_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(15),
      CE => tx_input_dinint_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_15_FFX_RST,
      O => tx_input_dinint(15)
    );
  tx_input_dinint_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_15_FFX_RST
    );
  rx_input_memio_RXCRCERR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0060,
      CE => rxfifowerr_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfifowerr_FFY_RST,
      O => rxcrcerr
    );
  rxfifowerr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfifowerr_FFY_RST
    );
  rx_input_memio_RXFIFOWERR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0061,
      CE => rxfifowerr_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxfifowerr_FFX_RST,
      O => rxfifowerr
    );
  rxfifowerr_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxfifowerr_FFX_RST
    );
  rx_output_cs_FFd17_1814 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd17_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd17_FFY_RST,
      O => rx_output_cs_FFd17
    );
  rx_output_cs_FFd17_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd17_FFY_RST
    );
  rx_input_memio_MD_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(25),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_25_FFX_RST,
      O => d1(25)
    );
  d1_25_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_25_FFX_RST
    );
  rx_input_memio_MD_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(16),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_17_FFY_RST,
      O => d1(16)
    );
  d1_17_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_17_FFY_RST
    );
  rx_input_memio_MD_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(17),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_17_FFX_RST,
      O => d1(17)
    );
  d1_17_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_17_FFX_RST
    );
  rx_input_memio_MD_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(26),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_27_FFY_RST,
      O => d1(26)
    );
  d1_27_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_27_FFY_RST
    );
  rx_input_memio_MD_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(27),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_27_FFX_RST,
      O => d1(27)
    );
  d1_27_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_27_FFX_RST
    );
  rx_input_memio_MD_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(18),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_19_FFY_RST,
      O => d1(18)
    );
  d1_19_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_19_FFY_RST
    );
  rx_input_memio_MD_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(19),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_19_FFX_RST,
      O => d1(19)
    );
  d1_19_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_19_FFX_RST
    );
  rx_input_memio_MD_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(28),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_29_FFY_RST,
      O => d1(28)
    );
  d1_29_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_29_FFY_RST
    );
  rx_output_fifodin_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(10),
      CE => rx_output_fifodin_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_11_FFY_RST,
      O => rx_output_fifodin(10)
    );
  rx_output_fifodin_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_11_FFY_RST
    );
  rx_input_memio_MD_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_lmd(29),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d1_29_FFX_RST,
      O => d1(29)
    );
  d1_29_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => d1_29_FFX_RST
    );
  tx_output_cs_FFd16_1815 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd16_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd16_FFX_RST,
      O => tx_output_cs_FFd16
    );
  tx_output_cs_FFd16_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd16_FFX_RST
    );
  rx_output_fifodin_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(0),
      CE => rx_output_fifodin_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_1_FFY_RST,
      O => rx_output_fifodin(0)
    );
  rx_output_fifodin_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_1_FFY_RST
    );
  rx_output_fifodin_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(1),
      CE => rx_output_fifodin_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_1_FFX_RST,
      O => rx_output_fifodin(1)
    );
  rx_output_fifodin_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_1_FFX_RST
    );
  rx_output_fifodin_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(2),
      CE => rx_output_fifodin_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_3_FFY_RST,
      O => rx_output_fifodin(2)
    );
  rx_output_fifodin_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_3_FFY_RST
    );
  rx_output_fifodin_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(3),
      CE => rx_output_fifodin_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_3_FFX_RST,
      O => rx_output_fifodin(3)
    );
  rx_output_fifodin_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_3_FFX_RST
    );
  rx_output_fifodin_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(4),
      CE => rx_output_fifodin_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_5_FFY_RST,
      O => rx_output_fifodin(4)
    );
  rx_output_fifodin_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_5_FFY_RST
    );
  rx_output_fifodin_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(5),
      CE => rx_output_fifodin_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_5_FFX_RST,
      O => rx_output_fifodin(5)
    );
  rx_output_fifodin_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_5_FFX_RST
    );
  rx_output_fifodin_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(6),
      CE => rx_output_fifodin_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_7_FFY_RST,
      O => rx_output_fifodin(6)
    );
  rx_output_fifodin_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_7_FFY_RST
    );
  rx_output_fifodin_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(7),
      CE => rx_output_fifodin_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_7_FFX_RST,
      O => rx_output_fifodin(7)
    );
  rx_output_fifodin_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_7_FFX_RST
    );
  rx_output_fifodin_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(8),
      CE => rx_output_fifodin_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_9_FFY_RST,
      O => rx_output_fifodin(8)
    );
  rx_output_fifodin_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_9_FFY_RST
    );
  rx_input_memio_cs_FFd2_1816 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd4,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd2_FFY_RST,
      O => rx_input_memio_cs_FFd2
    );
  rx_input_memio_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd2_FFY_RST
    );
  mac_control_txfifowerr_cntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(6),
      CE => mac_control_txfifowerr_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_7_FFY_RST,
      O => mac_control_txfifowerr_cntl(6)
    );
  mac_control_txfifowerr_cntl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_7_FFY_RST
    );
  mac_control_txfifowerr_cntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(7),
      CE => mac_control_txfifowerr_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_7_FFX_RST,
      O => mac_control_txfifowerr_cntl(7)
    );
  mac_control_txfifowerr_cntl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_7_FFX_RST
    );
  mac_control_txfifowerr_cntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(8),
      CE => mac_control_txfifowerr_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_9_FFY_RST,
      O => mac_control_txfifowerr_cntl(8)
    );
  mac_control_txfifowerr_cntl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_9_FFY_RST
    );
  mac_control_txfifowerr_cntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(9),
      CE => mac_control_txfifowerr_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_9_FFX_RST,
      O => mac_control_txfifowerr_cntl(9)
    );
  mac_control_txfifowerr_cntl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_9_FFX_RST
    );
  rx_input_memio_cs_FFd5_1817 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd6,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd6_FFY_RST,
      O => rx_input_memio_cs_FFd5
    );
  rx_input_memio_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd6_FFY_RST
    );
  rx_input_memio_cs_FFd6_1818 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd7,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd6_FFX_RST,
      O => rx_input_memio_cs_FFd6
    );
  rx_input_memio_cs_FFd6_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd6_FFX_RST
    );
  tx_output_crcl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_23_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_23_FFY_RST,
      O => tx_output_crcl(23)
    );
  tx_output_crcl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_23_FFY_RST
    );
  rx_input_memio_bcnt_88_1819 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bcnt_inst_sum_237,
      CE => rx_input_memio_n0102,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bcnt_88_FFY_RST,
      O => rx_input_memio_bcnt_88
    );
  rx_input_memio_bcnt_88_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_bcnt_88_FFY_RST
    );
  rx_input_memio_crcl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_10_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_10_FFY_RST,
      O => rx_input_memio_crcl(10)
    );
  rx_input_memio_crcl_10_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_10_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(2),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_3_FFY_RST,
      O => mac_control_phydo(2)
    );
  mac_control_phydo_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_3_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(0),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_1_FFY_RST,
      O => mac_control_phydo(0)
    );
  mac_control_phydo_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_1_FFY_RST
    );
  rx_output_fifodin_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(11),
      CE => rx_output_fifodin_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_11_FFX_RST,
      O => rx_output_fifodin(11)
    );
  rx_output_fifodin_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_11_FFX_RST
    );
  rx_output_fifodin_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(12),
      CE => rx_output_fifodin_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_13_FFY_RST,
      O => rx_output_fifodin(12)
    );
  rx_output_fifodin_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_13_FFY_RST
    );
  rx_output_fifodin_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(13),
      CE => rx_output_fifodin_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_13_FFX_RST,
      O => rx_output_fifodin(13)
    );
  rx_output_fifodin_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_13_FFX_RST
    );
  rx_output_fifodin_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(14),
      CE => rx_output_fifodin_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_15_FFY_RST,
      O => rx_output_fifodin(14)
    );
  rx_output_fifodin_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_15_FFY_RST
    );
  rx_output_fifodin_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_lma(15),
      CE => rx_output_fifodin_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifodin_15_FFX_RST,
      O => rx_output_fifodin(15)
    );
  rx_output_fifodin_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_fifodin_15_FFX_RST
    );
  tx_input_enableintl_1820 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_enableintl_GSHIFT,
      CE => tx_input_enableintl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_enableintl_FFY_RST,
      O => tx_input_enableintl
    );
  tx_input_enableintl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_enableintl_FFY_RST
    );
  mac_control_PHY_status_cs_FFd1_1821 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd1_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd2_FFY_RST,
      O => mac_control_PHY_status_cs_FFd1
    );
  mac_control_PHY_status_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd2_FFY_RST
    );
  mac_control_PHY_status_cs_FFd3_1822 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd4_FFY_RST,
      O => mac_control_PHY_status_cs_FFd3
    );
  mac_control_PHY_status_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd4_FFY_RST
    );
  mac_control_PHY_status_cs_FFd2_1823 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd2_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd2_FFX_RST,
      O => mac_control_PHY_status_cs_FFd2
    );
  mac_control_PHY_status_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd2_FFX_RST
    );
  rx_output_cs_FFd19_1824 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_cs_FFd19_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_cs_FFd4_FFY_SET,
      RST => GND,
      O => rx_output_cs_FFd19
    );
  rx_output_cs_FFd4_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => rx_output_cs_FFd4_FFY_SET
    );
  rx_output_cs_FFd4_1825 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd4_FFX_RST,
      O => rx_output_cs_FFd4
    );
  rx_output_cs_FFd4_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd4_FFX_RST
    );
  rx_input_memio_RXPHYERR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0057,
      CE => rxoferr_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxoferr_FFY_RST,
      O => rxphyerr
    );
  rxoferr_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxoferr_FFY_RST
    );
  rx_input_memio_RXOFERR : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0058,
      CE => rxoferr_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxoferr_FFX_RST,
      O => rxoferr
    );
  rxoferr_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxoferr_FFX_RST
    );
  tx_input_cs_FFd11_1826 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd11_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd11_FFY_RST,
      O => tx_input_cs_FFd11
    );
  tx_input_cs_FFd11_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd11_FFY_RST
    );
  mac_control_txf_cross_1827 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cross_GROM,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_txf_cross_FFY_RST,
      O => mac_control_txf_cross
    );
  mac_control_txf_cross_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cross_FFY_RST
    );
  tx_input_CNT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(10),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_11_FFY_RST,
      O => tx_input_CNT(10)
    );
  tx_input_CNT_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_11_FFY_RST
    );
  tx_input_CNT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(11),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_11_FFX_RST,
      O => tx_input_CNT(11)
    );
  tx_input_CNT_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_11_FFX_RST
    );
  tx_input_CNT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(13),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_13_FFX_RST,
      O => tx_input_CNT(13)
    );
  tx_input_CNT_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_13_FFX_RST
    );
  tx_input_CNT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(12),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_13_FFY_RST,
      O => tx_input_CNT(12)
    );
  tx_input_CNT_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_13_FFY_RST
    );
  tx_input_CNT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(14),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_15_FFY_RST,
      O => tx_input_CNT(14)
    );
  tx_input_CNT_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_15_FFY_RST
    );
  mac_control_PHY_status_cs_FFd4_1828 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd4_FFX_RST,
      O => mac_control_PHY_status_cs_FFd4
    );
  mac_control_PHY_status_cs_FFd4_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd4_FFX_RST
    );
  mac_control_PHY_status_cs_FFd5_1829 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd5_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd6_FFY_RST,
      O => mac_control_PHY_status_cs_FFd5
    );
  mac_control_PHY_status_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd6_FFY_RST
    );
  mac_control_PHY_status_cs_FFd6_1830 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd6_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd6_FFX_RST,
      O => mac_control_PHY_status_cs_FFd6
    );
  mac_control_PHY_status_cs_FFd6_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd6_FFX_RST
    );
  mac_control_PHY_status_cs_FFd7_1831 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd7_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_cs_FFd8_FFY_RST,
      O => mac_control_PHY_status_cs_FFd7
    );
  mac_control_PHY_status_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => mac_control_PHY_status_cs_FFd8_FFY_RST
    );
  mac_control_PHY_status_cs_FFd8_1832 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => mac_control_PHY_status_cs_FFd8_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => mac_control_PHY_status_cs_FFd8_FFX_SET,
      RST => GND,
      O => mac_control_PHY_status_cs_FFd8
    );
  mac_control_PHY_status_cs_FFd8_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => mac_control_PHY_status_cs_FFd8_FFX_SET
    );
  rx_input_memio_crcen_1833 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0049,
      CE => rx_input_memio_crcen_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcen_FFY_RST,
      O => rx_input_memio_crcen
    );
  rx_input_memio_crcen_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcen_FFY_RST
    );
  tx_input_den_1834 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_lden,
      CE => tx_input_den_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_den_FFY_RST,
      O => tx_input_den
    );
  tx_input_den_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_den_FFY_RST
    );
  tx_input_CNT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(0),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_1_FFY_RST,
      O => tx_input_CNT(0)
    );
  tx_input_CNT_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_1_FFY_RST
    );
  tx_input_CNT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(2),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_3_FFY_RST,
      O => tx_input_CNT(2)
    );
  tx_input_CNT_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_3_FFY_RST
    );
  rx_input_memio_doutl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(7),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_7_FFX_RST,
      O => rx_input_memio_doutl(7)
    );
  rx_input_memio_doutl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_7_FFX_RST
    );
  rx_input_memio_doutl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(8),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_9_FFY_RST,
      O => rx_input_memio_doutl(8)
    );
  rx_input_memio_doutl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_9_FFY_RST
    );
  rx_input_memio_doutl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(9),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_9_FFX_RST,
      O => rx_input_memio_doutl(9)
    );
  rx_input_memio_doutl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_9_FFX_RST
    );
  rx_input_memio_wbpl_1835 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd2,
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_wbpl_FFY_RST,
      O => rx_input_memio_wbpl
    );
  rx_input_memio_wbpl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_wbpl_FFY_RST
    );
  rx_input_memio_crcl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_19_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_19_FFY_RST,
      O => rx_input_memio_crcl(19)
    );
  rx_input_memio_crcl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_19_FFY_RST
    );
  rx_input_memio_crcl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_13_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_13_FFY_RST,
      O => rx_input_memio_crcl(13)
    );
  rx_input_memio_crcl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_13_FFY_RST
    );
  tx_output_crcl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_27_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_27_FFY_RST,
      O => tx_output_crcl(27)
    );
  tx_output_crcl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_27_FFY_RST
    );
  rx_output_cs_FFd6_1836 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd6_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd6_FFY_RST,
      O => rx_output_cs_FFd6
    );
  rx_output_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd6_FFY_RST
    );
  rx_input_memio_crcl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_30_1_O,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_30_FFY_RST,
      O => rx_input_memio_crcl(30)
    );
  rx_input_memio_crcl_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_30_FFY_RST
    );
  tx_input_dinint_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(5),
      CE => tx_input_dinint_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_5_FFX_RST,
      O => tx_input_dinint(5)
    );
  tx_input_dinint_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_5_FFX_RST
    );
  tx_input_dinint_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(6),
      CE => tx_input_dinint_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_7_FFY_RST,
      O => tx_input_dinint(6)
    );
  tx_input_dinint_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_7_FFY_RST
    );
  tx_input_dinint_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(7),
      CE => tx_input_dinint_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_7_FFX_RST,
      O => tx_input_dinint(7)
    );
  tx_input_dinint_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_7_FFX_RST
    );
  tx_input_dinint_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(8),
      CE => tx_input_dinint_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_9_FFY_RST,
      O => tx_input_dinint(8)
    );
  tx_input_dinint_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_9_FFY_RST
    );
  tx_input_dinint_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(9),
      CE => tx_input_dinint_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_9_FFX_RST,
      O => tx_input_dinint(9)
    );
  tx_input_dinint_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_9_FFX_RST
    );
  rx_input_fifo_control_cs_FFd1_1837 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_cs_FFd1_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_cs_FFd2_FFY_RST,
      O => rx_input_fifo_control_cs_FFd1
    );
  rx_input_fifo_control_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_cs_FFd2_FFY_RST
    );
  rx_input_fifo_control_cs_FFd2_1838 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_cs_FFd2_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_cs_FFd2_FFX_RST,
      O => rx_input_fifo_control_cs_FFd2
    );
  rx_input_fifo_control_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_cs_FFd2_FFX_RST
    );
  rx_output_cs_FFd1_1839 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd1_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd2_FFY_RST,
      O => rx_output_cs_FFd1
    );
  rx_output_cs_FFd2_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd2_FFY_RST
    );
  rx_output_cs_FFd7_1840 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd7_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd8_FFY_RST,
      O => rx_output_cs_FFd7
    );
  rx_output_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd8_FFY_RST
    );
  rx_output_cs_FFd2_1841 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd2_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd2_FFX_RST,
      O => rx_output_cs_FFd2
    );
  rx_output_cs_FFd2_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd2_FFX_RST
    );
  tx_input_CNT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_n0032(15),
      CE => tx_input_N35872,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_CNT_15_FFX_RST,
      O => tx_input_CNT(15)
    );
  tx_input_CNT_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_CNT_15_FFX_RST
    );
  tx_output_cs_FFd5_1_1842 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd5_GROM,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd5_FFY_RST,
      O => tx_output_cs_FFd5_1
    );
  tx_output_cs_FFd5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd5_FFY_RST
    );
  tx_input_dinint_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(0),
      CE => tx_input_dinint_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_1_FFY_RST,
      O => tx_input_dinint(0)
    );
  tx_input_dinint_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_1_FFY_RST
    );
  tx_output_cs_FFd6_1_1843 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd6_GROM,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd6_FFY_RST,
      O => tx_output_cs_FFd6_1
    );
  tx_output_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd6_FFY_RST
    );
  tx_output_cs_FFd5_1844 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd5_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd5_FFX_RST,
      O => tx_output_cs_FFd5
    );
  tx_output_cs_FFd5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd5_FFX_RST
    );
  tx_output_cs_FFd6_1845 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd6_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd6_FFX_RST,
      O => tx_output_cs_FFd6
    );
  tx_output_cs_FFd6_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd6_FFX_RST
    );
  tx_input_dinint_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(1),
      CE => tx_input_dinint_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_1_FFX_RST,
      O => tx_input_dinint(1)
    );
  tx_input_dinint_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_1_FFX_RST
    );
  tx_input_dinint_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(2),
      CE => tx_input_dinint_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_3_FFY_RST,
      O => tx_input_dinint(2)
    );
  tx_input_dinint_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_3_FFY_RST
    );
  tx_input_dinint_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(3),
      CE => tx_input_dinint_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_3_FFX_RST,
      O => tx_input_dinint(3)
    );
  tx_input_dinint_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_3_FFX_RST
    );
  tx_input_dinint_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_ldinint(4),
      CE => tx_input_dinint_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dinint_5_FFY_RST,
      O => tx_input_dinint(4)
    );
  tx_input_dinint_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dinint_5_FFY_RST
    );
  rx_output_cs_FFd8_1846 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd8_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd8_FFX_RST,
      O => rx_output_cs_FFd8
    );
  rx_output_cs_FFd8_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd8_FFX_RST
    );
  rx_input_GMII_INCE : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_lince,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_ince_FFY_RST,
      O => rx_input_ince
    );
  rx_input_ince_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_ince_FFY_RST
    );
  tx_input_cs_FFd2_1847 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd2_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd4_FFY_RST,
      O => tx_input_cs_FFd2
    );
  tx_input_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd4_FFY_RST
    );
  tx_input_cs_FFd4_1848 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd8,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd4_FFX_RST,
      O => tx_input_cs_FFd4
    );
  tx_input_cs_FFd4_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd4_FFX_RST
    );
  tx_input_cs_FFd3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfifowerr_FFY_RST,
      O => txfifowerr
    );
  txfifowerr_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => txfifowerr_FFY_RST
    );
  tx_input_cs_FFd9_1849 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd9_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd10_FFY_RST,
      O => tx_input_cs_FFd9
    );
  tx_input_cs_FFd10_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd10_FFY_RST
    );
  tx_input_cs_FFd10_1850 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_cs_FFd10_In_O,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_cs_FFd10_FFX_RST,
      O => tx_input_cs_FFd10
    );
  tx_input_cs_FFd10_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => tx_input_cs_FFd10_FFX_RST
    );
  rx_input_memio_Mshreg_lbpout4_10_59_1851 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_10_net14,
      CE => rx_input_memio_Mshreg_lbpout4_10_59_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_10_59_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_10_59
    );
  rx_input_memio_Mshreg_lbpout4_10_59_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_10_59_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_11_58_1852 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_11_net12,
      CE => rx_input_memio_Mshreg_lbpout4_11_58_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_11_58_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_11_58
    );
  rx_input_memio_Mshreg_lbpout4_11_58_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_11_58_FFY_RST
    );
  rx_output_fifo_BU464 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N1589_FROM,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1589_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1589
    );
  rx_output_fifo_N1589_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1589_FFX_SET
    );
  rx_output_fifo_BU458 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3969,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1593_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1592
    );
  rx_output_fifo_N1593_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1593_FFY_SET
    );
  rx_output_fifo_BU456 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3968,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1593_FFX_SET,
      RST => GND,
      O => rx_output_fifo_N1593
    );
  rx_output_fifo_N1593_FFX_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1593_FFX_SET
    );
  tx_output_cs_FFd8_1853 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd8_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd8_FFX_RST,
      O => tx_output_cs_FFd8
    );
  tx_output_cs_FFd8_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd8_FFX_RST
    );
  tx_output_cs_FFd7_1854 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd7_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_cs_FFd8_FFY_RST,
      O => tx_output_cs_FFd7
    );
  tx_output_cs_FFd8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => tx_output_cs_FFd8_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_0_69_1855 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_0_net34,
      CE => rx_input_memio_Mshreg_lbpout4_0_69_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_0_69_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_0_69
    );
  rx_input_memio_Mshreg_lbpout4_0_69_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_0_69_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_1_68_1856 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_1_net32,
      CE => rx_input_memio_Mshreg_lbpout4_1_68_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_1_68_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_1_68
    );
  rx_input_memio_Mshreg_lbpout4_1_68_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_1_68_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_2_67_1857 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_2_net30,
      CE => rx_input_memio_Mshreg_lbpout4_2_67_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_2_67_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_2_67
    );
  rx_input_memio_Mshreg_lbpout4_2_67_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_2_67_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_3_66_1858 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_3_net28,
      CE => rx_input_memio_Mshreg_lbpout4_3_66_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_3_66_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_3_66
    );
  rx_input_memio_Mshreg_lbpout4_3_66_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_3_66_FFY_RST
    );
  rx_fifocheck_bpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_9_FFX_RST,
      O => rx_fifocheck_bpl(9)
    );
  rx_fifocheck_bpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_9_FFX_RST
    );
  tx_output_crcl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_13_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_13_FFY_RST,
      O => tx_output_crcl(13)
    );
  tx_output_crcl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_13_FFY_RST
    );
  rx_input_memio_crcl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_6_1_O,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_6_FFY_RST,
      O => rx_input_memio_crcl(6)
    );
  rx_input_memio_crcl_6_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_6_FFY_RST
    );
  rx_fifocheck_bpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_11_FFX_RST,
      O => rx_fifocheck_bpl(11)
    );
  rx_fifocheck_bpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_11_FFX_RST
    );
  rx_fifocheck_bpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_11_FFY_RST,
      O => rx_fifocheck_bpl(10)
    );
  rx_fifocheck_bpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_11_FFY_RST
    );
  rx_fifocheck_bpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_13_FFY_RST,
      O => rx_fifocheck_bpl(12)
    );
  rx_fifocheck_bpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_13_FFY_RST
    );
  rx_fifocheck_bpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_13_FFX_RST,
      O => rx_fifocheck_bpl(13)
    );
  rx_fifocheck_bpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_13_FFX_RST
    );
  rx_fifocheck_bpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_15_FFY_RST,
      O => rx_fifocheck_bpl(14)
    );
  rx_fifocheck_bpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_15_FFY_RST
    );
  rx_fifocheck_bpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_15_FFX_RST,
      O => rx_fifocheck_bpl(15)
    );
  rx_fifocheck_bpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_15_FFX_RST
    );
  tx_output_crcsell_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd3,
      CE => tx_output_crcsell_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcsell_3_FFY_RST,
      O => tx_output_crcsell(2)
    );
  tx_output_crcsell_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcsell_3_FFY_RST
    );
  tx_output_crcsell_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd7,
      CE => tx_output_crcsell_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcsell_3_FFX_RST,
      O => tx_output_crcsell(3)
    );
  tx_output_crcsell_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcsell_3_FFX_RST
    );
  memcontroller_dnl2_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(0),
      CE => memcontroller_dnl2_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_1_FFY_RST,
      O => memcontroller_dnl2(0)
    );
  memcontroller_dnl2_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_1_FFY_RST
    );
  rx_output_fifo_BU119 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2419,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1549_FFX_RST,
      O => rx_output_fifo_N1549
    );
  rx_output_fifo_N1549_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1549_FFX_RST
    );
  rx_output_fifo_BU266 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3267,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1615_FFX_RST,
      O => rx_output_fifo_N1615
    );
  rx_output_fifo_N1615_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1615_FFX_RST
    );
  rx_output_fifo_BU259 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3227,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1617_FFY_RST,
      O => rx_output_fifo_N1616
    );
  rx_output_fifo_N1617_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1617_FFY_RST
    );
  rx_output_fifo_BU252 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3187,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1617_FFX_RST,
      O => rx_output_fifo_N1617
    );
  rx_output_fifo_N1617_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1617_FFX_RST
    );
  rx_output_fifo_BU287 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3387,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1613_FFY_RST,
      O => rx_output_fifo_N1612
    );
  rx_output_fifo_N1613_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1613_FFY_RST
    );
  rx_output_fifo_BU280 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3347,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1613_FFX_RST,
      O => rx_output_fifo_N1613
    );
  rx_output_fifo_N1613_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1613_FFX_RST
    );
  rx_output_fifo_BU462 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3971,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1589_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1590
    );
  rx_output_fifo_N1589_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1589_FFY_SET
    );
  rx_output_fifo_BU466 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_output_fifo_N3973,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_output_fifo_N1588_FFY_SET,
      RST => GND,
      O => rx_output_fifo_N1588
    );
  rx_output_fifo_N1588_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_output_fifo_reset,
      O => rx_output_fifo_N1588_FFY_SET
    );
  rx_input_memio_Mshreg_lbpout4_12_57_1859 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_12_net10,
      CE => rx_input_memio_Mshreg_lbpout4_12_57_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_12_57_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_12_57
    );
  rx_input_memio_Mshreg_lbpout4_12_57_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_12_57_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_13_56_1860 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_13_net8,
      CE => rx_input_memio_Mshreg_lbpout4_13_56_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_13_56_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_13_56
    );
  rx_input_memio_Mshreg_lbpout4_13_56_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_13_56_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_14_55_1861 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_14_net6,
      CE => rx_input_memio_Mshreg_lbpout4_14_55_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_14_55_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_14_55
    );
  rx_input_memio_Mshreg_lbpout4_14_55_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_14_55_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_15_54_1862 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_15_net4,
      CE => rx_input_memio_Mshreg_lbpout4_15_54_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_15_54_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_15_54
    );
  rx_input_memio_Mshreg_lbpout4_15_54_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_15_54_FFY_RST
    );
  mac_control_Mshreg_sinlll_102_1863 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_Mshreg_sinlll_net185,
      CE => mac_control_Mshreg_sinlll_102_CEMUXNOT,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_Mshreg_sinlll_102_FFY_RST,
      O => mac_control_Mshreg_sinlll_102
    );
  mac_control_Mshreg_sinlll_102_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_Mshreg_sinlll_102_FFY_RST
    );
  rx_output_fifo_BU112 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2379,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1551_FFY_RST,
      O => rx_output_fifo_N1550
    );
  rx_output_fifo_N1551_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1551_FFY_RST
    );
  rx_output_fifo_BU105 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2339,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1551_FFX_RST,
      O => rx_output_fifo_N1551
    );
  rx_output_fifo_N1551_FFX_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1551_FFX_RST
    );
  rx_output_fifo_BU273 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N3307,
      CE => rx_output_fifo_N1517,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_fifo_N1615_FFY_RST,
      O => rx_output_fifo_N1614
    );
  rx_output_fifo_N1615_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1615_FFY_RST
    );
  rx_output_fifo_BU126 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_fifo_N2459,
      CE => rx_output_fifo_N1515,
      CLK => clkio,
      SET => GND,
      RST => rx_output_fifo_N1549_FFY_RST,
      O => rx_output_fifo_N1548
    );
  rx_output_fifo_N1549_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_output_fifo_reset,
      I1 => GSR,
      O => rx_output_fifo_N1549_FFY_RST
    );
  memcontroller_dnl2_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(1),
      CE => memcontroller_dnl2_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_1_FFX_RST,
      O => memcontroller_dnl2(1)
    );
  memcontroller_dnl2_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_1_FFX_RST
    );
  memcontroller_dnl2_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(2),
      CE => memcontroller_dnl2_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_3_FFY_RST,
      O => memcontroller_dnl2(2)
    );
  memcontroller_dnl2_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_3_FFY_RST
    );
  memcontroller_dnl2_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(3),
      CE => memcontroller_dnl2_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_3_FFX_RST,
      O => memcontroller_dnl2(3)
    );
  memcontroller_dnl2_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_3_FFX_RST
    );
  tx_output_crcl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_30_1_O,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_30_FFY_RST,
      O => tx_output_crcl(30)
    );
  tx_output_crcl_30_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_30_FFY_RST
    );
  memcontroller_dnl2_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(5),
      CE => memcontroller_dnl2_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_5_FFX_RST,
      O => memcontroller_dnl2(5)
    );
  memcontroller_dnl2_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_5_FFX_RST
    );
  memcontroller_dnl2_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(4),
      CE => memcontroller_dnl2_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_5_FFY_RST,
      O => memcontroller_dnl2(4)
    );
  memcontroller_dnl2_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_5_FFY_RST
    );
  memcontroller_dnl2_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(6),
      CE => memcontroller_dnl2_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_7_FFY_RST,
      O => memcontroller_dnl2(6)
    );
  memcontroller_dnl2_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_7_FFY_RST
    );
  memcontroller_dnl2_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(7),
      CE => memcontroller_dnl2_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_7_FFX_RST,
      O => memcontroller_dnl2(7)
    );
  memcontroller_dnl2_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_7_FFX_RST
    );
  memcontroller_dnl2_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(8),
      CE => memcontroller_dnl2_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_9_FFY_RST,
      O => memcontroller_dnl2(8)
    );
  memcontroller_dnl2_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_9_FFY_RST
    );
  memcontroller_dnl2_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(9),
      CE => memcontroller_dnl2_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_9_FFX_RST,
      O => memcontroller_dnl2(9)
    );
  memcontroller_dnl2_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_9_FFX_RST
    );
  tx_output_crcl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_14_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_14_FFY_RST,
      O => tx_output_crcl(14)
    );
  tx_output_crcl_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_14_FFY_RST
    );
  mac_control_sclkdeltal_1864 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_sclkdelta,
      CE => mac_control_sclkdeltal_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_sclkdeltal_FFY_RST,
      O => mac_control_sclkdeltal
    );
  mac_control_sclkdeltal_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_sclkdeltal_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_4_65_1865 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_4_net26,
      CE => rx_input_memio_Mshreg_lbpout4_4_65_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_4_65_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_4_65
    );
  rx_input_memio_Mshreg_lbpout4_4_65_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_4_65_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_5_64_1866 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_5_net24,
      CE => rx_input_memio_Mshreg_lbpout4_5_64_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_5_64_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_5_64
    );
  rx_input_memio_Mshreg_lbpout4_5_64_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_5_64_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_6_63_1867 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_6_net22,
      CE => rx_input_memio_Mshreg_lbpout4_6_63_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_6_63_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_6_63
    );
  rx_input_memio_Mshreg_lbpout4_6_63_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_6_63_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_7_62_1868 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_7_net20,
      CE => rx_input_memio_Mshreg_lbpout4_7_62_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_7_62_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_7_62
    );
  rx_input_memio_Mshreg_lbpout4_7_62_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_7_62_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_8_61_1869 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_8_net18,
      CE => rx_input_memio_Mshreg_lbpout4_8_61_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_8_61_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_8_61
    );
  rx_input_memio_Mshreg_lbpout4_8_61_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_8_61_FFY_RST
    );
  rx_input_memio_Mshreg_lbpout4_9_60_1870 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_9_net16,
      CE => rx_input_memio_Mshreg_lbpout4_9_60_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_Mshreg_lbpout4_9_60_FFY_RST,
      O => rx_input_memio_Mshreg_lbpout4_9_60
    );
  rx_input_memio_Mshreg_lbpout4_9_60_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_Mshreg_lbpout4_9_60_FFY_RST
    );
  tx_output_crcl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_20_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_21_FFY_RST,
      O => tx_output_crcl(20)
    );
  tx_output_crcl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_21_FFY_RST
    );
  tx_input_newfint_1871 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_lnewfint,
      CE => tx_input_newfint_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_newfint_FFY_RST,
      O => tx_input_newfint
    );
  tx_input_newfint_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_newfint_FFY_RST
    );
  tx_output_crcl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_21_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_21_FFX_RST,
      O => tx_output_crcl(21)
    );
  tx_output_crcl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_21_FFX_RST
    );
  tx_output_crcl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_22_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_22_FFY_RST,
      O => tx_output_crcl(22)
    );
  tx_output_crcl_22_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_22_FFY_RST
    );
  tx_output_crcl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_31_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_31_FFY_RST,
      O => tx_output_crcl(31)
    );
  tx_output_crcl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_31_FFY_RST
    );
  rx_fifocheck_bpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_1_FFY_RST,
      O => rx_fifocheck_bpl(0)
    );
  rx_fifocheck_bpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_1_FFY_RST
    );
  rx_fifocheck_bpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_1_FFX_RST,
      O => rx_fifocheck_bpl(1)
    );
  rx_fifocheck_bpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_1_FFX_RST
    );
  rx_fifocheck_bpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_3_FFY_RST,
      O => rx_fifocheck_bpl(2)
    );
  rx_fifocheck_bpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_3_FFY_RST
    );
  rx_fifocheck_bpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_3_FFX_RST,
      O => rx_fifocheck_bpl(3)
    );
  rx_fifocheck_bpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_3_FFX_RST
    );
  rx_fifocheck_bpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_5_FFY_RST,
      O => rx_fifocheck_bpl(4)
    );
  rx_fifocheck_bpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_5_FFY_RST
    );
  rx_fifocheck_bpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_5_FFX_RST,
      O => rx_fifocheck_bpl(5)
    );
  rx_fifocheck_bpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_5_FFX_RST
    );
  rx_fifocheck_bpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_7_FFY_RST,
      O => rx_fifocheck_bpl(6)
    );
  rx_fifocheck_bpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_7_FFY_RST
    );
  rx_fifocheck_bpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_7_FFX_RST,
      O => rx_fifocheck_bpl(7)
    );
  rx_fifocheck_bpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_7_FFX_RST
    );
  rx_fifocheck_bpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbp(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_bpl_9_FFY_RST,
      O => rx_fifocheck_bpl(8)
    );
  rx_fifocheck_bpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_bpl_9_FFY_RST
    );
  tx_output_crcl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_19_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_19_FFY_RST,
      O => tx_output_crcl(19)
    );
  tx_output_crcl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_19_FFY_RST
    );
  rx_input_memio_dout_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_23_FFX_RST,
      O => rx_input_memio_dout(23)
    );
  rx_input_memio_dout_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_23_FFX_RST
    );
  rx_input_memio_dout_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_15_FFX_RST,
      O => rx_input_memio_dout(15)
    );
  rx_input_memio_dout_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_15_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(13),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_14_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(14)
    );
  mac_control_PHY_status_MII_Interface_dreg_14_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_14_FFX_RST
    );
  rx_input_memio_dout_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_25_FFY_RST,
      O => rx_input_memio_dout(24)
    );
  rx_input_memio_dout_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_25_FFY_RST
    );
  rx_input_memio_dout_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_25_FFX_RST,
      O => rx_input_memio_dout(25)
    );
  rx_input_memio_dout_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_25_FFX_RST
    );
  rx_input_memio_dout_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_17_FFX_RST,
      O => rx_input_memio_dout(17)
    );
  rx_input_memio_dout_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_17_FFX_RST
    );
  rx_input_memio_dout_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_27_FFY_RST,
      O => rx_input_memio_dout(26)
    );
  rx_input_memio_dout_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_27_FFY_RST
    );
  rx_input_memio_dout_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_27_FFX_RST,
      O => rx_input_memio_dout(27)
    );
  rx_input_memio_dout_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_27_FFX_RST
    );
  rx_input_memio_dout_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_19_FFX_RST,
      O => rx_input_memio_dout(19)
    );
  rx_input_memio_dout_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_19_FFX_RST
    );
  rx_input_memio_dout_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_29_FFX_RST,
      O => rx_input_memio_dout(29)
    );
  rx_input_memio_dout_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_29_FFX_RST
    );
  rx_input_memio_crcl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_7_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_7_FFY_RST,
      O => rx_input_memio_crcl(7)
    );
  rx_input_memio_crcl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_7_FFY_RST
    );
  rx_input_memio_addrchk_datal_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_1_FFX_RST,
      O => rx_input_memio_addrchk_datal(1)
    );
  rx_input_memio_addrchk_datal_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_1_FFX_RST
    );
  rx_input_memio_addrchk_datal_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_1_FFY_RST,
      O => rx_input_memio_addrchk_datal(0)
    );
  rx_input_memio_addrchk_datal_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_1_FFY_RST
    );
  rx_input_memio_addrchk_datal_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_3_FFY_RST,
      O => rx_input_memio_addrchk_datal(2)
    );
  rx_input_memio_addrchk_datal_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_3_FFY_RST
    );
  rx_input_memio_addrchk_datal_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_3_FFX_RST,
      O => rx_input_memio_addrchk_datal(3)
    );
  rx_input_memio_addrchk_datal_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_3_FFX_RST
    );
  rx_input_memio_addrchk_datal_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_5_FFY_RST,
      O => rx_input_memio_addrchk_datal(4)
    );
  rx_input_memio_addrchk_datal_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_5_FFY_RST
    );
  rx_input_memio_addrchk_datal_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_5_FFX_RST,
      O => rx_input_memio_addrchk_datal(5)
    );
  rx_input_memio_addrchk_datal_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_5_FFX_RST
    );
  rx_input_memio_addrchk_datal_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_7_FFY_RST,
      O => rx_input_memio_addrchk_datal(6)
    );
  rx_input_memio_addrchk_datal_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_7_FFY_RST
    );
  rx_input_memio_addrchk_datal_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_7_FFX_RST,
      O => rx_input_memio_addrchk_datal(7)
    );
  rx_input_memio_addrchk_datal_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_7_FFX_RST
    );
  rx_input_fifo_control_cs_FFd4_1872 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_fifo_control_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_control_cs_FFd4_FFY_SET,
      RST => GND,
      O => rx_input_fifo_control_cs_FFd4
    );
  rx_input_fifo_control_cs_FFd4_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF_2,
      O => rx_input_fifo_control_cs_FFd4_FFY_SET
    );
  rx_input_memio_addrchk_datal_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_9_FFY_RST,
      O => rx_input_memio_addrchk_datal(8)
    );
  rx_input_memio_addrchk_datal_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_9_FFY_RST
    );
  rx_input_memio_addrchk_datal_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_9_FFX_RST,
      O => rx_input_memio_addrchk_datal(9)
    );
  rx_input_memio_addrchk_datal_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_9_FFX_RST
    );
  rx_fifocheck_fbbpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(0),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_1_FFY_RST,
      O => rx_fifocheck_fbbpl(0)
    );
  rx_fifocheck_fbbpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_1_FFY_RST
    );
  tx_input_dl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(15),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_15_FFX_RST,
      O => tx_input_dl(15)
    );
  tx_input_dl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_15_FFX_RST
    );
  tx_input_bp_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_30,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_15_FFY_RST,
      O => txbp(14)
    );
  txbp_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_15_FFY_RST
    );
  tx_input_bp_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_31,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_15_FFX_RST,
      O => txbp(15)
    );
  txbp_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_15_FFX_RST
    );
  rx_input_memio_addrchk_rxucastl_1873 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxucast,
      CE => rx_input_memio_addrchk_rxucastl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_rxucastl_FFY_RST,
      O => rx_input_memio_addrchk_rxucastl
    );
  rx_input_memio_addrchk_rxucastl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_rxucastl_FFY_RST
    );
  rx_input_memio_addrchk_cs_FFd1_1874 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd1_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd1_FFY_RST,
      O => rx_input_memio_addrchk_cs_FFd1
    );
  rx_input_memio_addrchk_cs_FFd1_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd1_FFY_RST
    );
  mac_control_lmacaddr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_11_FFX_RST,
      O => mac_control_lmacaddr(11)
    );
  mac_control_lmacaddr_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_11_FFX_RST
    );
  mac_control_lmacaddr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_11_FFY_RST,
      O => mac_control_lmacaddr(10)
    );
  mac_control_lmacaddr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_11_FFY_RST
    );
  mac_control_lmacaddr_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_13_FFY_RST,
      O => mac_control_lmacaddr(12)
    );
  mac_control_lmacaddr_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_13_FFY_RST
    );
  mac_control_lmacaddr_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_21_FFY_RST,
      O => mac_control_lmacaddr(20)
    );
  mac_control_lmacaddr_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_21_FFY_RST
    );
  mac_control_lmacaddr_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_21_FFX_RST,
      O => mac_control_lmacaddr(21)
    );
  mac_control_lmacaddr_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_21_FFX_RST
    );
  mac_control_lmacaddr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_13_FFX_RST,
      O => mac_control_lmacaddr(13)
    );
  mac_control_lmacaddr_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_13_FFX_RST
    );
  mac_control_lmacaddr_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_23_FFY_RST,
      O => mac_control_lmacaddr(22)
    );
  mac_control_lmacaddr_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_23_FFY_RST
    );
  mac_control_lmacaddr_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_23_FFX_RST,
      O => mac_control_lmacaddr(23)
    );
  mac_control_lmacaddr_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_23_FFX_RST
    );
  mac_control_lmacaddr_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_31_FFY_RST,
      O => mac_control_lmacaddr(30)
    );
  mac_control_lmacaddr_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_31_FFY_RST
    );
  rx_input_memio_addrchk_datal_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_27_FFX_RST,
      O => rx_input_memio_addrchk_datal(27)
    );
  rx_input_memio_addrchk_datal_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_27_FFX_RST
    );
  rx_input_memio_addrchk_datal_34 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_35_FFY_RST,
      O => rx_input_memio_addrchk_datal(34)
    );
  rx_input_memio_addrchk_datal_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_35_FFY_RST
    );
  rx_input_memio_addrchk_datal_35 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_35_FFX_RST,
      O => rx_input_memio_addrchk_datal(35)
    );
  rx_input_memio_addrchk_datal_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_35_FFX_RST
    );
  rx_input_memio_addrchk_datal_42 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_43_FFY_RST,
      O => rx_input_memio_addrchk_datal(42)
    );
  rx_input_memio_addrchk_datal_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_43_FFY_RST
    );
  rx_input_memio_addrchk_datal_43 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_43_FFX_RST,
      O => rx_input_memio_addrchk_datal(43)
    );
  rx_input_memio_addrchk_datal_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_43_FFX_RST
    );
  rx_input_memio_addrchk_datal_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_19_FFY_RST,
      O => rx_input_memio_addrchk_datal(18)
    );
  rx_input_memio_addrchk_datal_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_19_FFY_RST
    );
  rx_input_memio_addrchk_datal_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_19_FFX_RST,
      O => rx_input_memio_addrchk_datal(19)
    );
  rx_input_memio_addrchk_datal_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_19_FFX_RST
    );
  rx_input_memio_addrchk_datal_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_29_FFY_RST,
      O => rx_input_memio_addrchk_datal(28)
    );
  rx_input_memio_addrchk_datal_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_29_FFY_RST
    );
  rx_input_memio_addrchk_datal_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_29_FFX_RST,
      O => rx_input_memio_addrchk_datal(29)
    );
  rx_input_memio_addrchk_datal_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_29_FFX_RST
    );
  rx_input_memio_addrchk_datal_36 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_37_FFY_RST,
      O => rx_input_memio_addrchk_datal(36)
    );
  rx_input_memio_addrchk_datal_37_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_37_FFY_RST
    );
  rx_input_memio_addrchk_datal_37 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_37_FFX_RST,
      O => rx_input_memio_addrchk_datal(37)
    );
  rx_input_memio_addrchk_datal_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_37_FFX_RST
    );
  rx_input_memio_addrchk_datal_44 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_45_FFY_RST,
      O => rx_input_memio_addrchk_datal(44)
    );
  rx_input_memio_addrchk_datal_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_45_FFY_RST
    );
  rx_input_memio_addrchk_datal_45 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_45_FFX_RST,
      O => rx_input_memio_addrchk_datal(45)
    );
  rx_input_memio_addrchk_datal_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_45_FFX_RST
    );
  rx_input_memio_addrchk_datal_38 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_39_FFY_RST,
      O => rx_input_memio_addrchk_datal(38)
    );
  rx_input_memio_addrchk_datal_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_39_FFY_RST
    );
  rx_input_memio_addrchk_datal_39 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_39_FFX_RST,
      O => rx_input_memio_addrchk_datal(39)
    );
  rx_input_memio_addrchk_datal_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_39_FFX_RST
    );
  rx_input_memio_addrchk_datal_46 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_47_FFY_RST,
      O => rx_input_memio_addrchk_datal(46)
    );
  rx_input_memio_addrchk_datal_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_47_FFY_RST
    );
  rx_fifocheck_fbbpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(1),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_1_FFX_RST,
      O => rx_fifocheck_fbbpl(1)
    );
  rx_fifocheck_fbbpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_1_FFX_RST
    );
  rx_fifocheck_fbbpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(2),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_3_FFY_RST,
      O => rx_fifocheck_fbbpl(2)
    );
  rx_fifocheck_fbbpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_3_FFY_RST
    );
  rx_fifocheck_fbbpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(3),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_3_FFX_RST,
      O => rx_fifocheck_fbbpl(3)
    );
  rx_fifocheck_fbbpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_3_FFX_RST
    );
  rx_fifocheck_fbbpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(4),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_5_FFY_RST,
      O => rx_fifocheck_fbbpl(4)
    );
  rx_fifocheck_fbbpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_5_FFY_RST
    );
  rx_fifocheck_fbbpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(5),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_5_FFX_RST,
      O => rx_fifocheck_fbbpl(5)
    );
  rx_fifocheck_fbbpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_5_FFX_RST
    );
  rx_fifocheck_fbbpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(6),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_7_FFY_RST,
      O => rx_fifocheck_fbbpl(6)
    );
  rx_fifocheck_fbbpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_7_FFY_RST
    );
  rx_fifocheck_fbbpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(7),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_7_FFX_RST,
      O => rx_fifocheck_fbbpl(7)
    );
  rx_fifocheck_fbbpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_7_FFX_RST
    );
  rx_fifocheck_fbbpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(8),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_9_FFY_RST,
      O => rx_fifocheck_fbbpl(8)
    );
  rx_fifocheck_fbbpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_9_FFY_RST
    );
  rx_fifocheck_fbbpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(9),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_9_FFX_RST,
      O => rx_fifocheck_fbbpl(9)
    );
  rx_fifocheck_fbbpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_9_FFX_RST
    );
  mac_control_txfifowerr_cntl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(0),
      CE => mac_control_txfifowerr_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_1_FFY_RST,
      O => mac_control_txfifowerr_cntl(0)
    );
  mac_control_txfifowerr_cntl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_1_FFY_RST
    );
  mac_control_txfifowerr_cntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(1),
      CE => mac_control_txfifowerr_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_1_FFX_RST,
      O => mac_control_txfifowerr_cntl(1)
    );
  mac_control_txfifowerr_cntl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_1_FFX_RST
    );
  mac_control_txfifowerr_cntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(2),
      CE => mac_control_txfifowerr_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_3_FFY_RST,
      O => mac_control_txfifowerr_cntl(2)
    );
  mac_control_txfifowerr_cntl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_3_FFY_RST
    );
  mac_control_txfifowerr_cntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(3),
      CE => mac_control_txfifowerr_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_3_FFX_RST,
      O => mac_control_txfifowerr_cntl(3)
    );
  mac_control_txfifowerr_cntl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_3_FFX_RST
    );
  mac_control_txfifowerr_cntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(4),
      CE => mac_control_txfifowerr_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_5_FFY_RST,
      O => mac_control_txfifowerr_cntl(4)
    );
  mac_control_txfifowerr_cntl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_5_FFY_RST
    );
  rx_input_memio_cs_FFd1_1875 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd2,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd1_FFY_RST,
      O => rx_input_memio_cs_FFd1
    );
  rx_input_memio_cs_FFd1_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd1_FFY_RST
    );
  mac_control_txfifowerr_cntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txfifowerr_cnt(5),
      CE => mac_control_txfifowerr_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txfifowerr_cntl_5_FFX_RST,
      O => mac_control_txfifowerr_cntl(5)
    );
  mac_control_txfifowerr_cntl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txfifowerr_cntl_5_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(1),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_1_FFX_RST,
      O => mac_control_phydo(1)
    );
  mac_control_phydo_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_1_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(3),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_3_FFX_RST,
      O => mac_control_phydo(3)
    );
  mac_control_phydo_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_3_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(4),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_5_FFY_RST,
      O => mac_control_phydo(4)
    );
  mac_control_phydo_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_5_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(5),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_5_FFX_RST,
      O => mac_control_phydo(5)
    );
  mac_control_phydo_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_5_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(6),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_7_FFY_RST,
      O => mac_control_phydo(6)
    );
  mac_control_phydo_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_7_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(7),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_7_FFX_RST,
      O => mac_control_phydo(7)
    );
  mac_control_phydo_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_7_FFX_RST
    );
  mac_control_PHY_status_PHYDOUT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(8),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_9_FFY_RST,
      O => mac_control_phydo(8)
    );
  mac_control_phydo_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_9_FFY_RST
    );
  mac_control_PHY_status_PHYDOUT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_dout(9),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_phydo_9_FFX_RST,
      O => mac_control_phydo(9)
    );
  mac_control_phydo_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydo_9_FFX_RST
    );
  rx_input_memio_crcl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_8_1_O,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_8_FFY_RST,
      O => rx_input_memio_crcl(8)
    );
  rx_input_memio_crcl_8_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_8_FFY_RST
    );
  memcontroller_dnl2_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(11),
      CE => memcontroller_dnl2_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_11_FFX_RST,
      O => memcontroller_dnl2(11)
    );
  memcontroller_dnl2_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_11_FFX_RST
    );
  memcontroller_dnl2_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(10),
      CE => memcontroller_dnl2_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_11_FFY_RST,
      O => memcontroller_dnl2(10)
    );
  memcontroller_dnl2_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_11_FFY_RST
    );
  memcontroller_dnl2_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(20),
      CE => memcontroller_dnl2_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_21_FFY_RST,
      O => memcontroller_dnl2(20)
    );
  memcontroller_dnl2_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_21_FFY_RST
    );
  memcontroller_dnl2_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(21),
      CE => memcontroller_dnl2_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_21_FFX_RST,
      O => memcontroller_dnl2(21)
    );
  memcontroller_dnl2_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_21_FFX_RST
    );
  memcontroller_dnl2_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(12),
      CE => memcontroller_dnl2_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_13_FFY_RST,
      O => memcontroller_dnl2(12)
    );
  memcontroller_dnl2_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_13_FFY_RST
    );
  memcontroller_dnl2_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(19),
      CE => memcontroller_dnl2_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_19_FFX_RST,
      O => memcontroller_dnl2(19)
    );
  memcontroller_dnl2_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_19_FFX_RST
    );
  memcontroller_dnl2_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(28),
      CE => memcontroller_dnl2_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_29_FFY_RST,
      O => memcontroller_dnl2(28)
    );
  memcontroller_dnl2_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_29_FFY_RST
    );
  memcontroller_dnl2_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(29),
      CE => memcontroller_dnl2_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_29_FFX_RST,
      O => memcontroller_dnl2(29)
    );
  memcontroller_dnl2_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_29_FFX_RST
    );
  rx_input_memio_datal_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_datal_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_1_FFY_RST,
      O => rx_input_memio_datal(0)
    );
  rx_input_memio_datal_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_1_FFY_RST
    );
  rx_input_memio_datal_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_datal_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_1_FFX_RST,
      O => rx_input_memio_datal(1)
    );
  rx_input_memio_datal_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_1_FFX_RST
    );
  rx_input_memio_datal_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_datal_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_3_FFY_RST,
      O => rx_input_memio_datal(2)
    );
  rx_input_memio_datal_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_3_FFY_RST
    );
  rx_input_memio_datal_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_datal_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_3_FFX_RST,
      O => rx_input_memio_datal(3)
    );
  rx_input_memio_datal_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_3_FFX_RST
    );
  rx_input_memio_datal_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_datal_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_5_FFY_RST,
      O => rx_input_memio_datal(4)
    );
  rx_input_memio_datal_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_5_FFY_RST
    );
  rx_input_memio_datal_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_datal_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_5_FFX_RST,
      O => rx_input_memio_datal(5)
    );
  rx_input_memio_datal_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_5_FFX_RST
    );
  rx_input_memio_datal_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_datal_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_7_FFY_RST,
      O => rx_input_memio_datal(6)
    );
  rx_input_memio_datal_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_7_FFY_RST
    );
  rx_input_memio_datal_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_datal_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_datal_7_FFX_RST,
      O => rx_input_memio_datal(7)
    );
  rx_input_memio_datal_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_datal_7_FFX_RST
    );
  rx_input_memio_addrchk_maceq_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq(1),
      CE => rx_input_memio_addrchk_maceq_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_0_FFY_RST,
      O => rx_input_memio_addrchk_maceq(1)
    );
  rx_input_memio_addrchk_maceq_0_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_0_FFY_RST
    );
  rx_input_memio_addrchk_maceq_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq_0_rt,
      CE => rx_input_memio_addrchk_maceq_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_0_FFX_RST,
      O => rx_input_memio_addrchk_maceq(0)
    );
  rx_input_memio_addrchk_maceq_0_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_0_FFX_RST
    );
  memcontroller_dnl2_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(13),
      CE => memcontroller_dnl2_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_13_FFX_RST,
      O => memcontroller_dnl2(13)
    );
  memcontroller_dnl2_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_13_FFX_RST
    );
  memcontroller_dnl2_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(22),
      CE => memcontroller_dnl2_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_23_FFY_RST,
      O => memcontroller_dnl2(22)
    );
  memcontroller_dnl2_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_23_FFY_RST
    );
  memcontroller_dnl2_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(23),
      CE => memcontroller_dnl2_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_23_FFX_RST,
      O => memcontroller_dnl2(23)
    );
  memcontroller_dnl2_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_23_FFX_RST
    );
  memcontroller_dnl2_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(14),
      CE => memcontroller_dnl2_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_15_FFY_RST,
      O => memcontroller_dnl2(14)
    );
  memcontroller_dnl2_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_15_FFY_RST
    );
  memcontroller_dnl2_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(15),
      CE => memcontroller_dnl2_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_15_FFX_RST,
      O => memcontroller_dnl2(15)
    );
  memcontroller_dnl2_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_15_FFX_RST
    );
  memcontroller_dnl2_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(30),
      CE => memcontroller_dnl2_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_31_FFY_RST,
      O => memcontroller_dnl2(30)
    );
  memcontroller_dnl2_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_31_FFY_RST
    );
  memcontroller_dnl2_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(31),
      CE => memcontroller_dnl2_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_31_FFX_RST,
      O => memcontroller_dnl2(31)
    );
  memcontroller_dnl2_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_31_FFX_RST
    );
  memcontroller_dnl2_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(24),
      CE => memcontroller_dnl2_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_25_FFY_RST,
      O => memcontroller_dnl2(24)
    );
  memcontroller_dnl2_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_25_FFY_RST
    );
  memcontroller_dnl2_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(25),
      CE => memcontroller_dnl2_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_25_FFX_RST,
      O => memcontroller_dnl2(25)
    );
  memcontroller_dnl2_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_25_FFX_RST
    );
  memcontroller_dnl2_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(16),
      CE => memcontroller_dnl2_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_17_FFY_RST,
      O => memcontroller_dnl2(16)
    );
  memcontroller_dnl2_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_17_FFY_RST
    );
  memcontroller_dnl2_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(17),
      CE => memcontroller_dnl2_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_17_FFX_RST,
      O => memcontroller_dnl2(17)
    );
  memcontroller_dnl2_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_17_FFX_RST
    );
  memcontroller_dnl2_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(26),
      CE => memcontroller_dnl2_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_27_FFY_RST,
      O => memcontroller_dnl2(26)
    );
  memcontroller_dnl2_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_27_FFY_RST
    );
  memcontroller_dnl2_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(27),
      CE => memcontroller_dnl2_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_27_FFX_RST,
      O => memcontroller_dnl2(27)
    );
  memcontroller_dnl2_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_27_FFX_RST
    );
  memcontroller_dnl2_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_dnl1(18),
      CE => memcontroller_dnl2_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_dnl2_19_FFY_RST,
      O => memcontroller_dnl2(18)
    );
  memcontroller_dnl2_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_dnl2_19_FFY_RST
    );
  rx_input_memio_crcl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_9_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_9_FFY_RST,
      O => rx_input_memio_crcl(9)
    );
  rx_input_memio_crcl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_9_FFY_RST
    );
  mac_control_sclkdeltall_1876 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_sclkdeltal,
      CE => mac_control_sclkdeltall_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_sclkdeltall_FFY_RST,
      O => mac_control_sclkdeltall
    );
  mac_control_sclkdeltall_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_sclkdeltall_FFY_RST
    );
  mac_control_phyaddr_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_11_FFY_RST,
      O => mac_control_phyaddr(10)
    );
  mac_control_phyaddr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_11_FFY_RST
    );
  mac_control_phyaddr_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_11_FFX_RST,
      O => mac_control_phyaddr(11)
    );
  mac_control_phyaddr_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_11_FFX_RST
    );
  mac_control_phyaddr_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_13_FFX_RST,
      O => mac_control_phyaddr(13)
    );
  mac_control_phyaddr_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_13_FFX_RST
    );
  mac_control_phyaddr_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(21),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_21_FFX_RST,
      O => mac_control_phyaddr(21)
    );
  mac_control_phyaddr_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_21_FFX_RST
    );
  mac_control_phyaddr_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(22),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_23_FFY_RST,
      O => mac_control_phyaddr(22)
    );
  mac_control_phyaddr_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_23_FFY_RST
    );
  mac_control_phyaddr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_15_FFX_RST,
      O => mac_control_phyaddr(15)
    );
  mac_control_phyaddr_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_15_FFX_RST
    );
  rx_input_memio_addrchk_datal_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_13_FFX_RST,
      O => rx_input_memio_addrchk_datal(13)
    );
  rx_input_memio_addrchk_datal_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_13_FFX_RST
    );
  rx_input_memio_addrchk_datal_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_23_FFY_RST,
      O => rx_input_memio_addrchk_datal(22)
    );
  rx_input_memio_addrchk_datal_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_23_FFY_RST
    );
  rx_input_memio_addrchk_datal_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_31_FFY_RST,
      O => rx_input_memio_addrchk_datal(30)
    );
  rx_input_memio_addrchk_datal_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_31_FFY_RST
    );
  rx_input_memio_addrchk_datal_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_31_FFX_RST,
      O => rx_input_memio_addrchk_datal(31)
    );
  rx_input_memio_addrchk_datal_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_31_FFX_RST
    );
  rx_input_memio_addrchk_datal_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_23_FFX_RST,
      O => rx_input_memio_addrchk_datal(23)
    );
  rx_input_memio_addrchk_datal_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_23_FFX_RST
    );
  rx_input_memio_addrchk_datal_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_15_FFY_RST,
      O => rx_input_memio_addrchk_datal(14)
    );
  rx_input_memio_addrchk_datal_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_15_FFY_RST
    );
  rx_input_memio_addrchk_datal_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_15_FFX_RST,
      O => rx_input_memio_addrchk_datal(15)
    );
  rx_input_memio_addrchk_datal_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_15_FFX_RST
    );
  rx_input_memio_addrchk_datal_40 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_41_FFY_RST,
      O => rx_input_memio_addrchk_datal(40)
    );
  rx_input_memio_addrchk_datal_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_41_FFY_RST
    );
  rx_input_memio_addrchk_datal_32 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_33_FFY_RST,
      O => rx_input_memio_addrchk_datal(32)
    );
  rx_input_memio_addrchk_datal_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_33_FFY_RST
    );
  rx_input_memio_addrchk_datal_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_25_FFY_RST,
      O => rx_input_memio_addrchk_datal(24)
    );
  rx_input_memio_addrchk_datal_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_25_FFY_RST
    );
  rx_input_memio_addrchk_datal_33 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0028,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_33_FFX_RST,
      O => rx_input_memio_addrchk_datal(33)
    );
  rx_input_memio_addrchk_datal_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_33_FFX_RST
    );
  rx_input_memio_addrchk_datal_41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0027,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_41_FFX_RST,
      O => rx_input_memio_addrchk_datal(41)
    );
  rx_input_memio_addrchk_datal_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_41_FFX_RST
    );
  rx_input_memio_addrchk_datal_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_25_FFX_RST,
      O => rx_input_memio_addrchk_datal(25)
    );
  rx_input_memio_addrchk_datal_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_25_FFX_RST
    );
  rx_input_memio_addrchk_datal_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_17_FFY_RST,
      O => rx_input_memio_addrchk_datal(16)
    );
  rx_input_memio_addrchk_datal_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_17_FFY_RST
    );
  rx_input_memio_addrchk_datal_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_addrchk_n0029,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_27_FFY_RST,
      O => rx_input_memio_addrchk_datal(26)
    );
  rx_input_memio_addrchk_datal_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_27_FFY_RST
    );
  rx_input_memio_addrchk_datal_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_17_FFX_RST,
      O => rx_input_memio_addrchk_datal(17)
    );
  rx_input_memio_addrchk_datal_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_17_FFX_RST
    );
  rx_input_memio_addrchk_maceq_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq_2_rt,
      CE => rx_input_memio_addrchk_maceq_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_2_FFX_RST,
      O => rx_input_memio_addrchk_maceq(2)
    );
  rx_input_memio_addrchk_maceq_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_2_FFX_RST
    );
  rx_input_memio_addrchk_maceq_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_lmaceq_4_rt,
      CE => rx_input_memio_addrchk_maceq_4_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_maceq_4_FFX_RST,
      O => rx_input_memio_addrchk_maceq(4)
    );
  rx_input_memio_addrchk_maceq_4_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_maceq_4_FFX_RST
    );
  tx_output_crcl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_24_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_24_FFY_RST,
      O => tx_output_crcl(24)
    );
  tx_output_crcl_24_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_24_FFY_RST
    );
  tx_output_crcl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_16_1_O,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_16_FFY_RST,
      O => tx_output_crcl(16)
    );
  tx_output_crcl_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_16_FFY_RST
    );
  rx_input_memio_crcl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_11_1_O,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_11_FFY_RST,
      O => rx_input_memio_crcl(11)
    );
  rx_input_memio_crcl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_11_FFY_RST
    );
  rx_fifocheck_fbbpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_11_FFX_RST,
      O => rx_fifocheck_fbbpl(11)
    );
  rx_fifocheck_fbbpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_11_FFX_RST
    );
  rx_fifocheck_fbbpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_13_FFY_RST,
      O => rx_fifocheck_fbbpl(12)
    );
  rx_fifocheck_fbbpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_13_FFY_RST
    );
  rx_fifocheck_fbbpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_13_FFX_RST,
      O => rx_fifocheck_fbbpl(13)
    );
  rx_fifocheck_fbbpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_13_FFX_RST
    );
  rx_fifocheck_fbbpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_15_FFY_RST,
      O => rx_fifocheck_fbbpl(14)
    );
  rx_fifocheck_fbbpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_15_FFY_RST
    );
  rx_fifocheck_fbbpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfbbp(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_fifocheck_fbbpl_15_FFX_RST,
      O => rx_fifocheck_fbbpl(15)
    );
  rx_fifocheck_fbbpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_fifocheck_fbbpl_15_FFX_RST
    );
  rx_input_memio_dout_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_11_FFY_RST,
      O => rx_input_memio_dout(10)
    );
  rx_input_memio_dout_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_11_FFY_RST
    );
  rx_input_memio_dout_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_11_FFX_RST,
      O => rx_input_memio_dout(11)
    );
  rx_input_memio_dout_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_11_FFX_RST
    );
  rx_input_memio_dout_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_n0046,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_21_FFX_RST,
      O => rx_input_memio_dout(21)
    );
  rx_input_memio_dout_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_21_FFX_RST
    );
  rx_input_memio_dout_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_n0045,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_13_FFX_RST,
      O => rx_input_memio_dout(13)
    );
  rx_input_memio_dout_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_13_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_dreg_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(11),
      CE => mac_control_PHY_status_MII_Interface_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_MII_Interface_dreg_12_FFX_RST,
      O => mac_control_PHY_status_MII_Interface_dreg(12)
    );
  mac_control_PHY_status_MII_Interface_dreg_12_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_MII_Interface_dreg_12_FFX_RST
    );
  rx_input_memio_dout_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(6),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_31_FFY_RST,
      O => rx_input_memio_dout(30)
    );
  rx_input_memio_dout_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_31_FFY_RST
    );
  rx_input_memio_dout_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(7),
      CE => rx_input_memio_n0047,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_dout_31_FFX_RST,
      O => rx_input_memio_dout(31)
    );
  rx_input_memio_dout_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_dout_31_FFX_RST
    );
  mac_control_phyaddr_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(16),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_17_FFY_RST,
      O => mac_control_phyaddr(16)
    );
  mac_control_phyaddr_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_17_FFY_RST
    );
  mac_control_phyaddr_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(23),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_23_FFX_RST,
      O => mac_control_phyaddr(23)
    );
  mac_control_phyaddr_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_23_FFX_RST
    );
  mac_control_phyaddr_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(17),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_17_FFX_RST,
      O => mac_control_phyaddr(17)
    );
  mac_control_phyaddr_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_17_FFX_RST
    );
  mac_control_phyaddr_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(25),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_25_FFX_RST,
      O => mac_control_phyaddr(25)
    );
  mac_control_phyaddr_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_25_FFX_RST
    );
  mac_control_phyaddr_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(19),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_19_FFX_RST,
      O => mac_control_phyaddr(19)
    );
  mac_control_phyaddr_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_19_FFX_RST
    );
  mac_control_phyaddr_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(27),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_27_FFX_RST,
      O => mac_control_phyaddr(27)
    );
  mac_control_phyaddr_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_27_FFX_RST
    );
  mac_control_phyaddr_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(29),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_29_FFX_RST,
      O => mac_control_phyaddr(29)
    );
  mac_control_phyaddr_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_29_FFX_RST
    );
  rx_input_memio_addrchk_datal_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(3),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_11_FFX_RST,
      O => rx_input_memio_addrchk_datal(11)
    );
  rx_input_memio_addrchk_datal_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_11_FFX_RST
    );
  rx_input_memio_addrchk_datal_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0031,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_13_FFY_RST,
      O => rx_input_memio_addrchk_datal(12)
    );
  rx_input_memio_addrchk_datal_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_13_FFY_RST
    );
  rx_input_memio_addrchk_datal_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(4),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_21_FFY_RST,
      O => rx_input_memio_addrchk_datal(20)
    );
  rx_input_memio_addrchk_datal_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_21_FFY_RST
    );
  rx_input_memio_addrchk_datal_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(5),
      CE => rx_input_memio_addrchk_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_datal_21_FFX_RST,
      O => rx_input_memio_addrchk_datal(21)
    );
  rx_input_memio_addrchk_datal_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_datal_21_FFX_RST
    );
  tx_output_bpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(3),
      CE => tx_output_bpl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_3_FFX_RST,
      O => tx_output_bpl(3)
    );
  tx_output_bpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_3_FFX_RST
    );
  tx_output_bpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(4),
      CE => tx_output_bpl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_5_FFY_RST,
      O => tx_output_bpl(4)
    );
  tx_output_bpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_5_FFY_RST
    );
  tx_output_bpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(5),
      CE => tx_output_bpl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_5_FFX_RST,
      O => tx_output_bpl(5)
    );
  tx_output_bpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_5_FFX_RST
    );
  tx_output_bpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(6),
      CE => tx_output_bpl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_7_FFY_RST,
      O => tx_output_bpl(6)
    );
  tx_output_bpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_7_FFY_RST
    );
  tx_output_bpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(7),
      CE => tx_output_bpl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_7_FFX_RST,
      O => tx_output_bpl(7)
    );
  tx_output_bpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_7_FFX_RST
    );
  tx_output_bpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(8),
      CE => tx_output_bpl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_9_FFY_RST,
      O => tx_output_bpl(8)
    );
  tx_output_bpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_9_FFY_RST
    );
  tx_output_bpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(9),
      CE => tx_output_bpl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_9_FFX_RST,
      O => tx_output_bpl(9)
    );
  tx_output_bpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_9_FFX_RST
    );
  mac_control_MACADDR_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_11_FFY_RST,
      O => macaddr(10)
    );
  macaddr_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_11_FFY_RST
    );
  mac_control_MACADDR_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_11_FFX_RST,
      O => macaddr(11)
    );
  macaddr_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_11_FFX_RST
    );
  mac_control_MACADDR_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_13_FFX_RST,
      O => macaddr(13)
    );
  macaddr_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_13_FFX_RST
    );
  mac_control_MACADDR_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(21),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_21_FFX_RST,
      O => macaddr(21)
    );
  macaddr_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_21_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(19),
      CE => rx_input_memio_addrchk_macaddrl_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_19_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(19)
    );
  rx_input_memio_addrchk_macaddrl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_19_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_45 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(45),
      CE => rx_input_memio_addrchk_macaddrl_45_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_45_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(45)
    );
  rx_input_memio_addrchk_macaddrl_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_45_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_37 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(37),
      CE => rx_input_memio_addrchk_macaddrl_37_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_37_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(37)
    );
  rx_input_memio_addrchk_macaddrl_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_37_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(29),
      CE => rx_input_memio_addrchk_macaddrl_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_29_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(29)
    );
  rx_input_memio_addrchk_macaddrl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_29_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(47),
      CE => rx_input_memio_addrchk_macaddrl_47_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_47_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(47)
    );
  rx_input_memio_addrchk_macaddrl_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_47_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_39 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(39),
      CE => rx_input_memio_addrchk_macaddrl_39_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_39_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(39)
    );
  rx_input_memio_addrchk_macaddrl_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_39_FFX_RST
    );
  mac_control_phydi_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_1_FFX_RST,
      O => mac_control_phydi(1)
    );
  mac_control_phydi_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_1_FFX_RST
    );
  mac_control_phydi_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_1_FFY_RST,
      O => mac_control_phydi(0)
    );
  mac_control_phydi_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_1_FFY_RST
    );
  rx_input_memio_addrchk_validucast_1877 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_n0052,
      CE => rx_input_memio_addrchk_validucast_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_validucast_FFY_RST,
      O => rx_input_memio_addrchk_validucast
    );
  rx_input_memio_addrchk_validucast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_validucast_FFY_RST
    );
  mac_control_phydi_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_3_FFX_RST,
      O => mac_control_phydi(3)
    );
  mac_control_phydi_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_3_FFX_RST
    );
  mac_control_phydi_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_3_FFY_RST,
      O => mac_control_phydi(2)
    );
  mac_control_phydi_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_3_FFY_RST
    );
  mac_control_phydi_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_5_FFY_RST,
      O => mac_control_phydi(4)
    );
  mac_control_phydi_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_5_FFY_RST
    );
  mac_control_phydi_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_5_FFX_RST,
      O => mac_control_phydi(5)
    );
  mac_control_phydi_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_5_FFX_RST
    );
  mac_control_phydi_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_7_FFY_RST,
      O => mac_control_phydi(6)
    );
  mac_control_phydi_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_7_FFY_RST
    );
  mac_control_phydi_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_7_FFX_RST,
      O => mac_control_phydi(7)
    );
  mac_control_phydi_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_7_FFX_RST
    );
  mac_control_phydi_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_9_FFY_RST,
      O => mac_control_phydi(8)
    );
  mac_control_phydi_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_9_FFY_RST
    );
  mac_control_phydi_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_9_FFX_RST,
      O => mac_control_phydi(9)
    );
  mac_control_phydi_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_9_FFX_RST
    );
  rx_input_memio_bpen_1878 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd2,
      CE => rx_input_memio_bpen_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpen_FFY_RST,
      O => rx_input_memio_bpen
    );
  rx_input_memio_bpen_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpen_FFY_RST
    );
  rx_input_memio_addrchk_DESTOK : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_n0053,
      CE => rx_input_memio_destok_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_destok_FFY_RST,
      O => rx_input_memio_destok
    );
  rx_input_memio_destok_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_destok_FFY_RST
    );
  rx_output_cs_FFd10_1879 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd10_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd10_FFY_RST,
      O => rx_output_cs_FFd10
    );
  rx_output_cs_FFd10_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd10_FFY_RST
    );
  tx_output_crcl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_18_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_18_FFY_RST,
      O => tx_output_crcl(18)
    );
  tx_output_crcl_18_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_18_FFY_RST
    );
  tx_output_crcl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_26_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_26_FFY_RST,
      O => tx_output_crcl(26)
    );
  tx_output_crcl_26_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_26_FFY_RST
    );
  rx_input_memio_doutl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(1),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_1_FFX_RST,
      O => rx_input_memio_doutl(1)
    );
  rx_input_memio_doutl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_1_FFX_RST
    );
  rx_input_memio_doutl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(0),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_1_FFY_RST,
      O => rx_input_memio_doutl(0)
    );
  rx_input_memio_doutl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_1_FFY_RST
    );
  rx_input_memio_doutl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(2),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_2_FFY_RST,
      O => rx_input_memio_doutl(2)
    );
  rx_input_memio_doutl_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_2_FFY_RST
    );
  rx_input_memio_doutl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(3),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_3_FFY_RST,
      O => rx_input_memio_doutl(3)
    );
  rx_input_memio_doutl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_3_FFY_RST
    );
  rx_input_memio_doutl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(4),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_5_FFY_RST,
      O => rx_input_memio_doutl(4)
    );
  rx_input_memio_doutl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_5_FFY_RST
    );
  mac_control_lrxallf_1880 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0014,
      CLK => mac_control_CLKSL_5,
      SET => mac_control_lrxallf_FFY_SET,
      RST => GND,
      O => mac_control_lrxallf
    );
  mac_control_lrxallf_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => mac_control_lrxallf_FFY_SET
    );
  rx_input_memio_doutl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(6),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_7_FFY_RST,
      O => rx_input_memio_doutl(6)
    );
  rx_input_memio_doutl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_7_FFY_RST
    );
  rx_input_memio_doutl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(5),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_5_FFX_RST,
      O => rx_input_memio_doutl(5)
    );
  rx_input_memio_doutl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_5_FFX_RST
    );
  rx_input_memio_crcl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_14_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_14_FFY_RST,
      O => rx_input_memio_crcl(14)
    );
  rx_input_memio_crcl_14_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_14_FFY_RST
    );
  tx_input_cs_FFd12_1881 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => tx_input_cs_FFd12_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => tx_input_cs_FFd12_FFY_SET,
      RST => GND,
      O => tx_input_cs_FFd12
    );
  tx_input_cs_FFd12_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF_1,
      O => tx_input_cs_FFd12_FFY_SET
    );
  mac_control_rxcrcerr_cntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(1),
      CE => mac_control_rxcrcerr_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_1_FFX_RST,
      O => mac_control_rxcrcerr_cntl(1)
    );
  mac_control_rxcrcerr_cntl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_1_FFX_RST
    );
  mac_control_rxcrcerr_cntl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(0),
      CE => mac_control_rxcrcerr_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_1_FFY_RST,
      O => mac_control_rxcrcerr_cntl(0)
    );
  mac_control_rxcrcerr_cntl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_1_FFY_RST
    );
  mac_control_rxcrcerr_cntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(2),
      CE => mac_control_rxcrcerr_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_3_FFY_RST,
      O => mac_control_rxcrcerr_cntl(2)
    );
  mac_control_rxcrcerr_cntl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_3_FFY_RST
    );
  mac_control_rxcrcerr_cntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(3),
      CE => mac_control_rxcrcerr_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_3_FFX_RST,
      O => mac_control_rxcrcerr_cntl(3)
    );
  mac_control_rxcrcerr_cntl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_3_FFX_RST
    );
  mac_control_rxcrcerr_cntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(4),
      CE => mac_control_rxcrcerr_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_5_FFY_RST,
      O => mac_control_rxcrcerr_cntl(4)
    );
  mac_control_rxcrcerr_cntl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_5_FFY_RST
    );
  mac_control_rxcrcerr_cntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(5),
      CE => mac_control_rxcrcerr_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_5_FFX_RST,
      O => mac_control_rxcrcerr_cntl(5)
    );
  mac_control_rxcrcerr_cntl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_5_FFX_RST
    );
  mac_control_rxcrcerr_cntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(6),
      CE => mac_control_rxcrcerr_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_7_FFY_RST,
      O => mac_control_rxcrcerr_cntl(6)
    );
  mac_control_rxcrcerr_cntl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_7_FFY_RST
    );
  mac_control_rxcrcerr_cntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(7),
      CE => mac_control_rxcrcerr_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_7_FFX_RST,
      O => mac_control_rxcrcerr_cntl(7)
    );
  mac_control_rxcrcerr_cntl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_7_FFX_RST
    );
  mac_control_rxcrcerr_cntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(8),
      CE => mac_control_rxcrcerr_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_9_FFY_RST,
      O => mac_control_rxcrcerr_cntl(8)
    );
  mac_control_rxcrcerr_cntl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_9_FFY_RST
    );
  mac_control_rxcrcerr_cntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(9),
      CE => mac_control_rxcrcerr_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_9_FFX_RST,
      O => mac_control_rxcrcerr_cntl(9)
    );
  mac_control_rxcrcerr_cntl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_9_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(10),
      CE => rx_input_memio_addrchk_macaddrl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_11_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(10)
    );
  rx_input_memio_addrchk_macaddrl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_11_FFY_RST
    );
  rx_input_memio_addrchk_macaddrl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(11),
      CE => rx_input_memio_addrchk_macaddrl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_11_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(11)
    );
  rx_input_memio_addrchk_macaddrl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_11_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(21),
      CE => rx_input_memio_addrchk_macaddrl_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_21_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(21)
    );
  rx_input_memio_addrchk_macaddrl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_21_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(13),
      CE => rx_input_memio_addrchk_macaddrl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_13_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(13)
    );
  rx_input_memio_addrchk_macaddrl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_13_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(31),
      CE => rx_input_memio_addrchk_macaddrl_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_31_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(31)
    );
  rx_input_memio_addrchk_macaddrl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_31_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(23),
      CE => rx_input_memio_addrchk_macaddrl_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_23_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(23)
    );
  rx_input_memio_addrchk_macaddrl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_23_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(15),
      CE => rx_input_memio_addrchk_macaddrl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_15_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(15)
    );
  rx_input_memio_addrchk_macaddrl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_15_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_40 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(40),
      CE => rx_input_memio_addrchk_macaddrl_41_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_41_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(40)
    );
  rx_input_memio_addrchk_macaddrl_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_41_FFY_RST
    );
  mac_control_PHY_status_phyaddrws_1882 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_phyaddrws_BYMUXNOT,
      CE => mac_control_PHY_status_n00151_O,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_phyaddrws_FFY_RST,
      O => mac_control_PHY_status_phyaddrws
    );
  mac_control_PHY_status_phyaddrws_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_phyaddrws_FFY_RST
    );
  mac_control_dout_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0016(31),
      CE => mac_control_n0012,
      CLK => clksl,
      SET => GND,
      RST => mac_control_dout_31_FFY_RST,
      O => mac_control_dout(31)
    );
  mac_control_dout_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_dout_31_FFY_RST
    );
  mac_control_rxcrcerr_rst_1883 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_n0052,
      CE => mac_control_rxcrcerr_rst_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_rst_FFY_RST,
      O => mac_control_rxcrcerr_rst
    );
  mac_control_rxcrcerr_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_rst_FFY_RST
    );
  tx_output_bpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(0),
      CE => tx_output_bpl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_1_FFY_RST,
      O => tx_output_bpl(0)
    );
  tx_output_bpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_1_FFY_RST
    );
  tx_output_bpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(2),
      CE => tx_output_bpl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_3_FFY_RST,
      O => tx_output_bpl(2)
    );
  tx_output_bpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_3_FFY_RST
    );
  tx_output_bpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(1),
      CE => tx_output_bpl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_1_FFX_RST,
      O => tx_output_bpl(1)
    );
  tx_output_bpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_1_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(41),
      CE => rx_input_memio_addrchk_macaddrl_41_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_41_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(41)
    );
  rx_input_memio_addrchk_macaddrl_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_41_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_33 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(33),
      CE => rx_input_memio_addrchk_macaddrl_33_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_33_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(33)
    );
  rx_input_memio_addrchk_macaddrl_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_33_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(25),
      CE => rx_input_memio_addrchk_macaddrl_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_25_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(25)
    );
  rx_input_memio_addrchk_macaddrl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_25_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(17),
      CE => rx_input_memio_addrchk_macaddrl_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_17_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(17)
    );
  rx_input_memio_addrchk_macaddrl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_17_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_43 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(43),
      CE => rx_input_memio_addrchk_macaddrl_43_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_43_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(43)
    );
  rx_input_memio_addrchk_macaddrl_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_43_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_35 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(35),
      CE => rx_input_memio_addrchk_macaddrl_35_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_35_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(35)
    );
  rx_input_memio_addrchk_macaddrl_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_35_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(27),
      CE => rx_input_memio_addrchk_macaddrl_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_27_FFX_RST,
      O => rx_input_memio_addrchk_macaddrl(27)
    );
  rx_input_memio_addrchk_macaddrl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_27_FFX_RST
    );
  rx_input_memio_addrchk_macaddrl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => macaddr(18),
      CE => rx_input_memio_addrchk_macaddrl_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_macaddrl_19_FFY_RST,
      O => rx_input_memio_addrchk_macaddrl(18)
    );
  rx_input_memio_addrchk_macaddrl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_macaddrl_19_FFY_RST
    );
  tx_output_crcl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_28_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_28_FFY_RST,
      O => tx_output_crcl(28)
    );
  tx_output_crcl_28_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_28_FFY_RST
    );
  rx_input_memio_crcl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_23_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_23_FFY_RST,
      O => rx_input_memio_crcl(23)
    );
  rx_input_memio_crcl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_23_FFY_RST
    );
  rx_input_memio_addrchk_rxallfl_1884 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxallf,
      CE => rx_input_memio_addrchk_rxallfl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_rxallfl_FFY_RST,
      O => rx_input_memio_addrchk_rxallfl
    );
  rx_input_memio_addrchk_rxallfl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_rxallfl_FFY_RST
    );
  rx_input_memio_crcll_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(13),
      CE => rx_input_memio_crcll_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_13_FFX_RST,
      O => rx_input_memio_crcll(13)
    );
  rx_input_memio_crcll_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_13_FFX_RST
    );
  rx_input_memio_crcll_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(20),
      CE => rx_input_memio_crcll_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_21_FFY_RST,
      O => rx_input_memio_crcll(20)
    );
  rx_input_memio_crcll_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_21_FFY_RST
    );
  rx_input_memio_crcll_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(21),
      CE => rx_input_memio_crcll_21_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_21_FFX_RST,
      O => rx_input_memio_crcll(21)
    );
  rx_input_memio_crcll_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_21_FFX_RST
    );
  rx_input_memio_crcll_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(14),
      CE => rx_input_memio_crcll_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_15_FFY_RST,
      O => rx_input_memio_crcll(14)
    );
  rx_input_memio_crcll_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_15_FFY_RST
    );
  rx_input_memio_crcll_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(15),
      CE => rx_input_memio_crcll_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_15_FFX_RST,
      O => rx_input_memio_crcll(15)
    );
  rx_input_memio_crcll_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_15_FFX_RST
    );
  rx_input_memio_crcll_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(30),
      CE => rx_input_memio_crcll_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_31_FFY_RST,
      O => rx_input_memio_crcll(30)
    );
  rx_input_memio_crcll_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_31_FFY_RST
    );
  rx_input_memio_crcll_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(31),
      CE => rx_input_memio_crcll_31_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_31_FFX_RST,
      O => rx_input_memio_crcll(31)
    );
  rx_input_memio_crcll_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_31_FFX_RST
    );
  rx_input_memio_crcll_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(22),
      CE => rx_input_memio_crcll_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_23_FFY_RST,
      O => rx_input_memio_crcll(22)
    );
  rx_input_memio_crcll_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_23_FFY_RST
    );
  rx_input_memio_crcll_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(23),
      CE => rx_input_memio_crcll_23_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_23_FFX_RST,
      O => rx_input_memio_crcll(23)
    );
  rx_input_memio_crcll_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_23_FFX_RST
    );
  rx_input_memio_crcll_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(16),
      CE => rx_input_memio_crcll_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_17_FFY_RST,
      O => rx_input_memio_crcll(16)
    );
  rx_input_memio_crcll_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_17_FFY_RST
    );
  rx_input_memio_crcll_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(17),
      CE => rx_input_memio_crcll_17_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_17_FFX_RST,
      O => rx_input_memio_crcll(17)
    );
  rx_input_memio_crcll_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_17_FFX_RST
    );
  rx_input_memio_crcll_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(26),
      CE => rx_input_memio_crcll_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_27_FFY_RST,
      O => rx_input_memio_crcll(26)
    );
  rx_input_memio_crcll_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_27_FFY_RST
    );
  rx_input_memio_crcll_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(25),
      CE => rx_input_memio_crcll_25_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_25_FFX_RST,
      O => rx_input_memio_crcll(25)
    );
  rx_input_memio_crcll_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_25_FFX_RST
    );
  mac_control_PHY_status_addrl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(1),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_addrl_1_FFX_RST,
      O => mac_control_PHY_status_addrl(1)
    );
  mac_control_PHY_status_addrl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_addrl_1_FFX_RST
    );
  mac_control_PHY_status_addrl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(3),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_addrl_3_FFX_RST,
      O => mac_control_PHY_status_addrl(3)
    );
  mac_control_PHY_status_addrl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_addrl_3_FFX_RST
    );
  tx_output_outsell_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_outsel_1_Q,
      CE => tx_output_outsell_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outsell_1_FFY_RST,
      O => tx_output_outsell(1)
    );
  tx_output_outsell_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outsell_1_FFY_RST
    );
  mac_control_din_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_1_FFX_RST,
      O => mac_control_din(1)
    );
  mac_control_din_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_1_FFX_RST
    );
  rx_input_memio_crcl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_17_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_17_FFY_RST,
      O => rx_input_memio_crcl(17)
    );
  rx_input_memio_crcl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_17_FFY_RST
    );
  mac_control_din_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_Mshreg_sinlll_102,
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_1_FFY_RST,
      O => mac_control_din(0)
    );
  mac_control_din_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_1_FFY_RST
    );
  mac_control_din_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_3_FFY_RST,
      O => mac_control_din(2)
    );
  mac_control_din_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_3_FFY_RST
    );
  mac_control_din_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_3_FFX_RST,
      O => mac_control_din(3)
    );
  mac_control_din_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_3_FFX_RST
    );
  mac_control_din_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_5_FFY_RST,
      O => mac_control_din(4)
    );
  mac_control_din_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_5_FFY_RST
    );
  mac_control_din_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_7_FFY_RST,
      O => mac_control_din(6)
    );
  mac_control_din_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_7_FFY_RST
    );
  mac_control_din_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_5_FFX_RST,
      O => mac_control_din(5)
    );
  mac_control_din_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_5_FFX_RST
    );
  mac_control_rxcrcerr_cntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(11),
      CE => mac_control_rxcrcerr_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_11_FFX_RST,
      O => mac_control_rxcrcerr_cntl(11)
    );
  mac_control_rxcrcerr_cntl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_11_FFX_RST
    );
  mac_control_rxcrcerr_cntl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(20),
      CE => mac_control_rxcrcerr_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_21_FFY_RST,
      O => mac_control_rxcrcerr_cntl(20)
    );
  mac_control_rxcrcerr_cntl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_21_FFY_RST
    );
  mac_control_rxcrcerr_cntl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(21),
      CE => mac_control_rxcrcerr_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_21_FFX_RST,
      O => mac_control_rxcrcerr_cntl(21)
    );
  mac_control_rxcrcerr_cntl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_21_FFX_RST
    );
  mac_control_rxcrcerr_cntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(12),
      CE => mac_control_rxcrcerr_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_13_FFY_RST,
      O => mac_control_rxcrcerr_cntl(12)
    );
  mac_control_rxcrcerr_cntl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_13_FFY_RST
    );
  mac_control_rxcrcerr_cntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(13),
      CE => mac_control_rxcrcerr_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_13_FFX_RST,
      O => mac_control_rxcrcerr_cntl(13)
    );
  mac_control_rxcrcerr_cntl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_13_FFX_RST
    );
  mac_control_rxcrcerr_cntl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(22),
      CE => mac_control_rxcrcerr_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_23_FFY_RST,
      O => mac_control_rxcrcerr_cntl(22)
    );
  mac_control_rxcrcerr_cntl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_23_FFY_RST
    );
  mac_control_rxcrcerr_cntl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(23),
      CE => mac_control_rxcrcerr_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_23_FFX_RST,
      O => mac_control_rxcrcerr_cntl(23)
    );
  mac_control_rxcrcerr_cntl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_23_FFX_RST
    );
  mac_control_rxcrcerr_cntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(14),
      CE => mac_control_rxcrcerr_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_15_FFY_RST,
      O => mac_control_rxcrcerr_cntl(14)
    );
  mac_control_rxcrcerr_cntl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_15_FFY_RST
    );
  mac_control_rxcrcerr_cntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(15),
      CE => mac_control_rxcrcerr_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_15_FFX_RST,
      O => mac_control_rxcrcerr_cntl(15)
    );
  mac_control_rxcrcerr_cntl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_15_FFX_RST
    );
  mac_control_rxcrcerr_cntl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(30),
      CE => mac_control_rxcrcerr_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_31_FFY_RST,
      O => mac_control_rxcrcerr_cntl(30)
    );
  mac_control_rxcrcerr_cntl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_31_FFY_RST
    );
  mac_control_rxcrcerr_cntl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(31),
      CE => mac_control_rxcrcerr_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_31_FFX_RST,
      O => mac_control_rxcrcerr_cntl(31)
    );
  mac_control_rxcrcerr_cntl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_31_FFX_RST
    );
  mac_control_rxcrcerr_cntl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(16),
      CE => mac_control_rxcrcerr_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_17_FFY_RST,
      O => mac_control_rxcrcerr_cntl(16)
    );
  mac_control_rxcrcerr_cntl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_17_FFY_RST
    );
  mac_control_rxcrcerr_cntl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(24),
      CE => mac_control_rxcrcerr_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_25_FFY_RST,
      O => mac_control_rxcrcerr_cntl(24)
    );
  mac_control_rxcrcerr_cntl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_25_FFY_RST
    );
  mac_control_rxcrcerr_cntl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(17),
      CE => mac_control_rxcrcerr_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_17_FFX_RST,
      O => mac_control_rxcrcerr_cntl(17)
    );
  mac_control_rxcrcerr_cntl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_17_FFX_RST
    );
  mac_control_lrxmcast_1885 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0026,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lrxmcast_FFY_RST,
      O => mac_control_lrxmcast
    );
  mac_control_lrxmcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lrxmcast_FFY_RST
    );
  mac_control_rxoferr_cntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(10),
      CE => mac_control_rxoferr_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_11_FFY_RST,
      O => mac_control_rxoferr_cntl(10)
    );
  mac_control_rxoferr_cntl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_11_FFY_RST
    );
  mac_control_rxoferr_cntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(11),
      CE => mac_control_rxoferr_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_11_FFX_RST,
      O => mac_control_rxoferr_cntl(11)
    );
  mac_control_rxoferr_cntl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_11_FFX_RST
    );
  mac_control_rxoferr_cntl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(20),
      CE => mac_control_rxoferr_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_21_FFY_RST,
      O => mac_control_rxoferr_cntl(20)
    );
  mac_control_rxoferr_cntl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_21_FFY_RST
    );
  mac_control_rxoferr_cntl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(21),
      CE => mac_control_rxoferr_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_21_FFX_RST,
      O => mac_control_rxoferr_cntl(21)
    );
  mac_control_rxoferr_cntl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_21_FFX_RST
    );
  mac_control_rxoferr_cntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(12),
      CE => mac_control_rxoferr_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_13_FFY_RST,
      O => mac_control_rxoferr_cntl(12)
    );
  mac_control_rxoferr_cntl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_13_FFY_RST
    );
  mac_control_rxoferr_cntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(13),
      CE => mac_control_rxoferr_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_13_FFX_RST,
      O => mac_control_rxoferr_cntl(13)
    );
  mac_control_rxoferr_cntl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_13_FFX_RST
    );
  mac_control_rxoferr_cntl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(30),
      CE => mac_control_rxoferr_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_31_FFY_RST,
      O => mac_control_rxoferr_cntl(30)
    );
  mac_control_rxoferr_cntl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_31_FFY_RST
    );
  mac_control_rxoferr_cntl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(31),
      CE => mac_control_rxoferr_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_31_FFX_RST,
      O => mac_control_rxoferr_cntl(31)
    );
  mac_control_rxoferr_cntl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_31_FFX_RST
    );
  mac_control_rxoferr_cntl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(22),
      CE => mac_control_rxoferr_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_23_FFY_RST,
      O => mac_control_rxoferr_cntl(22)
    );
  mac_control_rxoferr_cntl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_23_FFY_RST
    );
  mac_control_rxoferr_cntl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(23),
      CE => mac_control_rxoferr_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_23_FFX_RST,
      O => mac_control_rxoferr_cntl(23)
    );
  mac_control_rxoferr_cntl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_23_FFX_RST
    );
  mac_control_rxoferr_cntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(14),
      CE => mac_control_rxoferr_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_15_FFY_RST,
      O => mac_control_rxoferr_cntl(14)
    );
  mac_control_rxoferr_cntl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_15_FFY_RST
    );
  mac_control_rxoferr_cntl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(24),
      CE => mac_control_rxoferr_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_25_FFY_RST,
      O => mac_control_rxoferr_cntl(24)
    );
  mac_control_rxoferr_cntl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_25_FFY_RST
    );
  mac_control_rxoferr_cntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(15),
      CE => mac_control_rxoferr_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_15_FFX_RST,
      O => mac_control_rxoferr_cntl(15)
    );
  mac_control_rxoferr_cntl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_15_FFX_RST
    );
  rx_input_memio_crcll_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(27),
      CE => rx_input_memio_crcll_27_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_27_FFX_RST,
      O => rx_input_memio_crcll(27)
    );
  rx_input_memio_crcll_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_27_FFX_RST
    );
  rx_input_memio_crcll_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(18),
      CE => rx_input_memio_crcll_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_19_FFY_RST,
      O => rx_input_memio_crcll(18)
    );
  rx_input_memio_crcll_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_19_FFY_RST
    );
  rx_input_memio_crcll_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(28),
      CE => rx_input_memio_crcll_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_29_FFY_RST,
      O => rx_input_memio_crcll(28)
    );
  rx_input_memio_crcll_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_29_FFY_RST
    );
  rx_input_memio_crcll_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(19),
      CE => rx_input_memio_crcll_19_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_19_FFX_RST,
      O => rx_input_memio_crcll(19)
    );
  rx_input_memio_crcll_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_19_FFX_RST
    );
  rx_input_memio_crcll_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_crcl(29),
      CE => rx_input_memio_crcll_29_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcll_29_FFX_RST,
      O => rx_input_memio_crcll(29)
    );
  rx_input_memio_crcll_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcll_29_FFX_RST
    );
  rx_input_memio_crcl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_24_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_24_FFY_RST,
      O => rx_input_memio_crcl(24)
    );
  rx_input_memio_crcl_24_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_24_FFY_RST
    );
  rx_input_memio_crcl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_16_1_O,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_16_FFY_RST,
      O => rx_input_memio_crcl(16)
    );
  rx_input_memio_crcl_16_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_16_FFY_RST
    );
  mac_control_din_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_7_FFX_RST,
      O => mac_control_din(7)
    );
  mac_control_din_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_7_FFX_RST
    );
  tx_output_outsell_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => tx_output_outsel_0_Q,
      CE => tx_output_outsell_0_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => tx_output_outsell_0_FFY_SET,
      RST => GND,
      O => tx_output_outsell(0)
    );
  tx_output_outsell_0_FFY_SETOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outsell_0_FFY_SET
    );
  memcontroller_oel_1886 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_oel_BYMUXNOT,
      CE => memcontroller_oel_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_oel_FFY_RST,
      O => memcontroller_oel
    );
  memcontroller_oel_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_oel_FFY_RST
    );
  mac_control_din_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_9_FFY_RST,
      O => mac_control_din(8)
    );
  mac_control_din_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_9_FFY_RST
    );
  mac_control_din_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_9_FFX_RST,
      O => mac_control_din(9)
    );
  mac_control_din_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_9_FFX_RST
    );
  rx_input_memio_macnt_72_1887 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_macnt_inst_sum_221,
      CE => rx_input_memio_n0101,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_macnt_72_FFY_RST,
      O => rx_input_memio_macnt_72
    );
  rx_input_memio_macnt_72_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_macnt_72_FFY_RST
    );
  rx_output_cs_FFd18_1888 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_cs_FFd18_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_cs_FFd18_FFY_RST,
      O => rx_output_cs_FFd18
    );
  rx_output_cs_FFd18_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => rx_output_cs_FFd18_FFY_RST
    );
  mac_control_phydi_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_11_FFY_RST,
      O => mac_control_phydi(10)
    );
  mac_control_phydi_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_11_FFY_RST
    );
  mac_control_phydi_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(20),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_21_FFY_RST,
      O => mac_control_phydi(20)
    );
  mac_control_phydi_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_21_FFY_RST
    );
  mac_control_phydi_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_11_FFX_RST,
      O => mac_control_phydi(11)
    );
  mac_control_phydi_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_11_FFX_RST
    );
  mac_control_MACADDR_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(31),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_31_FFX_RST,
      O => macaddr(31)
    );
  macaddr_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_31_FFX_RST
    );
  mac_control_MACADDR_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(23),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_23_FFX_RST,
      O => macaddr(23)
    );
  macaddr_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_23_FFX_RST
    );
  mac_control_MACADDR_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_15_FFX_RST,
      O => macaddr(15)
    );
  macaddr_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_15_FFX_RST
    );
  mac_control_MACADDR_33 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(33),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_33_FFX_RST,
      O => macaddr(33)
    );
  macaddr_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_33_FFX_RST
    );
  mac_control_MACADDR_41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(41),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_41_FFX_RST,
      O => macaddr(41)
    );
  macaddr_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_41_FFX_RST
    );
  mac_control_MACADDR_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(25),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_25_FFX_RST,
      O => macaddr(25)
    );
  macaddr_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_25_FFX_RST
    );
  mac_control_MACADDR_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(17),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_17_FFX_RST,
      O => macaddr(17)
    );
  macaddr_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_17_FFX_RST
    );
  mac_control_MACADDR_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(27),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_27_FFX_RST,
      O => macaddr(27)
    );
  macaddr_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_27_FFX_RST
    );
  mac_control_MACADDR_42 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(42),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_43_FFY_RST,
      O => macaddr(42)
    );
  macaddr_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_43_FFY_RST
    );
  mac_control_din_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(20),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_21_FFX_RST,
      O => mac_control_din(21)
    );
  mac_control_din_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_21_FFX_RST
    );
  mac_control_din_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_15_FFY_RST,
      O => mac_control_din(14)
    );
  mac_control_din_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_15_FFY_RST
    );
  mac_control_din_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_15_FFX_RST,
      O => mac_control_din(15)
    );
  mac_control_din_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_15_FFX_RST
    );
  mac_control_din_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(21),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_23_FFY_RST,
      O => mac_control_din(22)
    );
  mac_control_din_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_23_FFY_RST
    );
  mac_control_din_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(22),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_23_FFX_RST,
      O => mac_control_din(23)
    );
  mac_control_din_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_23_FFX_RST
    );
  mac_control_din_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(29),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_31_FFY_RST,
      O => mac_control_din(30)
    );
  mac_control_din_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_31_FFY_RST
    );
  mac_control_din_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(30),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_31_FFX_RST,
      O => mac_control_din(31)
    );
  mac_control_din_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_31_FFX_RST
    );
  mac_control_din_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_17_FFY_RST,
      O => mac_control_din(16)
    );
  mac_control_din_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_17_FFY_RST
    );
  mac_control_din_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(16),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_17_FFX_RST,
      O => mac_control_din(17)
    );
  mac_control_din_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_17_FFX_RST
    );
  mac_control_din_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(23),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_25_FFY_RST,
      O => mac_control_din(24)
    );
  mac_control_din_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_25_FFY_RST
    );
  mac_control_din_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(24),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_25_FFX_RST,
      O => mac_control_din(25)
    );
  mac_control_din_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_25_FFX_RST
    );
  mac_control_din_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(17),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_19_FFY_RST,
      O => mac_control_din(18)
    );
  mac_control_din_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_19_FFY_RST
    );
  mac_control_din_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(18),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_19_FFX_RST,
      O => mac_control_din(19)
    );
  mac_control_din_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_19_FFX_RST
    );
  mac_control_din_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(25),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_27_FFY_RST,
      O => mac_control_din(26)
    );
  mac_control_din_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_27_FFY_RST
    );
  mac_control_din_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(26),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_27_FFX_RST,
      O => mac_control_din(27)
    );
  mac_control_din_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_27_FFX_RST
    );
  mac_control_din_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(27),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_29_FFY_RST,
      O => mac_control_din(28)
    );
  mac_control_din_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_29_FFY_RST
    );
  mac_control_MACADDR_35 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(35),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_35_FFX_RST,
      O => macaddr(35)
    );
  macaddr_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_35_FFX_RST
    );
  mac_control_MACADDR_43 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(43),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_43_FFX_RST,
      O => macaddr(43)
    );
  macaddr_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_43_FFX_RST
    );
  mac_control_MACADDR_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(19),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_19_FFX_RST,
      O => macaddr(19)
    );
  macaddr_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_19_FFX_RST
    );
  mac_control_MACADDR_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(29),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_29_FFX_RST,
      O => macaddr(29)
    );
  macaddr_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_29_FFX_RST
    );
  mac_control_MACADDR_37 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(37),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_37_FFX_RST,
      O => macaddr(37)
    );
  macaddr_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_37_FFX_RST
    );
  mac_control_MACADDR_45 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(45),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_45_FFX_RST,
      O => macaddr(45)
    );
  macaddr_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_45_FFX_RST
    );
  mac_control_MACADDR_39 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(39),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_39_FFX_RST,
      O => macaddr(39)
    );
  macaddr_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_39_FFX_RST
    );
  mac_control_MACADDR_47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_lmacaddr(47),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => macaddr_47_FFX_RST,
      O => macaddr(47)
    );
  macaddr_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => macaddr_47_FFX_RST
    );
  mac_control_PHY_status_addrl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phyaddr(2),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_addrl_3_FFY_RST,
      O => mac_control_PHY_status_addrl(2)
    );
  mac_control_PHY_status_addrl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_addrl_3_FFY_RST
    );
  rx_input_memio_addrchk_rxmcastl_1889 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxmcast,
      CE => rx_input_memio_addrchk_rxmcastl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_rxmcastl_FFY_RST,
      O => rx_input_memio_addrchk_rxmcastl
    );
  rx_input_memio_addrchk_rxmcastl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_rxmcastl_FFY_RST
    );
  rx_input_fifo_control_dinl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(0),
      CE => rx_input_fifo_control_dinl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_1_FFY_RST,
      O => rx_input_fifo_control_dinl(0)
    );
  rx_input_fifo_control_dinl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_1_FFY_RST
    );
  rx_input_fifo_control_dinl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(1),
      CE => rx_input_fifo_control_dinl_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_1_FFX_RST,
      O => rx_input_fifo_control_dinl(1)
    );
  rx_input_fifo_control_dinl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_1_FFX_RST
    );
  rx_input_fifo_control_dinl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(2),
      CE => rx_input_fifo_control_dinl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_3_FFY_RST,
      O => rx_input_fifo_control_dinl(2)
    );
  rx_input_fifo_control_dinl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_3_FFY_RST
    );
  rx_input_fifo_control_dinl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(3),
      CE => rx_input_fifo_control_dinl_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_3_FFX_RST,
      O => rx_input_fifo_control_dinl(3)
    );
  rx_input_fifo_control_dinl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_3_FFX_RST
    );
  rx_input_fifo_control_dinl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(4),
      CE => rx_input_fifo_control_dinl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_5_FFY_RST,
      O => rx_input_fifo_control_dinl(4)
    );
  rx_input_fifo_control_dinl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_5_FFY_RST
    );
  rx_input_fifo_control_dinl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(5),
      CE => rx_input_fifo_control_dinl_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_5_FFX_RST,
      O => rx_input_fifo_control_dinl(5)
    );
  rx_input_fifo_control_dinl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_5_FFX_RST
    );
  rx_input_fifo_control_dinl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(6),
      CE => rx_input_fifo_control_dinl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_7_FFY_RST,
      O => rx_input_fifo_control_dinl(6)
    );
  rx_input_fifo_control_dinl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_7_FFY_RST
    );
  rx_input_fifo_control_dinl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(7),
      CE => rx_input_fifo_control_dinl_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_7_FFX_RST,
      O => rx_input_fifo_control_dinl(7)
    );
  rx_input_fifo_control_dinl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_7_FFX_RST
    );
  rx_input_fifo_control_dinl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_fifodout(8),
      CE => rx_input_fifo_control_dinl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_9_FFY_RST,
      O => rx_input_fifo_control_dinl(8)
    );
  rx_input_fifo_control_dinl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_9_FFY_RST
    );
  rx_input_fifo_control_dinl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_dout(9),
      CE => rx_input_fifo_control_dinl_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_dinl_9_FFX_RST,
      O => rx_input_fifo_control_dinl(9)
    );
  rx_input_fifo_control_dinl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_dinl_9_FFX_RST
    );
  mac_control_phydi_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(21),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_21_FFX_RST,
      O => mac_control_phydi(21)
    );
  mac_control_phydi_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_21_FFX_RST
    );
  mac_control_phydi_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_13_FFY_RST,
      O => mac_control_phydi(12)
    );
  mac_control_phydi_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_13_FFY_RST
    );
  mac_control_phydi_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_13_FFX_RST,
      O => mac_control_phydi(13)
    );
  mac_control_phydi_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_13_FFX_RST
    );
  mac_control_phydi_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(22),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_23_FFY_RST,
      O => mac_control_phydi(22)
    );
  mac_control_phydi_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_23_FFY_RST
    );
  mac_control_phydi_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(30),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_31_FFY_RST,
      O => mac_control_phydi(30)
    );
  mac_control_phydi_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_31_FFY_RST
    );
  mac_control_phydi_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(31),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_31_FFX_RST,
      O => mac_control_phydi(31)
    );
  mac_control_phydi_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_31_FFX_RST
    );
  mac_control_phydi_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(23),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_23_FFX_RST,
      O => mac_control_phydi(23)
    );
  mac_control_phydi_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_23_FFX_RST
    );
  mac_control_phydi_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_15_FFY_RST,
      O => mac_control_phydi(14)
    );
  mac_control_phydi_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_15_FFY_RST
    );
  mac_control_phydi_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_15_FFX_RST,
      O => mac_control_phydi(15)
    );
  mac_control_phydi_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_15_FFX_RST
    );
  mac_control_phydi_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(24),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_25_FFY_RST,
      O => mac_control_phydi(24)
    );
  mac_control_phydi_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_25_FFY_RST
    );
  mac_control_phydi_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(25),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_25_FFX_RST,
      O => mac_control_phydi(25)
    );
  mac_control_phydi_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_25_FFX_RST
    );
  mac_control_phydi_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(16),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_17_FFY_RST,
      O => mac_control_phydi(16)
    );
  mac_control_phydi_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_17_FFY_RST
    );
  mac_control_phydi_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(17),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_17_FFX_RST,
      O => mac_control_phydi(17)
    );
  mac_control_phydi_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_17_FFX_RST
    );
  mac_control_phydi_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(26),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_27_FFY_RST,
      O => mac_control_phydi(26)
    );
  mac_control_phydi_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_27_FFY_RST
    );
  mac_control_phydi_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(27),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_27_FFX_RST,
      O => mac_control_phydi(27)
    );
  mac_control_phydi_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_27_FFX_RST
    );
  mac_control_phydi_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(18),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_19_FFY_RST,
      O => mac_control_phydi(18)
    );
  mac_control_phydi_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_19_FFY_RST
    );
  mac_control_phydi_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(19),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_19_FFX_RST,
      O => mac_control_phydi(19)
    );
  mac_control_phydi_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_19_FFX_RST
    );
  mac_control_phydi_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(28),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_29_FFY_RST,
      O => mac_control_phydi(28)
    );
  mac_control_phydi_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_29_FFY_RST
    );
  mac_control_phydi_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(29),
      CE => mac_control_n0013,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phydi_29_FFX_RST,
      O => mac_control_phydi(29)
    );
  mac_control_phydi_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phydi_29_FFX_RST
    );
  rx_input_memio_bpl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(0),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_1_FFY_RST,
      O => rx_input_memio_bpl(0)
    );
  rx_input_memio_bpl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_1_FFY_RST
    );
  rx_input_memio_bpl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(1),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_1_FFX_RST,
      O => rx_input_memio_bpl(1)
    );
  rx_input_memio_bpl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_1_FFX_RST
    );
  rx_input_memio_bpl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(2),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_3_FFY_RST,
      O => rx_input_memio_bpl(2)
    );
  rx_input_memio_bpl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_3_FFY_RST
    );
  rx_input_memio_bpl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(3),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_3_FFX_RST,
      O => rx_input_memio_bpl(3)
    );
  rx_input_memio_bpl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_3_FFX_RST
    );
  rx_input_memio_bpl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(4),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_5_FFY_RST,
      O => rx_input_memio_bpl(4)
    );
  rx_input_memio_bpl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_5_FFY_RST
    );
  rx_input_memio_bpl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(5),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_5_FFX_RST,
      O => rx_input_memio_bpl(5)
    );
  rx_input_memio_bpl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_5_FFX_RST
    );
  rx_input_memio_bpl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(6),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_7_FFY_RST,
      O => rx_input_memio_bpl(6)
    );
  rx_input_memio_bpl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_7_FFY_RST
    );
  rx_input_memio_bpl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(7),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_7_FFX_RST,
      O => rx_input_memio_bpl(7)
    );
  rx_input_memio_bpl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_7_FFX_RST
    );
  rx_input_memio_bpl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(8),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_9_FFY_RST,
      O => rx_input_memio_bpl(8)
    );
  rx_input_memio_bpl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_9_FFY_RST
    );
  rx_input_memio_bpl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(9),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_9_FFX_RST,
      O => rx_input_memio_bpl(9)
    );
  rx_input_memio_bpl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_9_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_cs_FFd6_1890 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_cs_FFd6_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => mac_control_PHY_status_MII_Interface_cs_FFd6_FFY_SET,
      RST => GND,
      O => mac_control_PHY_status_MII_Interface_cs_FFd6
    );
  mac_control_PHY_status_MII_Interface_cs_FFd6_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => RESET_IBUF,
      O => mac_control_PHY_status_MII_Interface_cs_FFd6_FFY_SET
    );
  rx_input_memio_addrchk_cs_FFd6_1891 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_cs_FFd6_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_cs_FFd6_FFY_RST,
      O => rx_input_memio_addrchk_cs_FFd6
    );
  rx_input_memio_addrchk_cs_FFd6_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_memio_RESET_1,
      I1 => GSR,
      O => rx_input_memio_addrchk_cs_FFd6_FFY_RST
    );
  mac_control_PHY_status_din_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(10),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_11_FFY_RST,
      O => mac_control_PHY_status_din(10)
    );
  mac_control_PHY_status_din_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_11_FFY_RST
    );
  mac_control_PHY_status_din_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(11),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_11_FFX_RST,
      O => mac_control_PHY_status_din(11)
    );
  mac_control_PHY_status_din_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_11_FFX_RST
    );
  mac_control_PHY_status_din_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(12),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_13_FFY_RST,
      O => mac_control_PHY_status_din(12)
    );
  mac_control_PHY_status_din_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_13_FFY_RST
    );
  mac_control_PHY_status_din_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(13),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_13_FFX_RST,
      O => mac_control_PHY_status_din(13)
    );
  mac_control_PHY_status_din_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_13_FFX_RST
    );
  mac_control_PHY_status_din_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(14),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_15_FFY_RST,
      O => mac_control_PHY_status_din(14)
    );
  mac_control_PHY_status_din_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_15_FFY_RST
    );
  mac_control_PHY_status_din_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_phydi(15),
      CE => mac_control_PHY_status_n0011,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_din_15_FFX_RST,
      O => mac_control_PHY_status_din(15)
    );
  mac_control_PHY_status_din_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_din_15_FFX_RST
    );
  rx_input_memio_crcl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_18_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_18_FFY_RST,
      O => rx_input_memio_crcl(18)
    );
  rx_input_memio_crcl_18_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_18_FFY_RST
    );
  rx_input_memio_crcl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_26_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_26_FFY_RST,
      O => rx_input_memio_crcl(26)
    );
  rx_input_memio_crcl_26_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_26_FFY_RST
    );
  memcontroller_clknum_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_clknum_1_BYMUXNOT,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_clknum_1_FFY_RST,
      O => memcontroller_clknum(0)
    );
  memcontroller_clknum_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_1_FFY_RST
    );
  memcontroller_clknum_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_n0149,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => memcontroller_clknum_1_FFX_RST,
      O => memcontroller_clknum(1)
    );
  memcontroller_clknum_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF,
      I1 => GSR,
      O => memcontroller_clknum_1_FFX_RST
    );
  tx_output_FBBP_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(0),
      CE => txfbbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_1_FFY_RST,
      O => txfbbp(0)
    );
  txfbbp_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_1_FFY_RST
    );
  tx_output_FBBP_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(2),
      CE => txfbbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_3_FFY_RST,
      O => txfbbp(2)
    );
  txfbbp_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_3_FFY_RST
    );
  mac_control_rxf_cntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(1),
      CE => mac_control_rxf_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_1_FFX_RST,
      O => mac_control_rxf_cntl(1)
    );
  mac_control_rxf_cntl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_1_FFX_RST
    );
  mac_control_rxf_cntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(2),
      CE => mac_control_rxf_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_3_FFY_RST,
      O => mac_control_rxf_cntl(2)
    );
  mac_control_rxf_cntl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_3_FFY_RST
    );
  mac_control_rxf_cntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(3),
      CE => mac_control_rxf_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_3_FFX_RST,
      O => mac_control_rxf_cntl(3)
    );
  mac_control_rxf_cntl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_3_FFX_RST
    );
  mac_control_rxf_cntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(4),
      CE => mac_control_rxf_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_5_FFY_RST,
      O => mac_control_rxf_cntl(4)
    );
  mac_control_rxf_cntl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_5_FFY_RST
    );
  mac_control_rxf_cntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(5),
      CE => mac_control_rxf_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_5_FFX_RST,
      O => mac_control_rxf_cntl(5)
    );
  mac_control_rxf_cntl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_5_FFX_RST
    );
  mac_control_rxf_cntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(6),
      CE => mac_control_rxf_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_7_FFY_RST,
      O => mac_control_rxf_cntl(6)
    );
  mac_control_rxf_cntl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_7_FFY_RST
    );
  mac_control_rxf_cntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(7),
      CE => mac_control_rxf_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_7_FFX_RST,
      O => mac_control_rxf_cntl(7)
    );
  mac_control_rxf_cntl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_7_FFX_RST
    );
  mac_control_rxf_cntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(8),
      CE => mac_control_rxf_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_9_FFY_RST,
      O => mac_control_rxf_cntl(8)
    );
  mac_control_rxf_cntl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_9_FFY_RST
    );
  mac_control_rxf_cntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(9),
      CE => mac_control_rxf_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_9_FFX_RST,
      O => mac_control_rxf_cntl(9)
    );
  mac_control_rxf_cntl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_9_FFX_RST
    );
  rx_input_memio_addrchk_rxbcastl_1892 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxbcast,
      CE => rx_input_memio_addrchk_rxbcastl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_rxbcastl_FFY_RST,
      O => rx_input_memio_addrchk_rxbcastl
    );
  rx_input_memio_addrchk_rxbcastl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_rxbcastl_FFY_RST
    );
  mac_control_rxphyerr_cntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(10),
      CE => mac_control_rxphyerr_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_11_FFY_RST,
      O => mac_control_rxphyerr_cntl(10)
    );
  mac_control_rxphyerr_cntl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_11_FFY_RST
    );
  mac_control_rxphyerr_cntl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(11),
      CE => mac_control_rxphyerr_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_11_FFX_RST,
      O => mac_control_rxphyerr_cntl(11)
    );
  mac_control_rxphyerr_cntl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_11_FFX_RST
    );
  mac_control_rxphyerr_cntl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(20),
      CE => mac_control_rxphyerr_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_21_FFY_RST,
      O => mac_control_rxphyerr_cntl(20)
    );
  mac_control_rxphyerr_cntl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_21_FFY_RST
    );
  tx_output_FBBP_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(1),
      CE => txfbbp_1_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_1_FFX_RST,
      O => txfbbp(1)
    );
  txfbbp_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_1_FFX_RST
    );
  tx_output_FBBP_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(3),
      CE => txfbbp_3_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_3_FFX_RST,
      O => txfbbp(3)
    );
  txfbbp_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_3_FFX_RST
    );
  tx_output_FBBP_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(4),
      CE => txfbbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_5_FFY_RST,
      O => txfbbp(4)
    );
  txfbbp_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_5_FFY_RST
    );
  tx_output_FBBP_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(5),
      CE => txfbbp_5_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_5_FFX_RST,
      O => txfbbp(5)
    );
  txfbbp_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_5_FFX_RST
    );
  tx_output_FBBP_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(6),
      CE => txfbbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_7_FFY_RST,
      O => txfbbp(6)
    );
  txfbbp_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_7_FFY_RST
    );
  tx_output_FBBP_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(7),
      CE => txfbbp_7_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_7_FFX_RST,
      O => txfbbp(7)
    );
  txfbbp_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_7_FFX_RST
    );
  tx_output_FBBP_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(8),
      CE => txfbbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_9_FFY_RST,
      O => txfbbp(8)
    );
  txfbbp_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_9_FFY_RST
    );
  tx_output_FBBP_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => addr2ext(9),
      CE => txfbbp_9_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txfbbp_9_FFX_RST,
      O => txfbbp(9)
    );
  txfbbp_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txfbbp_9_FFX_RST
    );
  rx_input_memio_doutl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(10),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_11_FFY_RST,
      O => rx_input_memio_doutl(10)
    );
  rx_input_memio_doutl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_11_FFY_RST
    );
  rx_input_memio_doutl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(11),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_11_FFX_RST,
      O => rx_input_memio_doutl(11)
    );
  rx_input_memio_doutl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_11_FFX_RST
    );
  mac_control_lrxbcast_1893 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0025,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lrxbcast_FFY_RST,
      O => mac_control_lrxbcast
    );
  mac_control_lrxbcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lrxbcast_FFY_RST
    );
  rx_input_memio_doutl_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(20),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_21_FFY_RST,
      O => rx_input_memio_doutl(20)
    );
  rx_input_memio_doutl_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_21_FFY_RST
    );
  rx_input_memio_doutl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(21),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_21_FFX_RST,
      O => rx_input_memio_doutl(21)
    );
  rx_input_memio_doutl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_21_FFX_RST
    );
  rx_input_memio_doutl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(12),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_13_FFY_RST,
      O => rx_input_memio_doutl(12)
    );
  rx_input_memio_doutl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_13_FFY_RST
    );
  rx_input_fifo_control_d2_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(1),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_1_FFX_RST,
      O => rx_input_fifo_control_d2(1)
    );
  rx_input_fifo_control_d2_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_1_FFX_RST
    );
  rx_input_fifo_control_d1_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(6),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_7_FFY_RST,
      O => rx_input_fifo_control_d1(6)
    );
  rx_input_fifo_control_d1_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_7_FFY_RST
    );
  rx_input_fifo_control_d1_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(7),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_7_FFX_RST,
      O => rx_input_fifo_control_d1(7)
    );
  rx_input_fifo_control_d1_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_7_FFX_RST
    );
  rx_input_fifo_control_d2_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(2),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_3_FFY_RST,
      O => rx_input_fifo_control_d2(2)
    );
  rx_input_fifo_control_d2_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_3_FFY_RST
    );
  rx_input_fifo_control_d2_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(3),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_3_FFX_RST,
      O => rx_input_fifo_control_d2(3)
    );
  rx_input_fifo_control_d2_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_3_FFX_RST
    );
  rx_input_fifo_control_d2_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(4),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_5_FFY_RST,
      O => rx_input_fifo_control_d2(4)
    );
  rx_input_fifo_control_d2_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_5_FFY_RST
    );
  rx_input_fifo_control_d1_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0(8),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d1_8_FFY_RST,
      O => rx_input_fifo_control_d1(8)
    );
  rx_input_fifo_control_d1_8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d1_8_FFY_RST
    );
  rx_input_fifo_control_d2_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(5),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_5_FFX_RST,
      O => rx_input_fifo_control_d2(5)
    );
  rx_input_fifo_control_d2_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_5_FFX_RST
    );
  rx_input_fifo_control_d3_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(0),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_1_FFY_RST,
      O => rx_input_fifo_control_d3(0)
    );
  rx_input_fifo_control_d3_1_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_1_FFY_RST
    );
  rx_input_fifo_control_d3_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(1),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_1_FFX_RST,
      O => rx_input_fifo_control_d3(1)
    );
  rx_input_fifo_control_d3_1_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_1_FFX_RST
    );
  rx_input_fifo_control_d1_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d0_9_rt,
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_control_d1_9_FFY_SET,
      RST => rx_input_fifo_control_d1_9_FFY_RST,
      O => rx_input_fifo_control_d1(9)
    );
  rx_input_fifo_control_d1_9_FFY_SETOR : X_BUF
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_d1_9_FFY_SET
    );
  rx_input_fifo_control_d1_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_control_d1_9_LOGIC_ZERO,
      I1 => GSR,
      O => rx_input_fifo_control_d1_9_FFY_RST
    );
  rx_input_fifo_control_d2_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(6),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_7_FFY_RST,
      O => rx_input_fifo_control_d2(6)
    );
  rx_input_fifo_control_d2_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_7_FFY_RST
    );
  rx_input_memio_doutl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(13),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_13_FFX_RST,
      O => rx_input_memio_doutl(13)
    );
  rx_input_memio_doutl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_13_FFX_RST
    );
  rx_input_memio_doutl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(30),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_31_FFY_RST,
      O => rx_input_memio_doutl(30)
    );
  rx_input_memio_doutl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_31_FFY_RST
    );
  rx_input_memio_doutl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(31),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_31_FFX_RST,
      O => rx_input_memio_doutl(31)
    );
  rx_input_memio_doutl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_31_FFX_RST
    );
  rx_input_memio_doutl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(22),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_23_FFY_RST,
      O => rx_input_memio_doutl(22)
    );
  rx_input_memio_doutl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_23_FFY_RST
    );
  rx_input_memio_doutl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(23),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_23_FFX_RST,
      O => rx_input_memio_doutl(23)
    );
  rx_input_memio_doutl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_23_FFX_RST
    );
  rx_input_memio_doutl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(14),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_15_FFY_RST,
      O => rx_input_memio_doutl(14)
    );
  rx_input_memio_doutl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_15_FFY_RST
    );
  rx_input_memio_doutl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(15),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_15_FFX_RST,
      O => rx_input_memio_doutl(15)
    );
  rx_input_memio_doutl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_15_FFX_RST
    );
  rx_input_memio_doutl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(24),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_25_FFY_RST,
      O => rx_input_memio_doutl(24)
    );
  rx_input_memio_doutl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_25_FFY_RST
    );
  rx_input_memio_doutl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(25),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_25_FFX_RST,
      O => rx_input_memio_doutl(25)
    );
  rx_input_memio_doutl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_25_FFX_RST
    );
  rx_input_memio_doutl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(16),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_17_FFY_RST,
      O => rx_input_memio_doutl(16)
    );
  rx_input_memio_doutl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_17_FFY_RST
    );
  rx_input_memio_doutl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(17),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_17_FFX_RST,
      O => rx_input_memio_doutl(17)
    );
  rx_input_memio_doutl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_17_FFX_RST
    );
  rx_input_memio_doutl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(26),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_27_FFY_RST,
      O => rx_input_memio_doutl(26)
    );
  rx_input_memio_doutl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_27_FFY_RST
    );
  rx_input_memio_doutl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(27),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_27_FFX_RST,
      O => rx_input_memio_doutl(27)
    );
  rx_input_memio_doutl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_27_FFX_RST
    );
  rx_input_memio_doutl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(18),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_19_FFY_RST,
      O => rx_input_memio_doutl(18)
    );
  rx_input_memio_doutl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_19_FFY_RST
    );
  rx_input_memio_doutl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(19),
      CE => rx_input_memio_n0033,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_19_FFX_RST,
      O => rx_input_memio_doutl(19)
    );
  rx_input_memio_doutl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_19_FFX_RST
    );
  rx_input_memio_doutl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_dout(28),
      CE => rx_input_memio_n00331_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_doutl_29_FFY_RST,
      O => rx_input_memio_doutl(28)
    );
  rx_input_memio_doutl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_doutl_29_FFY_RST
    );
  rx_input_fifo_control_d2_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(7),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_7_FFX_RST,
      O => rx_input_fifo_control_d2(7)
    );
  rx_input_fifo_control_d2_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_7_FFX_RST
    );
  rx_input_fifo_control_d3_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(2),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_3_FFY_RST,
      O => rx_input_fifo_control_d3(2)
    );
  rx_input_fifo_control_d3_3_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_3_FFY_RST
    );
  rx_input_fifo_control_d3_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(3),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_3_FFX_RST,
      O => rx_input_fifo_control_d3(3)
    );
  rx_input_fifo_control_d3_3_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_3_FFX_RST
    );
  rx_input_fifo_control_d3_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(4),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_5_FFY_RST,
      O => rx_input_fifo_control_d3(4)
    );
  rx_input_fifo_control_d3_5_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_5_FFY_RST
    );
  rx_input_fifo_control_d2_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1(8),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d2_8_FFY_RST,
      O => rx_input_fifo_control_d2(8)
    );
  rx_input_fifo_control_d2_8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d2_8_FFY_RST
    );
  rx_input_fifo_control_d3_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(5),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_5_FFX_RST,
      O => rx_input_fifo_control_d3(5)
    );
  rx_input_fifo_control_d3_5_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_5_FFX_RST
    );
  rx_input_fifo_control_d2_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d1_9_rt,
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_control_d2_9_FFY_SET,
      RST => rx_input_fifo_control_d2_9_FFY_RST,
      O => rx_input_fifo_control_d2(9)
    );
  rx_input_fifo_control_d2_9_FFY_SETOR : X_BUF
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_d2_9_FFY_SET
    );
  rx_input_fifo_control_d2_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_control_d2_9_LOGIC_ZERO,
      I1 => GSR,
      O => rx_input_fifo_control_d2_9_FFY_RST
    );
  rx_input_fifo_control_d3_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(6),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_7_FFY_RST,
      O => rx_input_fifo_control_d3(6)
    );
  rx_input_fifo_control_d3_7_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_7_FFY_RST
    );
  rx_input_fifo_control_d3_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(7),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_7_FFX_RST,
      O => rx_input_fifo_control_d3(7)
    );
  rx_input_fifo_control_d3_7_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_7_FFX_RST
    );
  rx_input_fifo_control_d3_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2_9_rt,
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_fifo_control_d3_9_FFY_SET,
      RST => rx_input_fifo_control_d3_9_FFY_RST,
      O => rx_input_fifo_control_d3(9)
    );
  rx_input_fifo_control_d3_9_FFY_SETOR : X_BUF
    port map (
      I => RESET_IBUF_2,
      O => rx_input_fifo_control_d3_9_FFY_SET
    );
  rx_input_fifo_control_d3_9_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_fifo_control_d3_9_LOGIC_ZERO,
      I1 => GSR,
      O => rx_input_fifo_control_d3_9_FFY_RST
    );
  rx_input_fifo_control_d3_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_d2(8),
      CE => rx_input_fifo_control_celll,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_d3_8_FFY_RST,
      O => rx_input_fifo_control_d3(8)
    );
  rx_input_fifo_control_d3_8_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_2,
      I1 => GSR,
      O => rx_input_fifo_control_d3_8_FFY_RST
    );
  rx_input_memio_crcl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_27_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_27_FFY_RST,
      O => rx_input_memio_crcl(27)
    );
  rx_input_memio_crcl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_27_FFY_RST
    );
  rx_input_memio_crcl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_28_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_28_FFY_RST,
      O => rx_input_memio_crcl(28)
    );
  rx_input_memio_crcl_28_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_28_FFY_RST
    );
  rx_input_memio_crcl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_n0048_29_Q,
      CE => rx_input_memio_n0034,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_crcl_29_FFY_RST,
      O => rx_input_memio_crcl(29)
    );
  rx_input_memio_crcl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_crcl_29_FFY_RST
    );
  rx_input_fifo_control_celll_1894 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_control_cell,
      CE => rx_input_fifo_control_celll_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_celll_FFY_RST,
      O => rx_input_fifo_control_celll
    );
  rx_input_fifo_control_celll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_celll_FFY_RST
    );
  mac_control_rxcrcerr_cntl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(10),
      CE => mac_control_rxcrcerr_cntl_11_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_11_FFY_RST,
      O => mac_control_rxcrcerr_cntl(10)
    );
  mac_control_rxcrcerr_cntl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_11_FFY_RST
    );
  mac_control_rxoferr_cntl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(25),
      CE => mac_control_rxoferr_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_25_FFX_RST,
      O => mac_control_rxoferr_cntl(25)
    );
  mac_control_rxoferr_cntl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_25_FFX_RST
    );
  mac_control_rxoferr_cntl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(16),
      CE => mac_control_rxoferr_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_17_FFY_RST,
      O => mac_control_rxoferr_cntl(16)
    );
  mac_control_rxoferr_cntl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_17_FFY_RST
    );
  mac_control_rxoferr_cntl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(17),
      CE => mac_control_rxoferr_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_17_FFX_RST,
      O => mac_control_rxoferr_cntl(17)
    );
  mac_control_rxoferr_cntl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_17_FFX_RST
    );
  mac_control_rxoferr_cntl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(26),
      CE => mac_control_rxoferr_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_27_FFY_RST,
      O => mac_control_rxoferr_cntl(26)
    );
  mac_control_rxoferr_cntl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_27_FFY_RST
    );
  mac_control_rxoferr_cntl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(27),
      CE => mac_control_rxoferr_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_27_FFX_RST,
      O => mac_control_rxoferr_cntl(27)
    );
  mac_control_rxoferr_cntl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_27_FFX_RST
    );
  mac_control_rxoferr_cntl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(18),
      CE => mac_control_rxoferr_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_19_FFY_RST,
      O => mac_control_rxoferr_cntl(18)
    );
  mac_control_rxoferr_cntl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_19_FFY_RST
    );
  mac_control_rxoferr_cntl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(19),
      CE => mac_control_rxoferr_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_19_FFX_RST,
      O => mac_control_rxoferr_cntl(19)
    );
  mac_control_rxoferr_cntl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_19_FFX_RST
    );
  mac_control_rxoferr_cntl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(28),
      CE => mac_control_rxoferr_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_29_FFY_RST,
      O => mac_control_rxoferr_cntl(28)
    );
  mac_control_rxoferr_cntl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_29_FFY_RST
    );
  mac_control_rxoferr_cntl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxoferr_cnt(29),
      CE => mac_control_rxoferr_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxoferr_cntl_29_FFX_RST,
      O => mac_control_rxoferr_cntl(29)
    );
  mac_control_rxoferr_cntl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxoferr_cntl_29_FFX_RST
    );
  rx_input_GMII_rx_dvll_1895 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_GMII_rx_dvl,
      CE => VCC,
      CLK => clkrx,
      SET => GND,
      RST => rx_input_GMII_rx_dvll_FFY_RST,
      O => rx_input_GMII_rx_dvll
    );
  rx_input_GMII_rx_dvll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_GMII_rx_dvll_FFY_RST
    );
  mac_control_lrxucast_1896 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0027,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lrxucast_FFY_RST,
      O => mac_control_lrxucast
    );
  mac_control_lrxucast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lrxucast_FFY_RST
    );
  rx_input_fifo_control_cell_1897 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_fifo_rd_en,
      CE => rx_input_fifo_control_cell_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_fifo_control_cell_FFY_RST,
      O => rx_input_fifo_control_cell
    );
  rx_input_fifo_control_cell_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_fifo_control_cell_FFY_RST
    );
  tx_input_MA_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_26,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_11_FFY_RST,
      O => addr4ext(10)
    );
  addr4ext_11_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_11_FFY_RST
    );
  tx_input_MA_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_27,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_11_FFX_RST,
      O => addr4ext(11)
    );
  addr4ext_11_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_11_FFX_RST
    );
  tx_input_MA_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_28,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_13_FFY_RST,
      O => addr4ext(12)
    );
  addr4ext_13_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_13_FFY_RST
    );
  tx_input_MA_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_29,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_13_FFX_RST,
      O => addr4ext(13)
    );
  addr4ext_13_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_13_FFX_RST
    );
  tx_input_MA_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_30,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_15_FFY_RST,
      O => addr4ext(14)
    );
  addr4ext_15_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_15_FFY_RST
    );
  tx_input_MA_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_31,
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => addr4ext_15_FFX_RST,
      O => addr4ext(15)
    );
  addr4ext_15_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => addr4ext_15_FFX_RST
    );
  tx_input_MD_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(10),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_11_FFY_RST,
      O => d4(10)
    );
  d4_11_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_11_FFY_RST
    );
  tx_input_MD_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(11),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_11_FFX_RST,
      O => d4(11)
    );
  d4_11_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_11_FFX_RST
    );
  tx_input_MD_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(4),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_21_FFY_RST,
      O => d4(20)
    );
  d4_21_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_21_FFY_RST
    );
  tx_input_MD_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(5),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_21_FFX_RST,
      O => d4(21)
    );
  d4_21_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_21_FFX_RST
    );
  tx_input_MD_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(12),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_13_FFY_RST,
      O => d4(12)
    );
  d4_13_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_13_FFY_RST
    );
  tx_input_MD_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(13),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_13_FFX_RST,
      O => d4(13)
    );
  d4_13_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_13_FFX_RST
    );
  tx_input_MD_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(14),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_15_FFY_RST,
      O => d4(14)
    );
  d4_15_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_15_FFY_RST
    );
  mac_control_rxphyerr_cntl_21 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(21),
      CE => mac_control_rxphyerr_cntl_21_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_21_FFX_RST,
      O => mac_control_rxphyerr_cntl(21)
    );
  mac_control_rxphyerr_cntl_21_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_21_FFX_RST
    );
  mac_control_rxphyerr_cntl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(12),
      CE => mac_control_rxphyerr_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_13_FFY_RST,
      O => mac_control_rxphyerr_cntl(12)
    );
  mac_control_rxphyerr_cntl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_13_FFY_RST
    );
  mac_control_rxphyerr_cntl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(13),
      CE => mac_control_rxphyerr_cntl_13_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_13_FFX_RST,
      O => mac_control_rxphyerr_cntl(13)
    );
  mac_control_rxphyerr_cntl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_13_FFX_RST
    );
  mac_control_rxphyerr_cntl_30 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(30),
      CE => mac_control_rxphyerr_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_31_FFY_RST,
      O => mac_control_rxphyerr_cntl(30)
    );
  mac_control_rxphyerr_cntl_31_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_31_FFY_RST
    );
  mac_control_rxphyerr_cntl_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(31),
      CE => mac_control_rxphyerr_cntl_31_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_31_FFX_RST,
      O => mac_control_rxphyerr_cntl(31)
    );
  mac_control_rxphyerr_cntl_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_31_FFX_RST
    );
  mac_control_rxphyerr_cntl_22 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(22),
      CE => mac_control_rxphyerr_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_23_FFY_RST,
      O => mac_control_rxphyerr_cntl(22)
    );
  mac_control_rxphyerr_cntl_23_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_23_FFY_RST
    );
  mac_control_rxphyerr_cntl_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(23),
      CE => mac_control_rxphyerr_cntl_23_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_23_FFX_RST,
      O => mac_control_rxphyerr_cntl(23)
    );
  mac_control_rxphyerr_cntl_23_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_23_FFX_RST
    );
  mac_control_rxphyerr_cntl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(14),
      CE => mac_control_rxphyerr_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_15_FFY_RST,
      O => mac_control_rxphyerr_cntl(14)
    );
  mac_control_rxphyerr_cntl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_15_FFY_RST
    );
  mac_control_rxphyerr_cntl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(15),
      CE => mac_control_rxphyerr_cntl_15_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_15_FFX_RST,
      O => mac_control_rxphyerr_cntl(15)
    );
  mac_control_rxphyerr_cntl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_15_FFX_RST
    );
  mac_control_rxphyerr_cntl_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(24),
      CE => mac_control_rxphyerr_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_25_FFY_RST,
      O => mac_control_rxphyerr_cntl(24)
    );
  mac_control_rxphyerr_cntl_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_25_FFY_RST
    );
  mac_control_rxphyerr_cntl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(25),
      CE => mac_control_rxphyerr_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_25_FFX_RST,
      O => mac_control_rxphyerr_cntl(25)
    );
  mac_control_rxphyerr_cntl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_25_FFX_RST
    );
  mac_control_rxphyerr_cntl_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(16),
      CE => mac_control_rxphyerr_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_17_FFY_RST,
      O => mac_control_rxphyerr_cntl(16)
    );
  mac_control_rxphyerr_cntl_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_17_FFY_RST
    );
  mac_control_rxphyerr_cntl_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(17),
      CE => mac_control_rxphyerr_cntl_17_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_17_FFX_RST,
      O => mac_control_rxphyerr_cntl(17)
    );
  mac_control_rxphyerr_cntl_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_17_FFX_RST
    );
  mac_control_rxphyerr_cntl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(26),
      CE => mac_control_rxphyerr_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_27_FFY_RST,
      O => mac_control_rxphyerr_cntl(26)
    );
  mac_control_rxphyerr_cntl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_27_FFY_RST
    );
  mac_control_rxcrcerr_cntl_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(25),
      CE => mac_control_rxcrcerr_cntl_25_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_25_FFX_RST,
      O => mac_control_rxcrcerr_cntl(25)
    );
  mac_control_rxcrcerr_cntl_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_25_FFX_RST
    );
  mac_control_rxcrcerr_cntl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(18),
      CE => mac_control_rxcrcerr_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_19_FFY_RST,
      O => mac_control_rxcrcerr_cntl(18)
    );
  mac_control_rxcrcerr_cntl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_19_FFY_RST
    );
  mac_control_rxcrcerr_cntl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(19),
      CE => mac_control_rxcrcerr_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_19_FFX_RST,
      O => mac_control_rxcrcerr_cntl(19)
    );
  mac_control_rxcrcerr_cntl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_19_FFX_RST
    );
  mac_control_rxcrcerr_cntl_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(26),
      CE => mac_control_rxcrcerr_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_27_FFY_RST,
      O => mac_control_rxcrcerr_cntl(26)
    );
  mac_control_rxcrcerr_cntl_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_27_FFY_RST
    );
  mac_control_rxcrcerr_cntl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(27),
      CE => mac_control_rxcrcerr_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_27_FFX_RST,
      O => mac_control_rxcrcerr_cntl(27)
    );
  mac_control_rxcrcerr_cntl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_27_FFX_RST
    );
  mac_control_rxcrcerr_cntl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(28),
      CE => mac_control_rxcrcerr_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_29_FFY_RST,
      O => mac_control_rxcrcerr_cntl(28)
    );
  mac_control_rxcrcerr_cntl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_29_FFY_RST
    );
  mac_control_rxcrcerr_cntl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxcrcerr_cnt(29),
      CE => mac_control_rxcrcerr_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxcrcerr_cntl_29_FFX_RST,
      O => mac_control_rxcrcerr_cntl(29)
    );
  mac_control_rxcrcerr_cntl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxcrcerr_cntl_29_FFX_RST
    );
  rx_input_memio_cs_FFd3_1898 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd3_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd3_FFY_RST,
      O => rx_input_memio_cs_FFd3
    );
  rx_input_memio_cs_FFd3_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd3_FFY_RST
    );
  mac_control_ledrx_rst_1899 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cross,
      CE => mac_control_ledrx_rst_CEMUXNOT,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledrx_rst_FFY_RST,
      O => mac_control_ledrx_rst
    );
  mac_control_ledrx_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledrx_rst_FFY_RST
    );
  rx_input_memio_addrchk_validmcast_1900 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_addrchk_mcast(0),
      CE => rx_input_memio_addrchk_validmcast_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_addrchk_validmcast_FFY_RST,
      O => rx_input_memio_addrchk_validmcast
    );
  rx_input_memio_addrchk_validmcast_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_addrchk_validmcast_FFY_RST
    );
  mac_control_ledtx_rst_1901 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cross,
      CE => mac_control_ledtx_rst_CEMUXNOT,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_ledtx_rst_FFY_RST,
      O => mac_control_ledtx_rst
    );
  mac_control_ledtx_rst_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_ledtx_rst_FFY_RST
    );
  rx_input_memio_cs_FFd4_1902 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd4_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_cs_FFd4_FFY_RST,
      O => rx_input_memio_cs_FFd4
    );
  rx_input_memio_cs_FFd4_FFY_RSTOR : X_OR2
    port map (
      I0 => rx_input_RESET_1,
      I1 => GSR,
      O => rx_input_memio_cs_FFd4_FFY_RST
    );
  tx_input_MD_23 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(7),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_23_FFX_RST,
      O => d4(23)
    );
  d4_23_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_23_FFX_RST
    );
  tx_input_MD_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dl(15),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_15_FFX_RST,
      O => d4(15)
    );
  d4_15_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_15_FFX_RST
    );
  tx_input_MD_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(15),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_31_FFX_RST,
      O => d4(31)
    );
  d4_31_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_31_FFX_RST
    );
  tx_input_MD_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(1),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_17_FFX_RST,
      O => d4(17)
    );
  d4_17_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_17_FFX_RST
    );
  tx_input_MD_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(8),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_25_FFY_RST,
      O => d4(24)
    );
  d4_25_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_25_FFY_RST
    );
  tx_input_MD_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(9),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_25_FFX_RST,
      O => d4(25)
    );
  d4_25_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_25_FFX_RST
    );
  tx_input_MD_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(2),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_19_FFY_RST,
      O => d4(18)
    );
  d4_19_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_19_FFY_RST
    );
  tx_input_MD_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(3),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_19_FFX_RST,
      O => d4(19)
    );
  d4_19_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_19_FFX_RST
    );
  tx_input_MD_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(10),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_27_FFY_RST,
      O => d4(26)
    );
  d4_27_FFY_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_27_FFY_RST
    );
  tx_input_MD_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(11),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_27_FFX_RST,
      O => d4(27)
    );
  d4_27_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_27_FFX_RST
    );
  mac_control_rxf_cntl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxf_cnt(0),
      CE => mac_control_rxf_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_3,
      SET => GND,
      RST => mac_control_rxf_cntl_1_FFY_RST,
      O => mac_control_rxf_cntl(0)
    );
  mac_control_rxf_cntl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxf_cntl_1_FFY_RST
    );
  tx_input_MD_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dh(13),
      CE => tx_input_mrw,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => d4_29_FFX_RST,
      O => d4(29)
    );
  d4_29_FFX_RSTOR : X_OR2
    port map (
      I0 => RESET_IBUF_1,
      I1 => GSR,
      O => d4_29_FFX_RST
    );
  mac_control_txf_cntl_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(7),
      CE => mac_control_txf_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_7_FFX_RST,
      O => mac_control_txf_cntl(7)
    );
  mac_control_txf_cntl_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_7_FFX_RST
    );
  mac_control_txf_cntl_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(8),
      CE => mac_control_txf_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_9_FFY_RST,
      O => mac_control_txf_cntl(8)
    );
  mac_control_txf_cntl_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_9_FFY_RST
    );
  mac_control_txf_cntl_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(9),
      CE => mac_control_txf_cntl_9_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_9_FFX_RST,
      O => mac_control_txf_cntl(9)
    );
  mac_control_txf_cntl_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_9_FFX_RST
    );
  mac_control_addr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_Mshreg_sinlll_102,
      CE => mac_control_n0010,
      CLK => clksl,
      SET => GND,
      RST => mac_control_addr_1_FFY_RST,
      O => mac_control_addr(0)
    );
  mac_control_addr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_1_FFY_RST
    );
  mac_control_addr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr_0_1,
      CE => mac_control_n0010,
      CLK => clksl,
      SET => GND,
      RST => mac_control_addr_1_FFX_RST,
      O => mac_control_addr(1)
    );
  mac_control_addr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_1_FFX_RST
    );
  mac_control_addr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(1),
      CE => mac_control_n0010,
      CLK => clksl,
      SET => GND,
      RST => mac_control_addr_3_FFY_RST,
      O => mac_control_addr(2)
    );
  mac_control_addr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_3_FFY_RST
    );
  mac_control_addr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(2),
      CE => mac_control_n0010,
      CLK => clksl,
      SET => GND,
      RST => mac_control_addr_3_FFX_RST,
      O => mac_control_addr(3)
    );
  mac_control_addr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_3_FFX_RST
    );
  mac_control_addr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(3),
      CE => mac_control_n0010,
      CLK => clksl,
      SET => GND,
      RST => mac_control_addr_5_FFY_RST,
      O => mac_control_addr(4)
    );
  mac_control_addr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_5_FFY_RST
    );
  mac_control_addr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(4),
      CE => mac_control_n0010,
      CLK => clksl,
      SET => GND,
      RST => mac_control_addr_5_FFX_RST,
      O => mac_control_addr(5)
    );
  mac_control_addr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_5_FFX_RST
    );
  mac_control_din_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_11_FFY_RST,
      O => mac_control_din(10)
    );
  mac_control_din_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_11_FFY_RST
    );
  mac_control_addr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(5),
      CE => mac_control_n0010,
      CLK => clksl,
      SET => GND,
      RST => mac_control_addr_7_FFY_RST,
      O => mac_control_addr(6)
    );
  mac_control_addr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_7_FFY_RST
    );
  mac_control_addr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_addr(6),
      CE => mac_control_n0010,
      CLK => clksl,
      SET => GND,
      RST => mac_control_addr_7_FFX_RST,
      O => mac_control_addr(7)
    );
  mac_control_addr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_addr_7_FFX_RST
    );
  mac_control_din_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_11_FFX_RST,
      O => mac_control_din(11)
    );
  mac_control_din_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_11_FFX_RST
    );
  mac_control_din_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_13_FFY_RST,
      O => mac_control_din(12)
    );
  mac_control_din_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_13_FFY_RST
    );
  mac_control_din_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_13_FFX_RST,
      O => mac_control_din(13)
    );
  mac_control_din_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_13_FFX_RST
    );
  mac_control_din_20 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(19),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_21_FFY_RST,
      O => mac_control_din(20)
    );
  mac_control_din_21_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_21_FFY_RST
    );
  mac_control_rxphyerr_cntl_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(27),
      CE => mac_control_rxphyerr_cntl_27_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_27_FFX_RST,
      O => mac_control_rxphyerr_cntl(27)
    );
  mac_control_rxphyerr_cntl_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_27_FFX_RST
    );
  mac_control_rxphyerr_cntl_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(18),
      CE => mac_control_rxphyerr_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_19_FFY_RST,
      O => mac_control_rxphyerr_cntl(18)
    );
  mac_control_rxphyerr_cntl_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_19_FFY_RST
    );
  mac_control_rxphyerr_cntl_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(19),
      CE => mac_control_rxphyerr_cntl_19_CEMUXNOT,
      CLK => mac_control_CLKSL_2,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_19_FFX_RST,
      O => mac_control_rxphyerr_cntl(19)
    );
  mac_control_rxphyerr_cntl_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_19_FFX_RST
    );
  mac_control_rxphyerr_cntl_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(28),
      CE => mac_control_rxphyerr_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_29_FFY_RST,
      O => mac_control_rxphyerr_cntl(28)
    );
  mac_control_rxphyerr_cntl_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_29_FFY_RST
    );
  mac_control_rxphyerr_cntl_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_rxphyerr_cnt(29),
      CE => mac_control_rxphyerr_cntl_29_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_rxphyerr_cntl_29_FFX_RST,
      O => mac_control_rxphyerr_cntl(29)
    );
  mac_control_rxphyerr_cntl_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_rxphyerr_cntl_29_FFX_RST
    );
  tx_fifocheck_bpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(10),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_11_FFY_RST,
      O => tx_fifocheck_bpl(10)
    );
  tx_fifocheck_bpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_11_FFY_RST
    );
  tx_fifocheck_bpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(11),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_11_FFX_RST,
      O => tx_fifocheck_bpl(11)
    );
  tx_fifocheck_bpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_11_FFX_RST
    );
  tx_fifocheck_bpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(12),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_13_FFY_RST,
      O => tx_fifocheck_bpl(12)
    );
  tx_fifocheck_bpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_13_FFY_RST
    );
  tx_fifocheck_bpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(13),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_13_FFX_RST,
      O => tx_fifocheck_bpl(13)
    );
  tx_fifocheck_bpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_13_FFX_RST
    );
  tx_fifocheck_bpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(14),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_15_FFY_RST,
      O => tx_fifocheck_bpl(14)
    );
  tx_fifocheck_bpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_15_FFY_RST
    );
  tx_fifocheck_bpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(15),
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_fifocheck_bpl_15_FFX_RST,
      O => tx_fifocheck_bpl(15)
    );
  tx_fifocheck_bpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_fifocheck_bpl_15_FFX_RST
    );
  mac_control_lmacaddr_19 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_19_FFX_RST,
      O => mac_control_lmacaddr(19)
    );
  mac_control_lmacaddr_19_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_19_FFX_RST
    );
  mac_control_lmacaddr_27 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_27_FFX_RST,
      O => mac_control_lmacaddr(27)
    );
  mac_control_lmacaddr_27_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_27_FFX_RST
    );
  mac_control_lmacaddr_36 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_37_FFY_RST,
      O => mac_control_lmacaddr(36)
    );
  mac_control_lmacaddr_37_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_37_FFY_RST
    );
  mac_control_lmacaddr_37 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_37_FFX_RST,
      O => mac_control_lmacaddr(37)
    );
  mac_control_lmacaddr_37_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_37_FFX_RST
    );
  mac_control_lmacaddr_44 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_45_FFY_RST,
      O => mac_control_lmacaddr(44)
    );
  mac_control_lmacaddr_45_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_45_FFY_RST
    );
  mac_control_lmacaddr_45 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_45_FFX_RST,
      O => mac_control_lmacaddr(45)
    );
  mac_control_lmacaddr_45_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_45_FFX_RST
    );
  mac_control_lmacaddr_28 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(12),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_29_FFY_RST,
      O => mac_control_lmacaddr(28)
    );
  mac_control_lmacaddr_29_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_29_FFY_RST
    );
  mac_control_lmacaddr_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(13),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_29_FFX_RST,
      O => mac_control_lmacaddr(29)
    );
  mac_control_lmacaddr_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_29_FFX_RST
    );
  mac_control_lmacaddr_38 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_39_FFY_RST,
      O => mac_control_lmacaddr(38)
    );
  mac_control_lmacaddr_39_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_39_FFY_RST
    );
  mac_control_lmacaddr_39 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_39_FFX_RST,
      O => mac_control_lmacaddr(39)
    );
  mac_control_lmacaddr_39_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_39_FFX_RST
    );
  mac_control_lmacaddr_46 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_47_FFY_RST,
      O => mac_control_lmacaddr(46)
    );
  mac_control_lmacaddr_47_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_47_FFY_RST
    );
  mac_control_lmacaddr_47 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_47_FFX_RST,
      O => mac_control_lmacaddr(47)
    );
  mac_control_lmacaddr_47_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_47_FFX_RST
    );
  rx_input_memio_BPOUT_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_10_59,
      CE => rxbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_11_FFY_RST,
      O => rxbp(10)
    );
  rxbp_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_11_FFY_RST
    );
  rx_input_memio_BPOUT_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_11_58,
      CE => rxbp_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_11_FFX_RST,
      O => rxbp(11)
    );
  rxbp_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_11_FFX_RST
    );
  rx_input_memio_BPOUT_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_12_57,
      CE => rxbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_13_FFY_RST,
      O => rxbp(12)
    );
  rxbp_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_13_FFY_RST
    );
  rx_input_memio_BPOUT_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_14_55,
      CE => rxbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_15_FFY_RST,
      O => rxbp(14)
    );
  rxbp_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_15_FFY_RST
    );
  mac_control_lmacaddr_31 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_31_FFX_RST,
      O => mac_control_lmacaddr(31)
    );
  mac_control_lmacaddr_31_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_31_FFX_RST
    );
  mac_control_lmacaddr_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(14),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_15_FFY_RST,
      O => mac_control_lmacaddr(14)
    );
  mac_control_lmacaddr_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_15_FFY_RST
    );
  mac_control_lmacaddr_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(15),
      CE => mac_control_n0028,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_15_FFX_RST,
      O => mac_control_lmacaddr(15)
    );
  mac_control_lmacaddr_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_15_FFX_RST
    );
  mac_control_lmacaddr_40 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_41_FFY_RST,
      O => mac_control_lmacaddr(40)
    );
  mac_control_lmacaddr_41_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_41_FFY_RST
    );
  mac_control_lmacaddr_32 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_33_FFY_RST,
      O => mac_control_lmacaddr(32)
    );
  mac_control_lmacaddr_33_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_33_FFY_RST
    );
  mac_control_lmacaddr_33 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_33_FFX_RST,
      O => mac_control_lmacaddr(33)
    );
  mac_control_lmacaddr_33_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_33_FFX_RST
    );
  mac_control_lmacaddr_41 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_41_FFX_RST,
      O => mac_control_lmacaddr(41)
    );
  mac_control_lmacaddr_41_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_41_FFX_RST
    );
  mac_control_lmacaddr_16 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_17_FFY_RST,
      O => mac_control_lmacaddr(16)
    );
  mac_control_lmacaddr_17_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_17_FFY_RST
    );
  mac_control_lmacaddr_17 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_17_FFX_RST,
      O => mac_control_lmacaddr(17)
    );
  mac_control_lmacaddr_17_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_17_FFX_RST
    );
  mac_control_lmacaddr_24 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(8),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_25_FFY_RST,
      O => mac_control_lmacaddr(24)
    );
  mac_control_lmacaddr_25_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_25_FFY_RST
    );
  mac_control_lmacaddr_25 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(9),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_25_FFX_RST,
      O => mac_control_lmacaddr(25)
    );
  mac_control_lmacaddr_25_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_25_FFX_RST
    );
  mac_control_lmacaddr_34 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_35_FFY_RST,
      O => mac_control_lmacaddr(34)
    );
  mac_control_lmacaddr_35_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_35_FFY_RST
    );
  mac_control_lmacaddr_35 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_35_FFX_RST,
      O => mac_control_lmacaddr(35)
    );
  mac_control_lmacaddr_35_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_35_FFX_RST
    );
  mac_control_lmacaddr_42 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_43_FFY_RST,
      O => mac_control_lmacaddr(42)
    );
  mac_control_lmacaddr_43_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_43_FFY_RST
    );
  mac_control_lmacaddr_43 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(11),
      CE => mac_control_n0030,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_43_FFX_RST,
      O => mac_control_lmacaddr(43)
    );
  mac_control_lmacaddr_43_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_43_FFX_RST
    );
  mac_control_lmacaddr_18 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_19_FFY_RST,
      O => mac_control_lmacaddr(18)
    );
  mac_control_lmacaddr_19_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_19_FFY_RST
    );
  mac_control_lmacaddr_26 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(10),
      CE => mac_control_n0029,
      CLK => mac_control_CLKSL_5,
      SET => GND,
      RST => mac_control_lmacaddr_27_FFY_RST,
      O => mac_control_lmacaddr(26)
    );
  mac_control_lmacaddr_27_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_lmacaddr_27_FFY_RST
    );
  tx_input_dh_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(10),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_11_FFY_RST,
      O => tx_input_dh(10)
    );
  tx_input_dh_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_11_FFY_RST
    );
  tx_input_dh_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(11),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_11_FFX_RST,
      O => tx_input_dh(11)
    );
  tx_input_dh_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_11_FFX_RST
    );
  tx_input_dh_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(12),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_13_FFY_RST,
      O => tx_input_dh(12)
    );
  tx_input_dh_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_13_FFY_RST
    );
  tx_input_dh_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(13),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_13_FFX_RST,
      O => tx_input_dh(13)
    );
  tx_input_dh_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_13_FFX_RST
    );
  tx_input_dh_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(14),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_15_FFY_RST,
      O => tx_input_dh(14)
    );
  tx_input_dh_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_15_FFY_RST
    );
  tx_input_dh_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(15),
      CE => tx_input_n0021,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dh_15_FFX_RST,
      O => tx_input_dh(15)
    );
  tx_input_dh_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dh_15_FFX_RST
    );
  tx_input_dl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(10),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_11_FFY_RST,
      O => tx_input_dl(10)
    );
  tx_input_dl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_11_FFY_RST
    );
  tx_input_dl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(11),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_11_FFX_RST,
      O => tx_input_dl(11)
    );
  tx_input_dl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_11_FFX_RST
    );
  tx_input_bp_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_26,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_11_FFY_RST,
      O => txbp(10)
    );
  txbp_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_11_FFY_RST
    );
  tx_input_bp_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_27,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_11_FFX_RST,
      O => txbp(11)
    );
  txbp_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_11_FFX_RST
    );
  tx_input_dl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(12),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_13_FFY_RST,
      O => tx_input_dl(12)
    );
  tx_input_dl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_13_FFY_RST
    );
  tx_input_dl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(13),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_13_FFX_RST,
      O => tx_input_dl(13)
    );
  tx_input_dl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_13_FFX_RST
    );
  tx_input_bp_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_28,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_13_FFY_RST,
      O => txbp(12)
    );
  txbp_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_13_FFY_RST
    );
  tx_input_dl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_dinint(14),
      CE => tx_input_n0020,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_input_dl_15_FFY_RST,
      O => tx_input_dl(14)
    );
  tx_input_dl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_input_dl_15_FFY_RST
    );
  tx_input_bp_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_input_addr_29,
      CE => tx_input_n0023,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => txbp_13_FFX_RST,
      O => txbp(13)
    );
  txbp_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => txbp_13_FFX_RST
    );
  tx_output_outsell_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_cs_FFd9,
      CE => tx_output_outsell_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outsell_2_FFX_RST,
      O => tx_output_outsell(2)
    );
  tx_output_outsell_2_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outsell_2_FFX_RST
    );
  rx_input_memio_fifofulll_1903 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rxfifofull,
      CE => rx_input_memio_fifofulll_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_fifofulll_FFY_RST,
      O => rx_input_memio_fifofulll
    );
  rx_input_memio_fifofulll_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_fifofulll_FFY_RST
    );
  rx_input_memio_endbyte_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(0),
      CE => rx_input_memio_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_endbyte_1_FFY_RST,
      O => rx_input_memio_endbyte(0)
    );
  rx_input_memio_endbyte_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_endbyte_1_FFY_RST
    );
  rx_input_memio_endbyte_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(2),
      CE => rx_input_memio_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_endbyte_2_FFY_RST,
      O => rx_input_memio_endbyte(2)
    );
  rx_input_memio_endbyte_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_endbyte_2_FFY_RST
    );
  rx_input_memio_endbyte_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_data(1),
      CE => rx_input_memio_n0032,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_endbyte_1_FFX_RST,
      O => rx_input_memio_endbyte(1)
    );
  rx_input_memio_endbyte_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_endbyte_1_FFX_RST
    );
  rx_output_nfl_1904 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_output_nf,
      CE => rx_output_nfl_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_output_nfl_FFY_RST,
      O => rx_output_nfl
    );
  rx_output_nfl_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_output_nfl_FFY_RST
    );
  mac_control_txf_cntl_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(0),
      CE => mac_control_txf_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_1_FFY_RST,
      O => mac_control_txf_cntl(0)
    );
  mac_control_txf_cntl_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_1_FFY_RST
    );
  mac_control_txf_cntl_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(1),
      CE => mac_control_txf_cntl_1_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_1_FFX_RST,
      O => mac_control_txf_cntl(1)
    );
  mac_control_txf_cntl_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_1_FFX_RST
    );
  mac_control_txf_cntl_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(2),
      CE => mac_control_txf_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_3_FFY_RST,
      O => mac_control_txf_cntl(2)
    );
  mac_control_txf_cntl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_3_FFY_RST
    );
  mac_control_txf_cntl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(3),
      CE => mac_control_txf_cntl_3_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_3_FFX_RST,
      O => mac_control_txf_cntl(3)
    );
  mac_control_txf_cntl_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_3_FFX_RST
    );
  mac_control_txf_cntl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(4),
      CE => mac_control_txf_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_5_FFY_RST,
      O => mac_control_txf_cntl(4)
    );
  mac_control_txf_cntl_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_5_FFY_RST
    );
  mac_control_txf_cntl_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(5),
      CE => mac_control_txf_cntl_5_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_5_FFX_RST,
      O => mac_control_txf_cntl(5)
    );
  mac_control_txf_cntl_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_5_FFX_RST
    );
  mac_control_txf_cntl_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_txf_cnt(6),
      CE => mac_control_txf_cntl_7_CEMUXNOT,
      CLK => mac_control_CLKSL_1,
      SET => GND,
      RST => mac_control_txf_cntl_7_FFY_RST,
      O => mac_control_txf_cntl(6)
    );
  mac_control_txf_cntl_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_txf_cntl_7_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(9),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_9_FFX_RST,
      O => mac_control_PHY_status_dout(9)
    );
  mac_control_PHY_status_dout_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_9_FFX_RST
    );
  rx_input_memio_bpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(10),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_11_FFY_RST,
      O => rx_input_memio_bpl(10)
    );
  rx_input_memio_bpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_11_FFY_RST
    );
  rx_input_memio_bpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(11),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_11_FFX_RST,
      O => rx_input_memio_bpl(11)
    );
  rx_input_memio_bpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_11_FFX_RST
    );
  rx_input_memio_bpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(12),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_13_FFY_RST,
      O => rx_input_memio_bpl(12)
    );
  rx_input_memio_bpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_13_FFY_RST
    );
  rx_input_memio_bpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(13),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_13_FFX_RST,
      O => rx_input_memio_bpl(13)
    );
  rx_input_memio_bpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_13_FFX_RST
    );
  rx_input_memio_bpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(14),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_15_FFY_RST,
      O => rx_input_memio_bpl(14)
    );
  rx_input_memio_bpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_15_FFY_RST
    );
  rx_input_memio_bpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_bp(15),
      CE => rx_input_memio_n0030,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rx_input_memio_bpl_15_FFX_RST,
      O => rx_input_memio_bpl(15)
    );
  rx_input_memio_bpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rx_input_memio_bpl_15_FFX_RST
    );
  rx_input_memio_RXF : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_cs_FFd1,
      CE => rxf_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxf_FFY_RST,
      O => rxf
    );
  rxf_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxf_FFY_RST
    );
  tx_output_crcl_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_4_1_O,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_4_FFY_RST,
      O => tx_output_crcl(4)
    );
  tx_output_crcl_4_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_4_FFY_RST
    );
  mac_control_phyaddr_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(1),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_1_FFX_RST,
      O => mac_control_phyaddr(1)
    );
  mac_control_phyaddr_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_1_FFX_RST
    );
  mac_control_phyaddr_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(0),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_1_FFY_RST,
      O => mac_control_phyaddr(0)
    );
  mac_control_phyaddr_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_1_FFY_RST
    );
  mac_control_phyaddr_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(2),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_3_FFY_RST,
      O => mac_control_phyaddr(2)
    );
  mac_control_phyaddr_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_3_FFY_RST
    );
  mac_control_phyaddr_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(4),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_5_FFY_RST,
      O => mac_control_phyaddr(4)
    );
  mac_control_phyaddr_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_5_FFY_RST
    );
  rx_input_memio_BPOUT_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_13_56,
      CE => rxbp_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_13_FFX_RST,
      O => rxbp(13)
    );
  rxbp_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_13_FFX_RST
    );
  rx_input_memio_BPOUT_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => rx_input_memio_Mshreg_lbpout4_15_54,
      CE => rxbp_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => rxbp_15_FFX_RST,
      O => rxbp(15)
    );
  rxbp_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => rxbp_15_FFX_RST
    );
  memcontroller_Q2_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(0),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_1_FFY_RST,
      O => q2(0)
    );
  q2_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_1_FFY_RST
    );
  memcontroller_Q2_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(1),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_1_FFX_RST,
      O => q2(1)
    );
  q2_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_1_FFX_RST
    );
  memcontroller_Q2_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(2),
      CE => memcontroller_n0005,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_2_FFY_RST,
      O => q2(2)
    );
  q2_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_2_FFY_RST
    );
  memcontroller_Q2_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(3),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_3_FFY_RST,
      O => q2(3)
    );
  q2_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_3_FFY_RST
    );
  memcontroller_Q2_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(4),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_5_FFY_RST,
      O => q2(4)
    );
  q2_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_5_FFY_RST
    );
  memcontroller_Q2_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(5),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_5_FFX_RST,
      O => q2(5)
    );
  q2_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_5_FFX_RST
    );
  memcontroller_Q3_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(0),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_1_FFY_RST,
      O => q3(0)
    );
  q3_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_1_FFY_RST
    );
  memcontroller_Q3_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(1),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_1_FFX_RST,
      O => q3(1)
    );
  q3_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_1_FFX_RST
    );
  memcontroller_Q2_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(6),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_7_FFY_RST,
      O => q2(6)
    );
  q2_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_7_FFY_RST
    );
  memcontroller_Q2_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(7),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_7_FFX_RST,
      O => q2(7)
    );
  q2_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_7_FFX_RST
    );
  memcontroller_Q3_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(2),
      CE => memcontroller_n0006,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_2_FFY_RST,
      O => q3(2)
    );
  q3_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_2_FFY_RST
    );
  memcontroller_Q3_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(3),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_3_FFY_RST,
      O => q3(3)
    );
  q3_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_3_FFY_RST
    );
  memcontroller_Q2_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(8),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_9_FFY_RST,
      O => q2(8)
    );
  q2_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_9_FFY_RST
    );
  memcontroller_Q2_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(9),
      CE => memcontroller_n00051_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q2_9_FFX_RST,
      O => q2(9)
    );
  q2_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q2_9_FFX_RST
    );
  memcontroller_Q3_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(4),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_5_FFY_RST,
      O => q3(4)
    );
  q3_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_5_FFY_RST
    );
  memcontroller_Q3_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(5),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_5_FFX_RST,
      O => q3(5)
    );
  q3_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_5_FFX_RST
    );
  memcontroller_Q3_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(6),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_7_FFY_RST,
      O => q3(6)
    );
  q3_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_7_FFY_RST
    );
  memcontroller_Q3_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(7),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_7_FFX_RST,
      O => q3(7)
    );
  q3_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_7_FFX_RST
    );
  memcontroller_Q3_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(8),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_9_FFY_RST,
      O => q3(8)
    );
  q3_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_9_FFY_RST
    );
  memcontroller_Q3_9 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => memcontroller_qn(9),
      CE => memcontroller_n00061_1,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => q3_9_FFX_RST,
      O => q3(9)
    );
  q3_9_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => q3_9_FFX_RST
    );
  tx_output_bpl_10 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(10),
      CE => tx_output_bpl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_11_FFY_RST,
      O => tx_output_bpl(10)
    );
  tx_output_bpl_11_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_11_FFY_RST
    );
  tx_output_bpl_11 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(11),
      CE => tx_output_bpl_11_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_11_FFX_RST,
      O => tx_output_bpl(11)
    );
  tx_output_bpl_11_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_11_FFX_RST
    );
  tx_output_bpl_12 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(12),
      CE => tx_output_bpl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_13_FFY_RST,
      O => tx_output_bpl(12)
    );
  tx_output_bpl_13_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_13_FFY_RST
    );
  tx_output_bpl_13 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(13),
      CE => tx_output_bpl_13_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_13_FFX_RST,
      O => tx_output_bpl(13)
    );
  tx_output_bpl_13_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_13_FFX_RST
    );
  tx_output_bpl_14 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(14),
      CE => tx_output_bpl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_15_FFY_RST,
      O => tx_output_bpl(14)
    );
  tx_output_bpl_15_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_15_FFY_RST
    );
  tx_output_bpl_15 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => txbp(15),
      CE => tx_output_bpl_15_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_bpl_15_FFX_RST,
      O => tx_output_bpl(15)
    );
  tx_output_bpl_15_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_bpl_15_FFX_RST
    );
  tx_output_outsell_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_outsel_3_Q,
      CE => tx_output_outsell_2_CEMUXNOT,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_outsell_2_FFY_RST,
      O => tx_output_outsell(3)
    );
  tx_output_outsell_2_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_outsell_2_FFY_RST
    );
  mac_control_phyaddr_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(3),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_3_FFX_RST,
      O => mac_control_phyaddr(3)
    );
  mac_control_phyaddr_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_3_FFX_RST
    );
  mac_control_phyaddr_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(5),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_5_FFX_RST,
      O => mac_control_phyaddr(5)
    );
  mac_control_phyaddr_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_5_FFX_RST
    );
  mac_control_phyaddr_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(6),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_7_FFY_RST,
      O => mac_control_phyaddr(6)
    );
  mac_control_phyaddr_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_7_FFY_RST
    );
  mac_control_phyaddr_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(7),
      CE => mac_control_n0024,
      CLK => mac_control_CLKSL_4,
      SET => GND,
      RST => mac_control_phyaddr_7_FFX_RST,
      O => mac_control_phyaddr(7)
    );
  mac_control_phyaddr_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_phyaddr_7_FFX_RST
    );
  mac_control_din_29 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_din(28),
      CE => mac_control_n0011,
      CLK => clksl,
      SET => GND,
      RST => mac_control_din_29_FFX_RST,
      O => mac_control_din(29)
    );
  mac_control_din_29_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_din_29_FFX_RST
    );
  memcontroller_ts_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => memcontroller_oel,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => memcontroller_ts_0_FFY_SET,
      RST => GND,
      O => memcontroller_ts(0)
    );
  memcontroller_ts_0_FFY_SETOR : X_BUF
    port map (
      I => GSR,
      O => memcontroller_ts_0_FFY_SET
    );
  tx_output_crcl_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => tx_output_n0034_3_Q,
      CE => tx_output_n0025,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => tx_output_crcl_3_FFY_RST,
      O => tx_output_crcl(3)
    );
  tx_output_crcl_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => tx_output_crcl_3_FFY_RST
    );
  rx_input_memio_cs_FFd16_2_1905 : X_FF
    generic map(
      XON => FALSE,
      INIT => '1'
    )
    port map (
      I => rx_input_memio_cs_FFd16_In,
      CE => VCC,
      CLK => GTX_CLK_OBUF,
      SET => rx_input_memio_cs_FFd16_2_FFY_SET,
      RST => GND,
      O => rx_input_memio_cs_FFd16_2
    );
  rx_input_memio_cs_FFd16_2_FFY_SETOR : X_OR2
    port map (
      I0 => GSR,
      I1 => rx_input_RESET_1,
      O => rx_input_memio_cs_FFd16_2_FFY_SET
    );
  mac_control_PHY_status_MII_Interface_DOUT_1 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(1),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_1_FFX_RST,
      O => mac_control_PHY_status_dout(1)
    );
  mac_control_PHY_status_dout_1_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_1_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_0 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(0),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_1_FFY_RST,
      O => mac_control_PHY_status_dout(0)
    );
  mac_control_PHY_status_dout_1_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_1_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_2 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(2),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_3_FFY_RST,
      O => mac_control_PHY_status_dout(2)
    );
  mac_control_PHY_status_dout_3_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_3_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_3 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(3),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_3_FFX_RST,
      O => mac_control_PHY_status_dout(3)
    );
  mac_control_PHY_status_dout_3_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_3_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_4 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(4),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_5_FFY_RST,
      O => mac_control_PHY_status_dout(4)
    );
  mac_control_PHY_status_dout_5_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_5_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_5 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(5),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_5_FFX_RST,
      O => mac_control_PHY_status_dout(5)
    );
  mac_control_PHY_status_dout_5_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_5_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_6 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(6),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_7_FFY_RST,
      O => mac_control_PHY_status_dout(6)
    );
  mac_control_PHY_status_dout_7_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_7_FFY_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_7 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(7),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_7_FFX_RST,
      O => mac_control_PHY_status_dout(7)
    );
  mac_control_PHY_status_dout_7_FFX_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_7_FFX_RST
    );
  mac_control_PHY_status_MII_Interface_DOUT_8 : X_FF
    generic map(
      XON => FALSE,
      INIT => '0'
    )
    port map (
      I => mac_control_PHY_status_MII_Interface_dreg(8),
      CE => mac_control_PHY_status_MII_Interface_n0015,
      CLK => GTX_CLK_OBUF,
      SET => GND,
      RST => mac_control_PHY_status_dout_9_FFY_RST,
      O => mac_control_PHY_status_dout(8)
    );
  mac_control_PHY_status_dout_9_FFY_RSTOR : X_BUF
    port map (
      I => GSR,
      O => mac_control_PHY_status_dout_9_FFY_RST
    );
  CLKIN_BUF : X_CKBUF
    port map (
      I => CLKIN,
      O => CLKIN_IBUFG
    );
  RX_CLK_BUF : X_CKBUF
    port map (
      I => RX_CLK,
      O => RX_CLK_IBUFG
    );
  CLKIOIN_BUF : X_CKBUF
    port map (
      I => CLKIOIN,
      O => CLKIOIN_IBUFG
    );
  clkio_bufg_BUF : X_CKBUF
    port map (
      I => clkio_to_bufg,
      O => clkio
    );
  clk_bufg_BUF : X_CKBUF
    port map (
      I => clk_to_bufg,
      O => GTX_CLK_OBUF
    );
  clkrx_bufg_BUF : X_CKBUF
    port map (
      I => clkrx_to_bufg,
      O => clkrx
    );
  PWR_GND_0_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_0_GROM
    );
  PWR_GND_0_YUSED : X_BUF
    port map (
      I => PWR_GND_0_GROM,
      O => GLOBAL_LOGIC0
    );
  PWR_GND_1_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_1_GROM
    );
  PWR_GND_1_YUSED : X_BUF
    port map (
      I => PWR_GND_1_GROM,
      O => GLOBAL_LOGIC0_0
    );
  PWR_GND_2_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_2_GROM
    );
  PWR_GND_2_YUSED : X_BUF
    port map (
      I => PWR_GND_2_GROM,
      O => GLOBAL_LOGIC0_1
    );
  PWR_GND_3_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_3_GROM
    );
  PWR_GND_3_YUSED : X_BUF
    port map (
      I => PWR_GND_3_GROM,
      O => GLOBAL_LOGIC0_2
    );
  PWR_GND_4_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_4_GROM
    );
  PWR_GND_4_YUSED : X_BUF
    port map (
      I => PWR_GND_4_GROM,
      O => GLOBAL_LOGIC0_3
    );
  PWR_GND_5_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_5_GROM
    );
  PWR_GND_5_YUSED : X_BUF
    port map (
      I => PWR_GND_5_GROM,
      O => GLOBAL_LOGIC0_4
    );
  PWR_GND_6_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_6_GROM
    );
  PWR_GND_6_YUSED : X_BUF
    port map (
      I => PWR_GND_6_GROM,
      O => GLOBAL_LOGIC0_5
    );
  PWR_GND_7_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_7_GROM
    );
  PWR_GND_7_YUSED : X_BUF
    port map (
      I => PWR_GND_7_GROM,
      O => GLOBAL_LOGIC0_6
    );
  PWR_GND_8_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_8_GROM
    );
  PWR_GND_8_YUSED : X_BUF
    port map (
      I => PWR_GND_8_GROM,
      O => GLOBAL_LOGIC0_7
    );
  PWR_GND_9_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_9_FROM
    );
  PWR_GND_9_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_9_GROM
    );
  PWR_GND_9_XUSED : X_BUF
    port map (
      I => PWR_GND_9_FROM,
      O => GLOBAL_LOGIC1
    );
  PWR_GND_9_YUSED : X_BUF
    port map (
      I => PWR_GND_9_GROM,
      O => GLOBAL_LOGIC0_8
    );
  PWR_GND_10_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_10_FROM
    );
  PWR_GND_10_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_10_GROM
    );
  PWR_GND_10_XUSED : X_BUF
    port map (
      I => PWR_GND_10_FROM,
      O => GLOBAL_LOGIC1_0
    );
  PWR_GND_10_YUSED : X_BUF
    port map (
      I => PWR_GND_10_GROM,
      O => GLOBAL_LOGIC0_9
    );
  PWR_GND_11_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_11_FROM
    );
  PWR_GND_11_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_11_GROM
    );
  PWR_GND_11_XUSED : X_BUF
    port map (
      I => PWR_GND_11_FROM,
      O => GLOBAL_LOGIC1_1
    );
  PWR_GND_11_YUSED : X_BUF
    port map (
      I => PWR_GND_11_GROM,
      O => GLOBAL_LOGIC0_10
    );
  PWR_GND_12_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_12_FROM
    );
  PWR_GND_12_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_12_GROM
    );
  PWR_GND_12_XUSED : X_BUF
    port map (
      I => PWR_GND_12_FROM,
      O => GLOBAL_LOGIC1_2
    );
  PWR_GND_12_YUSED : X_BUF
    port map (
      I => PWR_GND_12_GROM,
      O => GLOBAL_LOGIC0_11
    );
  PWR_GND_13_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_13_FROM
    );
  PWR_GND_13_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_13_GROM
    );
  PWR_GND_13_XUSED : X_BUF
    port map (
      I => PWR_GND_13_FROM,
      O => GLOBAL_LOGIC1_3
    );
  PWR_GND_13_YUSED : X_BUF
    port map (
      I => PWR_GND_13_GROM,
      O => GLOBAL_LOGIC0_12
    );
  PWR_GND_14_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_14_FROM
    );
  PWR_GND_14_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_14_GROM
    );
  PWR_GND_14_XUSED : X_BUF
    port map (
      I => PWR_GND_14_FROM,
      O => GLOBAL_LOGIC1_4
    );
  PWR_GND_14_YUSED : X_BUF
    port map (
      I => PWR_GND_14_GROM,
      O => GLOBAL_LOGIC0_13
    );
  PWR_GND_15_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_15_GROM
    );
  PWR_GND_15_YUSED : X_BUF
    port map (
      I => PWR_GND_15_GROM,
      O => GLOBAL_LOGIC0_14
    );
  PWR_GND_16_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_16_GROM
    );
  PWR_GND_16_YUSED : X_BUF
    port map (
      I => PWR_GND_16_GROM,
      O => GLOBAL_LOGIC0_15
    );
  PWR_GND_17_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_17_FROM
    );
  PWR_GND_17_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_17_GROM
    );
  PWR_GND_17_XUSED : X_BUF
    port map (
      I => PWR_GND_17_FROM,
      O => GLOBAL_LOGIC1_9
    );
  PWR_GND_17_YUSED : X_BUF
    port map (
      I => PWR_GND_17_GROM,
      O => GLOBAL_LOGIC0_16
    );
  PWR_GND_18_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_18_GROM
    );
  PWR_GND_18_YUSED : X_BUF
    port map (
      I => PWR_GND_18_GROM,
      O => GLOBAL_LOGIC0_17
    );
  PWR_GND_19_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_19_FROM
    );
  PWR_GND_19_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_19_GROM
    );
  PWR_GND_19_XUSED : X_BUF
    port map (
      I => PWR_GND_19_FROM,
      O => GLOBAL_LOGIC1_11
    );
  PWR_GND_19_YUSED : X_BUF
    port map (
      I => PWR_GND_19_GROM,
      O => GLOBAL_LOGIC0_18
    );
  PWR_GND_20_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_20_GROM
    );
  PWR_GND_20_YUSED : X_BUF
    port map (
      I => PWR_GND_20_GROM,
      O => GLOBAL_LOGIC0_19
    );
  PWR_GND_21_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_21_GROM
    );
  PWR_GND_21_YUSED : X_BUF
    port map (
      I => PWR_GND_21_GROM,
      O => GLOBAL_LOGIC0_20
    );
  PWR_GND_22_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_22_GROM
    );
  PWR_GND_22_YUSED : X_BUF
    port map (
      I => PWR_GND_22_GROM,
      O => GLOBAL_LOGIC0_21
    );
  PWR_GND_23_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_23_FROM
    );
  PWR_GND_23_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_23_GROM
    );
  PWR_GND_23_XUSED : X_BUF
    port map (
      I => PWR_GND_23_FROM,
      O => GLOBAL_LOGIC1_14
    );
  PWR_GND_23_YUSED : X_BUF
    port map (
      I => PWR_GND_23_GROM,
      O => GLOBAL_LOGIC0_22
    );
  PWR_GND_24_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_24_GROM
    );
  PWR_GND_24_YUSED : X_BUF
    port map (
      I => PWR_GND_24_GROM,
      O => GLOBAL_LOGIC0_23
    );
  PWR_GND_25_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_25_FROM
    );
  PWR_GND_25_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_25_GROM
    );
  PWR_GND_25_XUSED : X_BUF
    port map (
      I => PWR_GND_25_FROM,
      O => GLOBAL_LOGIC1_16
    );
  PWR_GND_25_YUSED : X_BUF
    port map (
      I => PWR_GND_25_GROM,
      O => GLOBAL_LOGIC0_24
    );
  PWR_GND_26_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_26_GROM
    );
  PWR_GND_26_YUSED : X_BUF
    port map (
      I => PWR_GND_26_GROM,
      O => GLOBAL_LOGIC0_25
    );
  PWR_GND_27_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_27_GROM
    );
  PWR_GND_27_YUSED : X_BUF
    port map (
      I => PWR_GND_27_GROM,
      O => GLOBAL_LOGIC0_26
    );
  PWR_GND_28_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_28_GROM
    );
  PWR_GND_28_YUSED : X_BUF
    port map (
      I => PWR_GND_28_GROM,
      O => GLOBAL_LOGIC0_27
    );
  PWR_GND_29_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_29_FROM
    );
  PWR_GND_29_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_29_GROM
    );
  PWR_GND_29_XUSED : X_BUF
    port map (
      I => PWR_GND_29_FROM,
      O => GLOBAL_LOGIC1_19
    );
  PWR_GND_29_YUSED : X_BUF
    port map (
      I => PWR_GND_29_GROM,
      O => GLOBAL_LOGIC0_28
    );
  PWR_GND_30_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_30_FROM
    );
  PWR_GND_30_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_30_GROM
    );
  PWR_GND_30_XUSED : X_BUF
    port map (
      I => PWR_GND_30_FROM,
      O => GLOBAL_LOGIC1_20
    );
  PWR_GND_30_YUSED : X_BUF
    port map (
      I => PWR_GND_30_GROM,
      O => GLOBAL_LOGIC0_29
    );
  PWR_GND_31_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_31_GROM
    );
  PWR_GND_31_YUSED : X_BUF
    port map (
      I => PWR_GND_31_GROM,
      O => GLOBAL_LOGIC0_30
    );
  PWR_GND_32_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_32_GROM
    );
  PWR_GND_32_YUSED : X_BUF
    port map (
      I => PWR_GND_32_GROM,
      O => GLOBAL_LOGIC0_31
    );
  PWR_GND_33_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_33_GROM
    );
  PWR_GND_33_YUSED : X_BUF
    port map (
      I => PWR_GND_33_GROM,
      O => GLOBAL_LOGIC0_32
    );
  PWR_GND_34_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_34_GROM
    );
  PWR_GND_34_YUSED : X_BUF
    port map (
      I => PWR_GND_34_GROM,
      O => GLOBAL_LOGIC0_33
    );
  PWR_GND_35_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_35_FROM
    );
  PWR_GND_35_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_35_GROM
    );
  PWR_GND_35_XUSED : X_BUF
    port map (
      I => PWR_GND_35_FROM,
      O => GLOBAL_LOGIC1_21
    );
  PWR_GND_35_YUSED : X_BUF
    port map (
      I => PWR_GND_35_GROM,
      O => GLOBAL_LOGIC0_34
    );
  PWR_GND_36_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_36_FROM
    );
  PWR_GND_36_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_36_GROM
    );
  PWR_GND_36_XUSED : X_BUF
    port map (
      I => PWR_GND_36_FROM,
      O => GLOBAL_LOGIC1_22
    );
  PWR_GND_36_YUSED : X_BUF
    port map (
      I => PWR_GND_36_GROM,
      O => GLOBAL_LOGIC0_35
    );
  PWR_GND_37_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_37_FROM
    );
  PWR_GND_37_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_37_GROM
    );
  PWR_GND_37_XUSED : X_BUF
    port map (
      I => PWR_GND_37_FROM,
      O => GLOBAL_LOGIC1_23
    );
  PWR_GND_37_YUSED : X_BUF
    port map (
      I => PWR_GND_37_GROM,
      O => GLOBAL_LOGIC0_36
    );
  PWR_GND_38_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_38_FROM
    );
  PWR_GND_38_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_38_GROM
    );
  PWR_GND_38_XUSED : X_BUF
    port map (
      I => PWR_GND_38_FROM,
      O => GLOBAL_LOGIC1_24
    );
  PWR_GND_38_YUSED : X_BUF
    port map (
      I => PWR_GND_38_GROM,
      O => GLOBAL_LOGIC0_37
    );
  PWR_GND_39_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_39_GROM
    );
  PWR_GND_39_YUSED : X_BUF
    port map (
      I => PWR_GND_39_GROM,
      O => GLOBAL_LOGIC0_38
    );
  PWR_GND_40_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_40_FROM
    );
  PWR_GND_40_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_40_GROM
    );
  PWR_GND_40_XUSED : X_BUF
    port map (
      I => PWR_GND_40_FROM,
      O => GLOBAL_LOGIC1_25
    );
  PWR_GND_40_YUSED : X_BUF
    port map (
      I => PWR_GND_40_GROM,
      O => GLOBAL_LOGIC0_39
    );
  PWR_GND_41_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_41_GROM
    );
  PWR_GND_41_YUSED : X_BUF
    port map (
      I => PWR_GND_41_GROM,
      O => GLOBAL_LOGIC0_40
    );
  PWR_GND_42_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_42_FROM
    );
  PWR_GND_42_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_42_GROM
    );
  PWR_GND_42_XUSED : X_BUF
    port map (
      I => PWR_GND_42_FROM,
      O => GLOBAL_LOGIC1_26
    );
  PWR_GND_42_YUSED : X_BUF
    port map (
      I => PWR_GND_42_GROM,
      O => GLOBAL_LOGIC0_41
    );
  PWR_GND_43_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_43_GROM
    );
  PWR_GND_43_YUSED : X_BUF
    port map (
      I => PWR_GND_43_GROM,
      O => GLOBAL_LOGIC0_42
    );
  PWR_GND_44_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_44_FROM
    );
  PWR_GND_44_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_44_GROM
    );
  PWR_GND_44_XUSED : X_BUF
    port map (
      I => PWR_GND_44_FROM,
      O => GLOBAL_LOGIC1_29
    );
  PWR_GND_44_YUSED : X_BUF
    port map (
      I => PWR_GND_44_GROM,
      O => GLOBAL_LOGIC0_43
    );
  PWR_GND_45_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_45_FROM
    );
  PWR_GND_45_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_45_GROM
    );
  PWR_GND_45_XUSED : X_BUF
    port map (
      I => PWR_GND_45_FROM,
      O => GLOBAL_LOGIC1_30
    );
  PWR_GND_45_YUSED : X_BUF
    port map (
      I => PWR_GND_45_GROM,
      O => GLOBAL_LOGIC0_44
    );
  PWR_GND_46_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_46_FROM
    );
  PWR_GND_46_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_46_GROM
    );
  PWR_GND_46_XUSED : X_BUF
    port map (
      I => PWR_GND_46_FROM,
      O => GLOBAL_LOGIC1_31
    );
  PWR_GND_46_YUSED : X_BUF
    port map (
      I => PWR_GND_46_GROM,
      O => GLOBAL_LOGIC0_45
    );
  PWR_GND_47_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_47_GROM
    );
  PWR_GND_47_YUSED : X_BUF
    port map (
      I => PWR_GND_47_GROM,
      O => GLOBAL_LOGIC0_46
    );
  PWR_GND_48_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_48_GROM
    );
  PWR_GND_48_YUSED : X_BUF
    port map (
      I => PWR_GND_48_GROM,
      O => GLOBAL_LOGIC0_47
    );
  PWR_GND_49_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_49_GROM
    );
  PWR_GND_49_YUSED : X_BUF
    port map (
      I => PWR_GND_49_GROM,
      O => GLOBAL_LOGIC0_48
    );
  PWR_GND_50_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_50_FROM
    );
  PWR_GND_50_G : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_50_GROM
    );
  PWR_GND_50_XUSED : X_BUF
    port map (
      I => PWR_GND_50_FROM,
      O => GLOBAL_LOGIC1_32
    );
  PWR_GND_50_YUSED : X_BUF
    port map (
      I => PWR_GND_50_GROM,
      O => GLOBAL_LOGIC0_49
    );
  PWR_VCC_0_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_0_FROM
    );
  PWR_VCC_0_XUSED : X_BUF
    port map (
      I => PWR_VCC_0_FROM,
      O => GLOBAL_LOGIC1_5
    );
  PWR_VCC_1_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_1_FROM
    );
  PWR_VCC_1_XUSED : X_BUF
    port map (
      I => PWR_VCC_1_FROM,
      O => GLOBAL_LOGIC1_6
    );
  PWR_VCC_2_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_2_FROM
    );
  PWR_VCC_2_XUSED : X_BUF
    port map (
      I => PWR_VCC_2_FROM,
      O => GLOBAL_LOGIC1_7
    );
  PWR_VCC_3_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_3_FROM
    );
  PWR_VCC_3_XUSED : X_BUF
    port map (
      I => PWR_VCC_3_FROM,
      O => GLOBAL_LOGIC1_8
    );
  PWR_VCC_4_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_4_FROM
    );
  PWR_VCC_4_XUSED : X_BUF
    port map (
      I => PWR_VCC_4_FROM,
      O => GLOBAL_LOGIC1_10
    );
  PWR_VCC_5_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_5_FROM
    );
  PWR_VCC_5_XUSED : X_BUF
    port map (
      I => PWR_VCC_5_FROM,
      O => GLOBAL_LOGIC1_12
    );
  PWR_VCC_6_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_6_FROM
    );
  PWR_VCC_6_XUSED : X_BUF
    port map (
      I => PWR_VCC_6_FROM,
      O => GLOBAL_LOGIC1_13
    );
  PWR_VCC_7_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_7_FROM
    );
  PWR_VCC_7_XUSED : X_BUF
    port map (
      I => PWR_VCC_7_FROM,
      O => GLOBAL_LOGIC1_15
    );
  PWR_VCC_8_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_8_FROM
    );
  PWR_VCC_8_XUSED : X_BUF
    port map (
      I => PWR_VCC_8_FROM,
      O => GLOBAL_LOGIC1_17
    );
  PWR_VCC_9_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_9_FROM
    );
  PWR_VCC_9_XUSED : X_BUF
    port map (
      I => PWR_VCC_9_FROM,
      O => GLOBAL_LOGIC1_18
    );
  PWR_VCC_10_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_10_FROM
    );
  PWR_VCC_10_XUSED : X_BUF
    port map (
      I => PWR_VCC_10_FROM,
      O => GLOBAL_LOGIC1_27
    );
  PWR_VCC_11_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_11_FROM
    );
  PWR_VCC_11_XUSED : X_BUF
    port map (
      I => PWR_VCC_11_FROM,
      O => GLOBAL_LOGIC1_28
    );
  PWR_VCC_12_F : X_LUT4
    generic map(
      INIT => X"FFFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_VCC_12_FROM
    );
  PWR_VCC_12_XUSED : X_BUF
    port map (
      I => PWR_VCC_12_FROM,
      O => GLOBAL_LOGIC1_33
    );
  NlwBlock_network_VCC : X_ONE
    port map (
      O => VCC
    );
  NlwBlock_network_GND : X_ZERO
    port map (
      O => GND
    );
  NlwBlockROC : X_ROC
    generic map (ROC_WIDTH => 100 ns)
    port map (O => GSR);
  NlwBlockTOC : X_TOC
    port map (O => GTS);

end Structure;

